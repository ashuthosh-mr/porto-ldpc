`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 25.11.2020 03:22:30
// Design Name: Check Node Processing
// Module Name: minmaxdecoding
// Project Name: ALPHA_INIT(v) + FB_init1
// Target Devices:
// Tool Versions: 1.0
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module minmaxdecoding(clk,reset,in, out,out_enable);


input clk;
input reset;
input [5:0]in;
output reg out_enable;
output reg[5:0] out;

reg[9:0]loop_var,l_v,l_v1,loop_var1,loop_var2, l_v2;

reg[9:0]col_row[255:0][2:0];
reg[5:0]H[255:0][383:0];
reg[3:0]inv_val[255:0],inv_val1[255:0];
reg[3:0]mul_val[255:0],mul_val1[255:0];

reg[5:0] state,next_state,cout;
reg[5:0]GAM,GAM1;
reg[9:0]row_state,col_state,row_state1,col_state1,address,row2,col2,row_ena,row_ena1,row1_ena,row1_ena1,col_ena,col_ena1;
reg[4:0] c,a_state1;
reg[3:0]address1;


reg[5:0]F[15:0][2:0][255:0];/////BASED ON RW AND CW
reg[5:0]B[15:0][2:0][255:0];


reg[5:0]F_[15:0][2:0][255:0];/////BASED ON RW AND CW
reg[5:0]B_[15:0][2:0][255:0];



reg[8:0]row_col[1:0][383:0];
reg alphaCSR[255:0][383:0];
//(* keep="true" *)reg[95:0] GAMMA[2:0];
reg reset1,reset_a;
reg enable,enable1,enable2,enable3,enable4,enable5,enable_copy,enable_even,enable_odd,enable_d1,enable_d2;
wire[12:0]reg_read_col,reg_read_a,count_copy;
wire[11:0]f_count,b_count;
wire[3:0]a_read_FB,a_write_FB;
wire[9:0]count_odd,count_even,count_d1,count_d2;

wire [3:0]count;
wire[4:0]bram_a;
reg enable_disable;
wire [9:0]bramid;
defparam gammain_counter.COUNT_LEN=4 ;
defparam counter3.COUNT_LEN=4 ;
defparam counter4.COUNT_LEN=4 ;
defparam counter5.COUNT_LEN=12 ;
defparam counter6.COUNT_LEN=12 ;
/*defparam  bram_out_a_counter.COUNT_LEN=5,bramid_counter.COUNT_LEN=10; */

/* counter_block bramid_counter(reset1,clk,enable1,bramid);
counter_block bram_out_a_counter(reset,clk,enable4,bram_a); */


counter_block gammain_counter(reset,clk,enable,count);
counter_block counter3(reset,clk,enable2,a_read_FB);
counter_block counter4(reset,clk,enable3,a_write_FB);
counter_block counter5(reset,clk,enable4,f_count);
counter_block counter6(reset,clk,enable5,b_count);


counter_even ce1(reset,clk,enable_even,count_even);
counter_odd co1(reset,clk,enable_odd,count_odd);

counter_disable_a d2(reset,clk,enable_d1,count_d1);
counter_disable_b d1(reset,clk,enable_d2,count_d2,enable_disable);

//counter_block gammain_counter_copy(reset,clk,enable_copy,count_copy);

  reg[3:0] addrA[767:0];
  reg[3:0] addrA_[767:0];
  reg weA[767:0];
  reg[5:0]dinA[767:0];
  wire[5:0]doutA[767:0];

 reg[3:0] addrA1[767:0];
  reg weA1[767:0];
  reg[5:0]dinA1[767:0];
  wire[5:0]doutA1[767:0];
  reg ena[767:0],enb[767:0];


  genvar i;
  generate
  for(i=0;i<768;i=i+1)
  begin
  blk_mem_gen_0 ALPHA (
    .clka(clk),    // input wire clka
    .ena(ena[i]),      // input wire ena
    .wea(weA[i]),      // input wire [0 : 0] wea
    .addra(addrA[i]),  // input wire [3 : 0] addra
    .dina(dinA[i]),    // input wire [5 : 0] dina
    .douta(doutA[i]),  // output wire [5 : 0] douta
    .clkb(clk),    // input wire clkb
    .enb(enb[i]),      // input wire enb
    .web(weA1[i]),      // input wire [0 : 0] web
    .addrb(addrA1[i]),  // input wire [3 : 0] addrb
    .dinb(dinA1[i]),    // input wire [5 : 0] dinb
    .doutb(doutA1[i])  // output wire [5 : 0] doutb
  );
  end
  endgenerate



`define RESET_STATE 6'd0
`define GAMMAIN0 6'd1
`define GAMMAIN1 6'd2
`define processing_state0 6'd3
`define processing_state1 6'd4
`define processing_state2 6'd5
`define FB_init1 6'd6
`define F_OUT 6'd7
`define B_OUT 6'd8
/* `define BRAM_OUT 6'D3
`define BRAM_OUT_WAIT0 6'd4
`define BRAM_OUT_WAIT1 6'd5
`define BRAM_OUT_WAIT2 6'd6
`define BRAM_OUT_WAIT3 6'd7
`define BETA_OUT 6'd8
`define ADD_CHECK 6'D9 */
`define END 6'd9




function[5:0] max;
    input[5:0] p,q;
    if(p<q) max=q;
    else max=p;
    endfunction

function[5:0] min;
        input[5:0] p,q;
        if(p<q) min=p;
        else min=q;
        endfunction


/* ALL THE TASKS ARE DEFINED BELOW*/
task mul_gf;// this one defines the multiplication for gf(16)
input[3:0] A;
input[3:0]B;
output [3:0]Y;
begin
Y={(A[3]&B[0])^(A[2]&B[1])^(A[1]&B[2])^(A[0]&B[3])^(A[3]&B[3]),(A[2]&B[0])^(A[1]&B[1])^(A[0]&B[2])^(A[3]&B[3])^(A[3]&B[2])^(A[2]&B[3]),(A[3]&B[2])^(A[3]&B[1])^(A[2]&B[3])^(A[2]&B[2])^(A[1]&B[3])^(A[1]&B[0])^(A[0]&B[1]),(A[1]&B[3])^(A[2]&B[2])^(A[3]&B[1])^(A[0]&B[0])};
end
endtask



task add_gf;// this one defines the addition for gf(16)
input[3:0] A;//this is simply xor operation of bits
input [3:0]Be;
output[3:0] out;
begin
out[0]=A[0]^Be[0];
out[1]=A[1]^Be[1];
out[2]=A[2]^Be[2];
out[3]=A[3]^Be[3];
end
endtask

task inv_gf;// this one defines the multiplication for gf(16)
input[3:0] A;
output [3:0]Y;
begin
case({A[3],A[2]})
2'd0: Y={A[1],A[1]&A[0],A[1]&A[0],((A[1]&(~A[0]))|((A[0]&(~A[1]))))};
2'd1: Y={~A[1],~A[0]|A[1],A[1]|A[0],~A[1]|(~A[0])};
2'd2: Y={~A[0],~A[0]|A[1],~A[1],~(A[1]^A[0])};
2'd3: Y={~(A[1]^A[0]),(~A[1])&A[0],~A[0],A[1]&(~A[0])};
endcase
end
endtask






//CODE TO REGISTER THE INPUT,IN
always@(posedge clk,posedge reset) begin
if(reset) begin
GAM=6'd0;
end
else begin
GAM=in;
end
end


/*
//BRAM_A ASSIGNEMENT
always@(state or reset)
begin
if(reset) enable4=1'b0;
else
begin
case(state)
`RESET_STATE: begin
enable4=1'b0;
end
`GAMMAIN0: begin
enable4=1'b0;
end

`BRAM_OUT: enable4=1'b1;


default: begin
enable4=0;
end

endcase
end
end

 */

//////// counter_odd
always@(state or reset)
begin
if(reset) enable_odd=1'b0;
else
begin
case(state)
`RESET_STATE: begin
enable_odd=1'b1;
end
`GAMMAIN0: begin
enable_odd=1'b0;
end
`GAMMAIN1: begin
enable_odd=1'b1;

end



default: begin
enable_odd=1'b0;
end

endcase
end
end


////counter_even
always@(state or reset)
begin
if(reset) enable_even=1'b0;
else
begin
case(state)
`RESET_STATE: begin
enable_even=1'b0;
end
`GAMMAIN0: begin
enable_even=1'b0;
end
`GAMMAIN1: begin
enable_even=1'b1;

end


default: begin
enable_even=1'b0;
end

endcase
end
end

//////counter_disable_a
always@(state or reset)
begin
if(reset) enable_d1=1'b0;
else
begin
case(state)
`RESET_STATE: begin
enable_d1=1'b1;
end
`GAMMAIN0: begin
enable_d1=1'b0;
end
`GAMMAIN1: begin
enable_d1=1'b1;

end



default: begin
enable_d1=1'b0;
end

endcase
end
end


/////counter_disable_b
always@(state or reset)
begin
if(reset) begin enable_d2=1'b0; enable_disable=1'b0; end
else
begin
case(state)
`RESET_STATE: begin
enable_d2=1'b1;
enable_disable=1'b0;
end
`GAMMAIN0: begin
enable_d2=1'b0;
enable_disable=1'b0;
end
`GAMMAIN1: begin
enable_d2=1'b1;
enable_disable=1'b1;
end



default: begin
enable_d2=1'b0;
enable_disable=1'b0;
end

endcase
end
end


//THIS IS FOR THE COUNTER REQD FOR GAMMAIN0
always@(state or reset)
begin
if(reset) enable=1'b0;
else
begin
case(state)
`RESET_STATE: begin
enable=1'b0;
end
`GAMMAIN0: begin
enable=1'b1;
end
`GAMMAIN1: begin
enable=1'b1;
end

default: begin
enable=1'b0;
end

endcase
end
end


//To make addrA a flip flop
always@(posedge clk or posedge reset) begin

if(reset) begin

for(l_v1=0;l_v1<768;l_v1=l_v1+1) begin
addrA_[l_v1]=4'd0;
end
end
else begin
for(l_v1=0;l_v1<768;l_v1=l_v1+1) begin
addrA_[l_v1]=addrA[l_v1];
end
end
end



// COUNTER TO READ FROM ALPHA FOR F/B_init1
always@(state or reset)
begin
if(reset) enable2=0;
else
begin
case(state)
`RESET_STATE: begin
enable2=0;
end
`GAMMAIN0: begin
enable2=0;
end
`processing_state0: begin
enable2=1;
end


`processing_state1: begin
enable2=1;
end
/*
`processing_state2: begin
enable2=1;
end
 */
`FB_init1: begin
enable2=1;
end

default: begin
enable2=0;
end

endcase
end
end


//COUNTER TO WRITE TO F/B
always@(state or reset)
begin
if(reset) enable3=0;
else
begin
case(state)
`RESET_STATE: begin
enable3=0;
end
`GAMMAIN0: begin
enable3=0;
end
`processing_state0: begin
enable3=0;
end


`processing_state1: begin
enable3=0;
end
/*
`processing_state2: begin
enable3=0;
end
 */
`FB_init1: begin
enable3=1;
end

default: begin
enable3=0;
end

endcase
end
end



//F_OUT COUNTER
always@(state or reset)
begin
if(reset) begin enable4=0;   end
else
begin
case(state)
`RESET_STATE: begin
enable4=0;
end
`F_OUT: begin
enable4=1;
end

default: begin
enable4=0;
end

endcase
end
end


//B_OUT COUNTER
always@(state or reset)
begin
if(reset) begin enable5=0;   end
else
begin
case(state)
`RESET_STATE: begin
enable5=0;
end
`B_OUT: begin
enable5=1;
end

default: begin
enable5=0;
end

endcase
end
end




/*
// RESET AND ENABLE FOR BRAMID COUNTER
always@(state or reset)
begin
if(reset) begin enable1=1'b0; reset1=1'b0;  end
else
begin
case(state)
`RESET_STATE: begin
enable1=1'b0;
reset1=1'b0;
end
`GAMMAIN0: begin
enable1=1'b0;
reset1=1'b1;
end

`BRAM_OUT_WAIT0: begin
reset1=1'b1;
enable1=1'b0;
end
`BRAM_OUT_WAIT1: begin
reset1=1'b0;
enable1=1'b0;
end
`BETA_OUT: begin
enable1=1'b1;
reset1=1'b0;
end

default: begin
enable1=1'b0;
reset1=1'b0;
end

endcase
end
end
 */


// ALWAYS BLOCK TO DETERMINE NEXT_STATE
always@(state,reset,count,bramid,bram_a,count_even,a_write_FB,f_count,b_count)
begin
if(reset)
begin
next_state=6'd0;
end
else begin
case(state)
`RESET_STATE: begin next_state=`GAMMAIN0; end
`GAMMAIN0: begin if(count==4'd14) begin next_state=`GAMMAIN1;  end else next_state=`GAMMAIN0; end
`GAMMAIN1: begin if(count_even==10'd766) begin next_state=`processing_state0; end else next_state=`GAMMAIN0; end
`processing_state0: begin next_state=`processing_state1; end
`processing_state1: begin next_state=`FB_init1; end
`FB_init1: begin if(a_write_FB==4'd15) next_state=`F_OUT; else begin next_state=`FB_init1; end   end
`F_OUT: begin if(f_count==12'b1111_1111_1111) next_state=`B_OUT; else next_state=`F_OUT;   end
`B_OUT: begin  if(b_count==12'b1111_1111_1111) next_state=`END; else next_state=`B_OUT; end






/* `BRAM_OUT: begin next_state=`BRAM_OUT_WAIT0;   end
`BRAM_OUT_WAIT0: begin  next_state=`BRAM_OUT_WAIT1;  end
`BRAM_OUT_WAIT1: begin  next_state=`BRAM_OUT_WAIT2;  end
`BRAM_OUT_WAIT2: begin  next_state=`BRAM_OUT_WAIT3;   end
`BRAM_OUT_WAIT3: begin next_state=`BETA_OUT; end
`BETA_OUT: begin if(bramid==10'b1_100_000_000) begin next_state=`ADD_CHECK;  end else next_state=`BETA_OUT; end
`ADD_CHECK: begin  if(bram_a==5'd16) next_state=`END; else next_state=`BRAM_OUT;  end
 */`END: begin   end
default: begin end
endcase
end
end

// to make F a flip flop
always@(posedge clk,posedge reset) begin
if(reset) begin
for(loop_var=0;loop_var<16;loop_var=loop_var+1) begin
for(loop_var1=0;loop_var1<3;loop_var1=loop_var1+1) begin
for(loop_var2=0;loop_var2<256;loop_var2=loop_var2+1) begin
F_[loop_var][loop_var1][loop_var2]=0;
end
end
end

end
else begin

for(loop_var=0;loop_var<16;loop_var=loop_var+1) begin
for(loop_var1=0;loop_var1<3;loop_var1=loop_var1+1) begin
for(loop_var2=0;loop_var2<256;loop_var2=loop_var2+1) begin
F_[loop_var][loop_var1][loop_var2]=F[loop_var][loop_var1][loop_var2];
end
end
end

end

end

//to make B a flip flop
always@(posedge clk,posedge reset) begin
if(reset) begin
for(loop_var=0;loop_var<16;loop_var=loop_var+1) begin
for(loop_var1=0;loop_var1<3;loop_var1=loop_var1+1) begin
for(loop_var2=0;loop_var2<256;loop_var2=loop_var2+1) begin
B_[loop_var][loop_var1][loop_var2]=0;
end
end
end

end
else begin

for(loop_var=0;loop_var<16;loop_var=loop_var+1) begin
for(loop_var1=0;loop_var1<3;loop_var1=loop_var1+1) begin
for(loop_var2=0;loop_var2<256;loop_var2=loop_var2+1) begin
B_[loop_var][loop_var1][loop_var2]=B[loop_var][loop_var1][loop_var2];
end
end
end

end

end


 // to enable and disable the brams as appropriate.
 always@(state,reset,count_even,count_odd,count_d1,count_d2) begin
 if(reset) begin
 for(l_v=0;l_v<768;l_v=l_v+1) begin
 ena[l_v]=1'b0;
 end
 end
 else begin
 case(state)
 `RESET_STATE: begin
  for(l_v=0;l_v<768;l_v=l_v+1) begin
 ena[l_v]=1'b0;
 end
 end
 `GAMMAIN0: begin
for(l_v=0;l_v<768;l_v=l_v+1) begin
if((l_v==count_even[9:0])||(l_v==count_odd[9:0]) ) begin
ena[l_v]=1'd1;
end
else
begin
ena[l_v]=1'd0;
end
end

 end
 `GAMMAIN1: begin
for(l_v=0;l_v<768;l_v=l_v+1) begin

 if((l_v==count_even[9:0])||(l_v==count_odd[9:0]) ) begin
 ena[l_v]=1'd1;
 end
 else
 begin
 ena[l_v]=1'd0;
 end
 end
 end

  `processing_state0: begin  for(l_v=0;l_v<768;l_v=l_v+1) begin ena[l_v]=1'b1;  end end
 `processing_state1: begin for(l_v=0;l_v<768;l_v=l_v+1) begin ena[l_v]=1'b1;  end  end
 `processing_state2: begin for(l_v=0;l_v<768;l_v=l_v+1) begin ena[l_v]=1'b1;  end  end
 `FB_init1: begin for(l_v=0;l_v<768;l_v=l_v+1) begin ena[l_v]=1'b1;  end  end
 `F_OUT: begin for(l_v=0;l_v<768;l_v=l_v+1) begin ena[l_v]=1'b1;  end  end
 `B_OUT: begin for(l_v=0;l_v<768;l_v=l_v+1) begin ena[l_v]=1'b1;  end  end





 default:
 begin
  for(l_v=0;l_v<768;l_v=l_v+1) begin
 ena[l_v]=1'b0;
 end

 end

 endcase
 end


 end



 // to enable and disable the brams PORT2 as appropriate.
 always@(state or reset) begin
 if(reset) begin
 for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin
 enb[l_v2]=1'b0;
 end
 end
 else begin
 case(state)
 `RESET_STATE: begin
  for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin
 enb[l_v2]=1'b0;
 end
 end
 `GAMMAIN0: begin
 for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin
 enb[l_v2]=1'b0;
 end
 end
 `GAMMAIN1: begin
 for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin
 enb[l_v2]=1'b0;
 end
 end

  `processing_state0: begin  for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin enb[l_v2]=1'b1;  end end
 `processing_state1: begin for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin enb[l_v2]=1'b1;  end  end
 `processing_state2: begin for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin enb[l_v2]=1'b1;  end  end
 `FB_init1: begin for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin enb[l_v2]=1'b1;  end  end
 `F_OUT: begin for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin enb[l_v2]=1'b1;  end  end
 `B_OUT: begin for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin enb[l_v2]=1'b1;  end  end





 default:
 begin
  for(l_v2=0;l_v2<768;l_v2=l_v2+1) begin
 enb[l_v2]=1'b0;
 end

 end

 endcase
 end


 end



// FUNCTIONALITY FOR EACH STATE
always@(state,reset,bramid,count,bram_a,GAM, count_even,count_odd,count_d1,count_d2,f_count,b_count,a_read_FB,a_write_FB,

row_col[1][ 0 ],
   row_col[0][ 1 ],
   row_col[1][ 1 ],
   row_col[0][ 2 ],
   row_col[1][ 2 ],
   row_col[0][ 3 ],
   row_col[1][ 3 ],
   row_col[0][ 4 ],
   row_col[1][ 4 ],
   row_col[0][ 5 ],
   row_col[1][ 5 ],
   row_col[0][ 6 ],
   row_col[1][ 6 ],
   row_col[0][ 7 ],
   row_col[1][ 7 ],
   row_col[0][ 8 ],
   row_col[1][ 8 ],
   row_col[0][ 9 ],
   row_col[1][ 9 ],
   row_col[0][ 10 ],
   row_col[1][ 10 ],
   row_col[0][ 11 ],
   row_col[1][ 11 ],
   row_col[0][ 12 ],
   row_col[1][ 12 ],
   row_col[0][ 13 ],
   row_col[1][ 13 ],
   row_col[0][ 14 ],
   row_col[1][ 14 ],
   row_col[0][ 15 ],
   row_col[1][ 15 ],
   row_col[0][ 16 ],
   row_col[1][ 16 ],
   row_col[0][ 17 ],
   row_col[1][ 17 ],
   row_col[0][ 18 ],
   row_col[1][ 18 ],
   row_col[0][ 19 ],
   row_col[1][ 19 ],
   row_col[0][ 20 ],
   row_col[1][ 20 ],
   row_col[0][ 21 ],
   row_col[1][ 21 ],
   row_col[0][ 22 ],
   row_col[1][ 22 ],
   row_col[0][ 23 ],
   row_col[1][ 23 ],
   row_col[0][ 24 ],
   row_col[1][ 24 ],
   row_col[0][ 25 ],
   row_col[1][ 25 ],
   row_col[0][ 26 ],
   row_col[1][ 26 ],
   row_col[0][ 27 ],
   row_col[1][ 27 ],
   row_col[0][ 28 ],
   row_col[1][ 28 ],
   row_col[0][ 29 ],
   row_col[1][ 29 ],
   row_col[0][ 30 ],
   row_col[1][ 30 ],
   row_col[0][ 31 ],
   row_col[1][ 31 ],
   row_col[0][ 32 ],
   row_col[1][ 32 ],
   row_col[0][ 33 ],
   row_col[1][ 33 ],
   row_col[0][ 34 ],
   row_col[1][ 34 ],
   row_col[0][ 35 ],
   row_col[1][ 35 ],
   row_col[0][ 36 ],
   row_col[1][ 36 ],
   row_col[0][ 37 ],
   row_col[1][ 37 ],
   row_col[0][ 38 ],
   row_col[1][ 38 ],
   row_col[0][ 39 ],
   row_col[1][ 39 ],
   row_col[0][ 40 ],
   row_col[1][ 40 ],
   row_col[0][ 41 ],
   row_col[1][ 41 ],
   row_col[0][ 42 ],
   row_col[1][ 42 ],
   row_col[0][ 43 ],
   row_col[1][ 43 ],
   row_col[0][ 44 ],
   row_col[1][ 44 ],
   row_col[0][ 45 ],
   row_col[1][ 45 ],
   row_col[0][ 46 ],
   row_col[1][ 46 ],
   row_col[0][ 47 ],
   row_col[1][ 47 ],
   row_col[0][ 48 ],
   row_col[1][ 48 ],
   row_col[0][ 49 ],
   row_col[1][ 49 ],
   row_col[0][ 50 ],
   row_col[1][ 50 ],
   row_col[0][ 51 ],
   row_col[1][ 51 ],
   row_col[0][ 52 ],
   row_col[1][ 52 ],
   row_col[0][ 53 ],
   row_col[1][ 53 ],
   row_col[0][ 54 ],
   row_col[1][ 54 ],
   row_col[0][ 55 ],
   row_col[1][ 55 ],
   row_col[0][ 56 ],
   row_col[1][ 56 ],
   row_col[0][ 57 ],
   row_col[1][ 57 ],
   row_col[0][ 58 ],
   row_col[1][ 58 ],
   row_col[0][ 59 ],
   row_col[1][ 59 ],
   row_col[0][ 60 ],
   row_col[1][ 60 ],
   row_col[0][ 61 ],
   row_col[1][ 61 ],
   row_col[0][ 62 ],
   row_col[1][ 62 ],
   row_col[0][ 63 ],
   row_col[1][ 63 ],
   row_col[0][ 64 ],
   row_col[1][ 64 ],
   row_col[0][ 65 ],
   row_col[1][ 65 ],
   row_col[0][ 66 ],
   row_col[1][ 66 ],
   row_col[0][ 67 ],
   row_col[1][ 67 ],
   row_col[0][ 68 ],
   row_col[1][ 68 ],
   row_col[0][ 69 ],
   row_col[1][ 69 ],
   row_col[0][ 70 ],
   row_col[1][ 70 ],
   row_col[0][ 71 ],
   row_col[1][ 71 ],
   row_col[0][ 72 ],
   row_col[1][ 72 ],
   row_col[0][ 73 ],
   row_col[1][ 73 ],
   row_col[0][ 74 ],
   row_col[1][ 74 ],
   row_col[0][ 75 ],
   row_col[1][ 75 ],
   row_col[0][ 76 ],
   row_col[1][ 76 ],
   row_col[0][ 77 ],
   row_col[1][ 77 ],
   row_col[0][ 78 ],
   row_col[1][ 78 ],
   row_col[0][ 79 ],
   row_col[1][ 79 ],
   row_col[0][ 80 ],
   row_col[1][ 80 ],
   row_col[0][ 81 ],
   row_col[1][ 81 ],
   row_col[0][ 82 ],
   row_col[1][ 82 ],
   row_col[0][ 83 ],
   row_col[1][ 83 ],
   row_col[0][ 84 ],
   row_col[1][ 84 ],
   row_col[0][ 85 ],
   row_col[1][ 85 ],
   row_col[0][ 86 ],
   row_col[1][ 86 ],
   row_col[0][ 87 ],
   row_col[1][ 87 ],
   row_col[0][ 88 ],
   row_col[1][ 88 ],
   row_col[0][ 89 ],
   row_col[1][ 89 ],
   row_col[0][ 90 ],
   row_col[1][ 90 ],
   row_col[0][ 91 ],
   row_col[1][ 91 ],
   row_col[0][ 92 ],
   row_col[1][ 92 ],
   row_col[0][ 93 ],
   row_col[1][ 93 ],
   row_col[0][ 94 ],
   row_col[1][ 94 ],
   row_col[0][ 95 ],
   row_col[1][ 95 ],
   row_col[0][ 96 ],
   row_col[1][ 96 ],
   row_col[0][ 97 ],
   row_col[1][ 97 ],
   row_col[0][ 98 ],
   row_col[1][ 98 ],
   row_col[0][ 99 ],
   row_col[1][ 99 ],
   row_col[0][ 100 ],
   row_col[1][ 100 ],
   row_col[0][ 101 ],
   row_col[1][ 101 ],
   row_col[0][ 102 ],
   row_col[1][ 102 ],
   row_col[0][ 103 ],
   row_col[1][ 103 ],
   row_col[0][ 104 ],
   row_col[1][ 104 ],
   row_col[0][ 105 ],
   row_col[1][ 105 ],
   row_col[0][ 106 ],
   row_col[1][ 106 ],
   row_col[0][ 107 ],
   row_col[1][ 107 ],
   row_col[0][ 108 ],
   row_col[1][ 108 ],
   row_col[0][ 109 ],
   row_col[1][ 109 ],
   row_col[0][ 110 ],
   row_col[1][ 110 ],
   row_col[0][ 111 ],
   row_col[1][ 111 ],
   row_col[0][ 112 ],
   row_col[1][ 112 ],
   row_col[0][ 113 ],
   row_col[1][ 113 ],
   row_col[0][ 114 ],
   row_col[1][ 114 ],
   row_col[0][ 115 ],
   row_col[1][ 115 ],
   row_col[0][ 116 ],
   row_col[1][ 116 ],
   row_col[0][ 117 ],
   row_col[1][ 117 ],
   row_col[0][ 118 ],
   row_col[1][ 118 ],
   row_col[0][ 119 ],
   row_col[1][ 119 ],
   row_col[0][ 120 ],
   row_col[1][ 120 ],
   row_col[0][ 121 ],
   row_col[1][ 121 ],
   row_col[0][ 122 ],
   row_col[1][ 122 ],
   row_col[0][ 123 ],
   row_col[1][ 123 ],
   row_col[0][ 124 ],
   row_col[1][ 124 ],
   row_col[0][ 125 ],
   row_col[1][ 125 ],
   row_col[0][ 126 ],
   row_col[1][ 126 ],
   row_col[0][ 127 ],
   row_col[1][ 127 ],
   row_col[0][ 128 ],
   row_col[1][ 128 ],
   row_col[0][ 129 ],
   row_col[1][ 129 ],
   row_col[0][ 130 ],
   row_col[1][ 130 ],
   row_col[0][ 131 ],
   row_col[1][ 131 ],
   row_col[0][ 132 ],
   row_col[1][ 132 ],
   row_col[0][ 133 ],
   row_col[1][ 133 ],
   row_col[0][ 134 ],
   row_col[1][ 134 ],
   row_col[0][ 135 ],
   row_col[1][ 135 ],
   row_col[0][ 136 ],
   row_col[1][ 136 ],
   row_col[0][ 137 ],
   row_col[1][ 137 ],
   row_col[0][ 138 ],
   row_col[1][ 138 ],
   row_col[0][ 139 ],
   row_col[1][ 139 ],
   row_col[0][ 140 ],
   row_col[1][ 140 ],
   row_col[0][ 141 ],
   row_col[1][ 141 ],
   row_col[0][ 142 ],
   row_col[1][ 142 ],
   row_col[0][ 143 ],
   row_col[1][ 143 ],
   row_col[0][ 144 ],
   row_col[1][ 144 ],
   row_col[0][ 145 ],
   row_col[1][ 145 ],
   row_col[0][ 146 ],
   row_col[1][ 146 ],
   row_col[0][ 147 ],
   row_col[1][ 147 ],
   row_col[0][ 148 ],
   row_col[1][ 148 ],
   row_col[0][ 149 ],
   row_col[1][ 149 ],
   row_col[0][ 150 ],
   row_col[1][ 150 ],
   row_col[0][ 151 ],
   row_col[1][ 151 ],
   row_col[0][ 152 ],
   row_col[1][ 152 ],
   row_col[0][ 153 ],
   row_col[1][ 153 ],
   row_col[0][ 154 ],
   row_col[1][ 154 ],
   row_col[0][ 155 ],
   row_col[1][ 155 ],
   row_col[0][ 156 ],
   row_col[1][ 156 ],
   row_col[0][ 157 ],
   row_col[1][ 157 ],
   row_col[0][ 158 ],
   row_col[1][ 158 ],
   row_col[0][ 159 ],
   row_col[1][ 159 ],
   row_col[0][ 160 ],
   row_col[1][ 160 ],
   row_col[0][ 161 ],
   row_col[1][ 161 ],
   row_col[0][ 162 ],
   row_col[1][ 162 ],
   row_col[0][ 163 ],
   row_col[1][ 163 ],
   row_col[0][ 164 ],
   row_col[1][ 164 ],
   row_col[0][ 165 ],
   row_col[1][ 165 ],
   row_col[0][ 166 ],
   row_col[1][ 166 ],
   row_col[0][ 167 ],
   row_col[1][ 167 ],
   row_col[0][ 168 ],
   row_col[1][ 168 ],
   row_col[0][ 169 ],
   row_col[1][ 169 ],
   row_col[0][ 170 ],
   row_col[1][ 170 ],
   row_col[0][ 171 ],
   row_col[1][ 171 ],
   row_col[0][ 172 ],
   row_col[1][ 172 ],
   row_col[0][ 173 ],
   row_col[1][ 173 ],
   row_col[0][ 174 ],
   row_col[1][ 174 ],
   row_col[0][ 175 ],
   row_col[1][ 175 ],
   row_col[0][ 176 ],
   row_col[1][ 176 ],
   row_col[0][ 177 ],
   row_col[1][ 177 ],
   row_col[0][ 178 ],
   row_col[1][ 178 ],
   row_col[0][ 179 ],
   row_col[1][ 179 ],
   row_col[0][ 180 ],
   row_col[1][ 180 ],
   row_col[0][ 181 ],
   row_col[1][ 181 ],
   row_col[0][ 182 ],
   row_col[1][ 182 ],
   row_col[0][ 183 ],
   row_col[1][ 183 ],
   row_col[0][ 184 ],
   row_col[1][ 184 ],
   row_col[0][ 185 ],
   row_col[1][ 185 ],
   row_col[0][ 186 ],
   row_col[1][ 186 ],
   row_col[0][ 187 ],
   row_col[1][ 187 ],
   row_col[0][ 188 ],
   row_col[1][ 188 ],
   row_col[0][ 189 ],
   row_col[1][ 189 ],
   row_col[0][ 190 ],
   row_col[1][ 190 ],
   row_col[0][ 191 ],
   row_col[1][ 191 ],
   row_col[0][ 192 ],
   row_col[1][ 192 ],
   row_col[0][ 193 ],
   row_col[1][ 193 ],
   row_col[0][ 194 ],
   row_col[1][ 194 ],
   row_col[0][ 195 ],
   row_col[1][ 195 ],
   row_col[0][ 196 ],
   row_col[1][ 196 ],
   row_col[0][ 197 ],
   row_col[1][ 197 ],
   row_col[0][ 198 ],
   row_col[1][ 198 ],
   row_col[0][ 199 ],
   row_col[1][ 199 ],
   row_col[0][ 200 ],
   row_col[1][ 200 ],
   row_col[0][ 201 ],
   row_col[1][ 201 ],
   row_col[0][ 202 ],
   row_col[1][ 202 ],
   row_col[0][ 203 ],
   row_col[1][ 203 ],
   row_col[0][ 204 ],
   row_col[1][ 204 ],
   row_col[0][ 205 ],
   row_col[1][ 205 ],
   row_col[0][ 206 ],
   row_col[1][ 206 ],
   row_col[0][ 207 ],
   row_col[1][ 207 ],
   row_col[0][ 208 ],
   row_col[1][ 208 ],
   row_col[0][ 209 ],
   row_col[1][ 209 ],
   row_col[0][ 210 ],
   row_col[1][ 210 ],
   row_col[0][ 211 ],
   row_col[1][ 211 ],
   row_col[0][ 212 ],
   row_col[1][ 212 ],
   row_col[0][ 213 ],
   row_col[1][ 213 ],
   row_col[0][ 214 ],
   row_col[1][ 214 ],
   row_col[0][ 215 ],
   row_col[1][ 215 ],
   row_col[0][ 216 ],
   row_col[1][ 216 ],
   row_col[0][ 217 ],
   row_col[1][ 217 ],
   row_col[0][ 218 ],
   row_col[1][ 218 ],
   row_col[0][ 219 ],
   row_col[1][ 219 ],
   row_col[0][ 220 ],
   row_col[1][ 220 ],
   row_col[0][ 221 ],
   row_col[1][ 221 ],
   row_col[0][ 222 ],
   row_col[1][ 222 ],
   row_col[0][ 223 ],
   row_col[1][ 223 ],
   row_col[0][ 224 ],
   row_col[1][ 224 ],
   row_col[0][ 225 ],
   row_col[1][ 225 ],
   row_col[0][ 226 ],
   row_col[1][ 226 ],
   row_col[0][ 227 ],
   row_col[1][ 227 ],
   row_col[0][ 228 ],
   row_col[1][ 228 ],
   row_col[0][ 229 ],
   row_col[1][ 229 ],
   row_col[0][ 230 ],
   row_col[1][ 230 ],
   row_col[0][ 231 ],
   row_col[1][ 231 ],
   row_col[0][ 232 ],
   row_col[1][ 232 ],
   row_col[0][ 233 ],
   row_col[1][ 233 ],
   row_col[0][ 234 ],
   row_col[1][ 234 ],
   row_col[0][ 235 ],
   row_col[1][ 235 ],
   row_col[0][ 236 ],
   row_col[1][ 236 ],
   row_col[0][ 237 ],
   row_col[1][ 237 ],
   row_col[0][ 238 ],
   row_col[1][ 238 ],
   row_col[0][ 239 ],
   row_col[1][ 239 ],
   row_col[0][ 240 ],
   row_col[1][ 240 ],
   row_col[0][ 241 ],
   row_col[1][ 241 ],
   row_col[0][ 242 ],
   row_col[1][ 242 ],
   row_col[0][ 243 ],
   row_col[1][ 243 ],
   row_col[0][ 244 ],
   row_col[1][ 244 ],
   row_col[0][ 245 ],
   row_col[1][ 245 ],
   row_col[0][ 246 ],
   row_col[1][ 246 ],
   row_col[0][ 247 ],
   row_col[1][ 247 ],
   row_col[0][ 248 ],
   row_col[1][ 248 ],
   row_col[0][ 249 ],
   row_col[1][ 249 ],
   row_col[0][ 250 ],
   row_col[1][ 250 ],
   row_col[0][ 251 ],
   row_col[1][ 251 ],
   row_col[0][ 252 ],
   row_col[1][ 252 ],
   row_col[0][ 253 ],
   row_col[1][ 253 ],
   row_col[0][ 254 ],
   row_col[1][ 254 ],
   row_col[0][ 255 ],
   row_col[1][ 255 ],
   row_col[0][ 256 ],
   row_col[1][ 256 ],
   row_col[0][ 257 ],
   row_col[1][ 257 ],
   row_col[0][ 258 ],
   row_col[1][ 258 ],
   row_col[0][ 259 ],
   row_col[1][ 259 ],
   row_col[0][ 260 ],
   row_col[1][ 260 ],
   row_col[0][ 261 ],
   row_col[1][ 261 ],
   row_col[0][ 262 ],
   row_col[1][ 262 ],
   row_col[0][ 263 ],
   row_col[1][ 263 ],
   row_col[0][ 264 ],
   row_col[1][ 264 ],
   row_col[0][ 265 ],
   row_col[1][ 265 ],
   row_col[0][ 266 ],
   row_col[1][ 266 ],
   row_col[0][ 267 ],
   row_col[1][ 267 ],
   row_col[0][ 268 ],
   row_col[1][ 268 ],
   row_col[0][ 269 ],
   row_col[1][ 269 ],
   row_col[0][ 270 ],
   row_col[1][ 270 ],
   row_col[0][ 271 ],
   row_col[1][ 271 ],
   row_col[0][ 272 ],
   row_col[1][ 272 ],
   row_col[0][ 273 ],
   row_col[1][ 273 ],
   row_col[0][ 274 ],
   row_col[1][ 274 ],
   row_col[0][ 275 ],
   row_col[1][ 275 ],
   row_col[0][ 276 ],
   row_col[1][ 276 ],
   row_col[0][ 277 ],
   row_col[1][ 277 ],
   row_col[0][ 278 ],
   row_col[1][ 278 ],
   row_col[0][ 279 ],
   row_col[1][ 279 ],
   row_col[0][ 280 ],
   row_col[1][ 280 ],
   row_col[0][ 281 ],
   row_col[1][ 281 ],
   row_col[0][ 282 ],
   row_col[1][ 282 ],
   row_col[0][ 283 ],
   row_col[1][ 283 ],
   row_col[0][ 284 ],
   row_col[1][ 284 ],
   row_col[0][ 285 ],
   row_col[1][ 285 ],
   row_col[0][ 286 ],
   row_col[1][ 286 ],
   row_col[0][ 287 ],
   row_col[1][ 287 ],
   row_col[0][ 288 ],
   row_col[1][ 288 ],
   row_col[0][ 289 ],
   row_col[1][ 289 ],
   row_col[0][ 290 ],
   row_col[1][ 290 ],
   row_col[0][ 291 ],
   row_col[1][ 291 ],
   row_col[0][ 292 ],
   row_col[1][ 292 ],
   row_col[0][ 293 ],
   row_col[1][ 293 ],
   row_col[0][ 294 ],
   row_col[1][ 294 ],
   row_col[0][ 295 ],
   row_col[1][ 295 ],
   row_col[0][ 296 ],
   row_col[1][ 296 ],
   row_col[0][ 297 ],
   row_col[1][ 297 ],
   row_col[0][ 298 ],
   row_col[1][ 298 ],
   row_col[0][ 299 ],
   row_col[1][ 299 ],
   row_col[0][ 300 ],
   row_col[1][ 300 ],
   row_col[0][ 301 ],
   row_col[1][ 301 ],
   row_col[0][ 302 ],
   row_col[1][ 302 ],
   row_col[0][ 303 ],
   row_col[1][ 303 ],
   row_col[0][ 304 ],
   row_col[1][ 304 ],
   row_col[0][ 305 ],
   row_col[1][ 305 ],
   row_col[0][ 306 ],
   row_col[1][ 306 ],
   row_col[0][ 307 ],
   row_col[1][ 307 ],
   row_col[0][ 308 ],
   row_col[1][ 308 ],
   row_col[0][ 309 ],
   row_col[1][ 309 ],
   row_col[0][ 310 ],
   row_col[1][ 310 ],
   row_col[0][ 311 ],
   row_col[1][ 311 ],
   row_col[0][ 312 ],
   row_col[1][ 312 ],
   row_col[0][ 313 ],
   row_col[1][ 313 ],
   row_col[0][ 314 ],
   row_col[1][ 314 ],
   row_col[0][ 315 ],
   row_col[1][ 315 ],
   row_col[0][ 316 ],
   row_col[1][ 316 ],
   row_col[0][ 317 ],
   row_col[1][ 317 ],
   row_col[0][ 318 ],
   row_col[1][ 318 ],
   row_col[0][ 319 ],
   row_col[1][ 319 ],
   row_col[0][ 320 ],
   row_col[1][ 320 ],
   row_col[0][ 321 ],
   row_col[1][ 321 ],
   row_col[0][ 322 ],
   row_col[1][ 322 ],
   row_col[0][ 323 ],
   row_col[1][ 323 ],
   row_col[0][ 324 ],
   row_col[1][ 324 ],
   row_col[0][ 325 ],
   row_col[1][ 325 ],
   row_col[0][ 326 ],
   row_col[1][ 326 ],
   row_col[0][ 327 ],
   row_col[1][ 327 ],
   row_col[0][ 328 ],
   row_col[1][ 328 ],
   row_col[0][ 329 ],
   row_col[1][ 329 ],
   row_col[0][ 330 ],
   row_col[1][ 330 ],
   row_col[0][ 331 ],
   row_col[1][ 331 ],
   row_col[0][ 332 ],
   row_col[1][ 332 ],
   row_col[0][ 333 ],
   row_col[1][ 333 ],
   row_col[0][ 334 ],
   row_col[1][ 334 ],
   row_col[0][ 335 ],
   row_col[1][ 335 ],
   row_col[0][ 336 ],
   row_col[1][ 336 ],
   row_col[0][ 337 ],
   row_col[1][ 337 ],
   row_col[0][ 338 ],
   row_col[1][ 338 ],
   row_col[0][ 339 ],
   row_col[1][ 339 ],
   row_col[0][ 340 ],
   row_col[1][ 340 ],
   row_col[0][ 341 ],
   row_col[1][ 341 ],
   row_col[0][ 342 ],
   row_col[1][ 342 ],
   row_col[0][ 343 ],
   row_col[1][ 343 ],
   row_col[0][ 344 ],
   row_col[1][ 344 ],
   row_col[0][ 345 ],
   row_col[1][ 345 ],
   row_col[0][ 346 ],
   row_col[1][ 346 ],
   row_col[0][ 347 ],
   row_col[1][ 347 ],
   row_col[0][ 348 ],
   row_col[1][ 348 ],
   row_col[0][ 349 ],
   row_col[1][ 349 ],
   row_col[0][ 350 ],
   row_col[1][ 350 ],
   row_col[0][ 351 ],
   row_col[1][ 351 ],
   row_col[0][ 352 ],
   row_col[1][ 352 ],
   row_col[0][ 353 ],
   row_col[1][ 353 ],
   row_col[0][ 354 ],
   row_col[1][ 354 ],
   row_col[0][ 355 ],
   row_col[1][ 355 ],
   row_col[0][ 356 ],
   row_col[1][ 356 ],
   row_col[0][ 357 ],
   row_col[1][ 357 ],
   row_col[0][ 358 ],
   row_col[1][ 358 ],
   row_col[0][ 359 ],
   row_col[1][ 359 ],
   row_col[0][ 360 ],
   row_col[1][ 360 ],
   row_col[0][ 361 ],
   row_col[1][ 361 ],
   row_col[0][ 362 ],
   row_col[1][ 362 ],
   row_col[0][ 363 ],
   row_col[1][ 363 ],
   row_col[0][ 364 ],
   row_col[1][ 364 ],
   row_col[0][ 365 ],
   row_col[1][ 365 ],
   row_col[0][ 366 ],
   row_col[1][ 366 ],
   row_col[0][ 367 ],
   row_col[1][ 367 ],
   row_col[0][ 368 ],
   row_col[1][ 368 ],
   row_col[0][ 369 ],
   row_col[1][ 369 ],
   row_col[0][ 370 ],
   row_col[1][ 370 ],
   row_col[0][ 371 ],
   row_col[1][ 371 ],
   row_col[0][ 372 ],
   row_col[1][ 372 ],
   row_col[0][ 373 ],
   row_col[1][ 373 ],
   row_col[0][ 374 ],
   row_col[1][ 374 ],
   row_col[0][ 375 ],
   row_col[1][ 375 ],
   row_col[0][ 376 ],
   row_col[1][ 376 ],
   row_col[0][ 377 ],
   row_col[1][ 377 ],
   row_col[0][ 378 ],
   row_col[1][ 378 ],
   row_col[0][ 379 ],
   row_col[1][ 379 ],
   row_col[0][ 380 ],
   row_col[1][ 380 ],
   row_col[0][ 381 ],
   row_col[1][ 381 ],
   row_col[0][ 382 ],
   row_col[1][ 382 ],
   row_col[0][383],
   row_col[1][383],
   alphaCSR[ 0 ][ 0 ],
   alphaCSR[ 0 ][ 1 ],
   alphaCSR[ 0 ][ 2 ],
   alphaCSR[ 0 ][ 3 ],
   alphaCSR[ 0 ][ 4 ],
   alphaCSR[ 0 ][ 5 ],
   alphaCSR[ 0 ][ 6 ],
   alphaCSR[ 0 ][ 7 ],
   alphaCSR[ 0 ][ 8 ],
   alphaCSR[ 0 ][ 9 ],
   alphaCSR[ 0 ][ 10 ],
   alphaCSR[ 0 ][ 11 ],
   alphaCSR[ 0 ][ 12 ],
   alphaCSR[ 0 ][ 13 ],
   alphaCSR[ 0 ][ 14 ],
   alphaCSR[ 0 ][ 15 ],
   alphaCSR[ 0 ][ 16 ],
   alphaCSR[ 0 ][ 17 ],
   alphaCSR[ 0 ][ 18 ],
   alphaCSR[ 0 ][ 19 ],
   alphaCSR[ 0 ][ 20 ],
   alphaCSR[ 0 ][ 21 ],
   alphaCSR[ 0 ][ 22 ],
   alphaCSR[ 0 ][ 23 ],
   alphaCSR[ 0 ][ 24 ],
   alphaCSR[ 0 ][ 25 ],
   alphaCSR[ 0 ][ 26 ],
   alphaCSR[ 0 ][ 27 ],
   alphaCSR[ 0 ][ 28 ],
   alphaCSR[ 0 ][ 29 ],
   alphaCSR[ 0 ][ 30 ],
   alphaCSR[ 0 ][ 31 ],
   alphaCSR[ 0 ][ 32 ],
   alphaCSR[ 0 ][ 33 ],
   alphaCSR[ 0 ][ 34 ],
   alphaCSR[ 0 ][ 35 ],
   alphaCSR[ 0 ][ 36 ],
   alphaCSR[ 0 ][ 37 ],
   alphaCSR[ 0 ][ 38 ],
   alphaCSR[ 0 ][ 39 ],
   alphaCSR[ 0 ][ 40 ],
   alphaCSR[ 0 ][ 41 ],
   alphaCSR[ 0 ][ 42 ],
   alphaCSR[ 0 ][ 43 ],
   alphaCSR[ 0 ][ 44 ],
   alphaCSR[ 0 ][ 45 ],
   alphaCSR[ 0 ][ 46 ],
   alphaCSR[ 0 ][ 47 ],
   alphaCSR[ 0 ][ 48 ],
   alphaCSR[ 0 ][ 49 ],
   alphaCSR[ 0 ][ 50 ],
   alphaCSR[ 0 ][ 51 ],
   alphaCSR[ 0 ][ 52 ],
   alphaCSR[ 0 ][ 53 ],
   alphaCSR[ 0 ][ 54 ],
   alphaCSR[ 0 ][ 55 ],
   alphaCSR[ 0 ][ 56 ],
   alphaCSR[ 0 ][ 57 ],
   alphaCSR[ 0 ][ 58 ],
   alphaCSR[ 0 ][ 59 ],
   alphaCSR[ 0 ][ 60 ],
   alphaCSR[ 0 ][ 61 ],
   alphaCSR[ 0 ][ 62 ],
   alphaCSR[ 0 ][ 63 ],
   alphaCSR[ 0 ][ 64 ],
   alphaCSR[ 0 ][ 65 ],
   alphaCSR[ 0 ][ 66 ],
   alphaCSR[ 0 ][ 67 ],
   alphaCSR[ 0 ][ 68 ],
   alphaCSR[ 0 ][ 69 ],
   alphaCSR[ 0 ][ 70 ],
   alphaCSR[ 0 ][ 71 ],
   alphaCSR[ 0 ][ 72 ],
   alphaCSR[ 0 ][ 73 ],
   alphaCSR[ 0 ][ 74 ],
   alphaCSR[ 0 ][ 75 ],
   alphaCSR[ 0 ][ 76 ],
   alphaCSR[ 0 ][ 77 ],
   alphaCSR[ 0 ][ 78 ],
   alphaCSR[ 0 ][ 79 ],
   alphaCSR[ 0 ][ 80 ],
   alphaCSR[ 0 ][ 81 ],
   alphaCSR[ 0 ][ 82 ],
   alphaCSR[ 0 ][ 83 ],
   alphaCSR[ 0 ][ 84 ],
   alphaCSR[ 0 ][ 85 ],
   alphaCSR[ 0 ][ 86 ],
   alphaCSR[ 0 ][ 87 ],
   alphaCSR[ 0 ][ 88 ],
   alphaCSR[ 0 ][ 89 ],
   alphaCSR[ 0 ][ 90 ],
   alphaCSR[ 0 ][ 91 ],
   alphaCSR[ 0 ][ 92 ],
   alphaCSR[ 0 ][ 93 ],
   alphaCSR[ 0 ][ 94 ],
   alphaCSR[ 0 ][ 95 ],
   alphaCSR[ 0 ][ 96 ],
   alphaCSR[ 0 ][ 97 ],
   alphaCSR[ 0 ][ 98 ],
   alphaCSR[ 0 ][ 99 ],
   alphaCSR[ 0 ][ 100 ],
   alphaCSR[ 0 ][ 101 ],
   alphaCSR[ 0 ][ 102 ],
   alphaCSR[ 0 ][ 103 ],
   alphaCSR[ 0 ][ 104 ],
   alphaCSR[ 0 ][ 105 ],
   alphaCSR[ 0 ][ 106 ],
   alphaCSR[ 0 ][ 107 ],
   alphaCSR[ 0 ][ 108 ],
   alphaCSR[ 0 ][ 109 ],
   alphaCSR[ 0 ][ 110 ],
   alphaCSR[ 0 ][ 111 ],
   alphaCSR[ 0 ][ 112 ],
   alphaCSR[ 0 ][ 113 ],
   alphaCSR[ 0 ][ 114 ],
   alphaCSR[ 0 ][ 115 ],
   alphaCSR[ 0 ][ 116 ],
   alphaCSR[ 0 ][ 117 ],
   alphaCSR[ 0 ][ 118 ],
   alphaCSR[ 0 ][ 119 ],
   alphaCSR[ 0 ][ 120 ],
   alphaCSR[ 0 ][ 121 ],
   alphaCSR[ 0 ][ 122 ],
   alphaCSR[ 0 ][ 123 ],
   alphaCSR[ 0 ][ 124 ],
   alphaCSR[ 0 ][ 125 ],
   alphaCSR[ 0 ][ 126 ],
   alphaCSR[ 0 ][ 127 ],
   alphaCSR[ 0 ][ 128 ],
   alphaCSR[ 0 ][ 129 ],
   alphaCSR[ 0 ][ 130 ],
   alphaCSR[ 0 ][ 131 ],
   alphaCSR[ 0 ][ 132 ],
   alphaCSR[ 0 ][ 133 ],
   alphaCSR[ 0 ][ 134 ],
   alphaCSR[ 0 ][ 135 ],
   alphaCSR[ 0 ][ 136 ],
   alphaCSR[ 0 ][ 137 ],
   alphaCSR[ 0 ][ 138 ],
   alphaCSR[ 0 ][ 139 ],
   alphaCSR[ 0 ][ 140 ],
   alphaCSR[ 0 ][ 141 ],
   alphaCSR[ 0 ][ 142 ],
   alphaCSR[ 0 ][ 143 ],
   alphaCSR[ 0 ][ 144 ],
   alphaCSR[ 0 ][ 145 ],
   alphaCSR[ 0 ][ 146 ],
   alphaCSR[ 0 ][ 147 ],
   alphaCSR[ 0 ][ 148 ],
   alphaCSR[ 0 ][ 149 ],
   alphaCSR[ 0 ][ 150 ],
   alphaCSR[ 0 ][ 151 ],
   alphaCSR[ 0 ][ 152 ],
   alphaCSR[ 0 ][ 153 ],
   alphaCSR[ 0 ][ 154 ],
   alphaCSR[ 0 ][ 155 ],
   alphaCSR[ 0 ][ 156 ],
   alphaCSR[ 0 ][ 157 ],
   alphaCSR[ 0 ][ 158 ],
   alphaCSR[ 0 ][ 159 ],
   alphaCSR[ 0 ][ 160 ],
   alphaCSR[ 0 ][ 161 ],
   alphaCSR[ 0 ][ 162 ],
   alphaCSR[ 0 ][ 163 ],
   alphaCSR[ 0 ][ 164 ],
   alphaCSR[ 0 ][ 165 ],
   alphaCSR[ 0 ][ 166 ],
   alphaCSR[ 0 ][ 167 ],
   alphaCSR[ 0 ][ 168 ],
   alphaCSR[ 0 ][ 169 ],
   alphaCSR[ 0 ][ 170 ],
   alphaCSR[ 0 ][ 171 ],
   alphaCSR[ 0 ][ 172 ],
   alphaCSR[ 0 ][ 173 ],
   alphaCSR[ 0 ][ 174 ],
   alphaCSR[ 0 ][ 175 ],
   alphaCSR[ 0 ][ 176 ],
   alphaCSR[ 0 ][ 177 ],
   alphaCSR[ 0 ][ 178 ],
   alphaCSR[ 0 ][ 179 ],
   alphaCSR[ 0 ][ 180 ],
   alphaCSR[ 0 ][ 181 ],
   alphaCSR[ 0 ][ 182 ],
   alphaCSR[ 0 ][ 183 ],
   alphaCSR[ 0 ][ 184 ],
   alphaCSR[ 0 ][ 185 ],
   alphaCSR[ 0 ][ 186 ],
   alphaCSR[ 0 ][ 187 ],
   alphaCSR[ 0 ][ 188 ],
   alphaCSR[ 0 ][ 189 ],
   alphaCSR[ 0 ][ 190 ],
   alphaCSR[ 0 ][ 191 ],
   alphaCSR[ 0 ][ 192 ],
   alphaCSR[ 0 ][ 193 ],
   alphaCSR[ 0 ][ 194 ],
   alphaCSR[ 0 ][ 195 ],
   alphaCSR[ 0 ][ 196 ],
   alphaCSR[ 0 ][ 197 ],
   alphaCSR[ 0 ][ 198 ],
   alphaCSR[ 0 ][ 199 ],
   alphaCSR[ 0 ][ 200 ],
   alphaCSR[ 0 ][ 201 ],
   alphaCSR[ 0 ][ 202 ],
   alphaCSR[ 0 ][ 203 ],
   alphaCSR[ 0 ][ 204 ],
   alphaCSR[ 0 ][ 205 ],
   alphaCSR[ 0 ][ 206 ],
   alphaCSR[ 0 ][ 207 ],
   alphaCSR[ 0 ][ 208 ],
   alphaCSR[ 0 ][ 209 ],
   alphaCSR[ 0 ][ 210 ],
   alphaCSR[ 0 ][ 211 ],
   alphaCSR[ 0 ][ 212 ],
   alphaCSR[ 0 ][ 213 ],
   alphaCSR[ 0 ][ 214 ],
   alphaCSR[ 0 ][ 215 ],
   alphaCSR[ 0 ][ 216 ],
   alphaCSR[ 0 ][ 217 ],
   alphaCSR[ 0 ][ 218 ],
   alphaCSR[ 0 ][ 219 ],
   alphaCSR[ 0 ][ 220 ],
   alphaCSR[ 0 ][ 221 ],
   alphaCSR[ 0 ][ 222 ],
   alphaCSR[ 0 ][ 223 ],
   alphaCSR[ 0 ][ 224 ],
   alphaCSR[ 0 ][ 225 ],
   alphaCSR[ 0 ][ 226 ],
   alphaCSR[ 0 ][ 227 ],
   alphaCSR[ 0 ][ 228 ],
   alphaCSR[ 0 ][ 229 ],
   alphaCSR[ 0 ][ 230 ],
   alphaCSR[ 0 ][ 231 ],
   alphaCSR[ 0 ][ 232 ],
   alphaCSR[ 0 ][ 233 ],
   alphaCSR[ 0 ][ 234 ],
   alphaCSR[ 0 ][ 235 ],
   alphaCSR[ 0 ][ 236 ],
   alphaCSR[ 0 ][ 237 ],
   alphaCSR[ 0 ][ 238 ],
   alphaCSR[ 0 ][ 239 ],
   alphaCSR[ 0 ][ 240 ],
   alphaCSR[ 0 ][ 241 ],
   alphaCSR[ 0 ][ 242 ],
   alphaCSR[ 0 ][ 243 ],
   alphaCSR[ 0 ][ 244 ],
   alphaCSR[ 0 ][ 245 ],
   alphaCSR[ 0 ][ 246 ],
   alphaCSR[ 0 ][ 247 ],
   alphaCSR[ 0 ][ 248 ],
   alphaCSR[ 0 ][ 249 ],
   alphaCSR[ 0 ][ 250 ],
   alphaCSR[ 0 ][ 251 ],
   alphaCSR[ 0 ][ 252 ],
   alphaCSR[ 0 ][ 253 ],
   alphaCSR[ 0 ][ 254 ],
   alphaCSR[ 0 ][ 255 ],
   alphaCSR[ 0 ][ 256 ],
   alphaCSR[ 0 ][ 257 ],
   alphaCSR[ 0 ][ 258 ],
   alphaCSR[ 0 ][ 259 ],
   alphaCSR[ 0 ][ 260 ],
   alphaCSR[ 0 ][ 261 ],
   alphaCSR[ 0 ][ 262 ],
   alphaCSR[ 0 ][ 263 ],
   alphaCSR[ 0 ][ 264 ],
   alphaCSR[ 0 ][ 265 ],
   alphaCSR[ 0 ][ 266 ],
   alphaCSR[ 0 ][ 267 ],
   alphaCSR[ 0 ][ 268 ],
   alphaCSR[ 0 ][ 269 ],
   alphaCSR[ 0 ][ 270 ],
   alphaCSR[ 0 ][ 271 ],
   alphaCSR[ 0 ][ 272 ],
   alphaCSR[ 0 ][ 273 ],
   alphaCSR[ 0 ][ 274 ],
   alphaCSR[ 0 ][ 275 ],
   alphaCSR[ 0 ][ 276 ],
   alphaCSR[ 0 ][ 277 ],
   alphaCSR[ 0 ][ 278 ],
   alphaCSR[ 0 ][ 279 ],
   alphaCSR[ 0 ][ 280 ],
   alphaCSR[ 0 ][ 281 ],
   alphaCSR[ 0 ][ 282 ],
   alphaCSR[ 0 ][ 283 ],
   alphaCSR[ 0 ][ 284 ],
   alphaCSR[ 0 ][ 285 ],
   alphaCSR[ 0 ][ 286 ],
   alphaCSR[ 0 ][ 287 ],
   alphaCSR[ 0 ][ 288 ],
   alphaCSR[ 0 ][ 289 ],
   alphaCSR[ 0 ][ 290 ],
   alphaCSR[ 0 ][ 291 ],
   alphaCSR[ 0 ][ 292 ],
   alphaCSR[ 0 ][ 293 ],
   alphaCSR[ 0 ][ 294 ],
   alphaCSR[ 0 ][ 295 ],
   alphaCSR[ 0 ][ 296 ],
   alphaCSR[ 0 ][ 297 ],
   alphaCSR[ 0 ][ 298 ],
   alphaCSR[ 0 ][ 299 ],
   alphaCSR[ 0 ][ 300 ],
   alphaCSR[ 0 ][ 301 ],
   alphaCSR[ 0 ][ 302 ],
   alphaCSR[ 0 ][ 303 ],
   alphaCSR[ 0 ][ 304 ],
   alphaCSR[ 0 ][ 305 ],
   alphaCSR[ 0 ][ 306 ],
   alphaCSR[ 0 ][ 307 ],
   alphaCSR[ 0 ][ 308 ],
   alphaCSR[ 0 ][ 309 ],
   alphaCSR[ 0 ][ 310 ],
   alphaCSR[ 0 ][ 311 ],
   alphaCSR[ 0 ][ 312 ],
   alphaCSR[ 0 ][ 313 ],
   alphaCSR[ 0 ][ 314 ],
   alphaCSR[ 0 ][ 315 ],
   alphaCSR[ 0 ][ 316 ],
   alphaCSR[ 0 ][ 317 ],
   alphaCSR[ 0 ][ 318 ],
   alphaCSR[ 0 ][ 319 ],
   alphaCSR[ 0 ][ 320 ],
   alphaCSR[ 0 ][ 321 ],
   alphaCSR[ 0 ][ 322 ],
   alphaCSR[ 0 ][ 323 ],
   alphaCSR[ 0 ][ 324 ],
   alphaCSR[ 0 ][ 325 ],
   alphaCSR[ 0 ][ 326 ],
   alphaCSR[ 0 ][ 327 ],
   alphaCSR[ 0 ][ 328 ],
   alphaCSR[ 0 ][ 329 ],
   alphaCSR[ 0 ][ 330 ],
   alphaCSR[ 0 ][ 331 ],
   alphaCSR[ 0 ][ 332 ],
   alphaCSR[ 0 ][ 333 ],
   alphaCSR[ 0 ][ 334 ],
   alphaCSR[ 0 ][ 335 ],
   alphaCSR[ 0 ][ 336 ],
   alphaCSR[ 0 ][ 337 ],
   alphaCSR[ 0 ][ 338 ],
   alphaCSR[ 0 ][ 339 ],
   alphaCSR[ 0 ][ 340 ],
   alphaCSR[ 0 ][ 341 ],
   alphaCSR[ 0 ][ 342 ],
   alphaCSR[ 0 ][ 343 ],
   alphaCSR[ 0 ][ 344 ],
   alphaCSR[ 0 ][ 345 ],
   alphaCSR[ 0 ][ 346 ],
   alphaCSR[ 0 ][ 347 ],
   alphaCSR[ 0 ][ 348 ],
   alphaCSR[ 0 ][ 349 ],
   alphaCSR[ 0 ][ 350 ],
   alphaCSR[ 0 ][ 351 ],
   alphaCSR[ 0 ][ 352 ],
   alphaCSR[ 0 ][ 353 ],
   alphaCSR[ 0 ][ 354 ],
   alphaCSR[ 0 ][ 355 ],
   alphaCSR[ 0 ][ 356 ],
   alphaCSR[ 0 ][ 357 ],
   alphaCSR[ 0 ][ 358 ],
   alphaCSR[ 0 ][ 359 ],
   alphaCSR[ 0 ][ 360 ],
   alphaCSR[ 0 ][ 361 ],
   alphaCSR[ 0 ][ 362 ],
   alphaCSR[ 0 ][ 363 ],
   alphaCSR[ 0 ][ 364 ],
   alphaCSR[ 0 ][ 365 ],
   alphaCSR[ 0 ][ 366 ],
   alphaCSR[ 0 ][ 367 ],
   alphaCSR[ 0 ][ 368 ],
   alphaCSR[ 0 ][ 369 ],
   alphaCSR[ 0 ][ 370 ],
   alphaCSR[ 0 ][ 371 ],
   alphaCSR[ 0 ][ 372 ],
   alphaCSR[ 0 ][ 373 ],
   alphaCSR[ 0 ][ 374 ],
   alphaCSR[ 0 ][ 375 ],
   alphaCSR[ 0 ][ 376 ],
   alphaCSR[ 0 ][ 377 ],
   alphaCSR[ 0 ][ 378 ],
   alphaCSR[ 0 ][ 379 ],
   alphaCSR[ 0 ][ 380 ],
   alphaCSR[ 0 ][ 381 ],
   alphaCSR[ 0 ][ 382 ],
   alphaCSR[ 0 ][ 383 ],
   alphaCSR[ 1 ][ 0 ],
   alphaCSR[ 1 ][ 1 ],
   alphaCSR[ 1 ][ 2 ],
   alphaCSR[ 1 ][ 3 ],
   alphaCSR[ 1 ][ 4 ],
   alphaCSR[ 1 ][ 5 ],
   alphaCSR[ 1 ][ 6 ],
   alphaCSR[ 1 ][ 7 ],
   alphaCSR[ 1 ][ 8 ],
   alphaCSR[ 1 ][ 9 ],
   alphaCSR[ 1 ][ 10 ],
   alphaCSR[ 1 ][ 11 ],
   alphaCSR[ 1 ][ 12 ],
   alphaCSR[ 1 ][ 13 ],
   alphaCSR[ 1 ][ 14 ],
   alphaCSR[ 1 ][ 15 ],
   alphaCSR[ 1 ][ 16 ],
   alphaCSR[ 1 ][ 17 ],
   alphaCSR[ 1 ][ 18 ],
   alphaCSR[ 1 ][ 19 ],
   alphaCSR[ 1 ][ 20 ],
   alphaCSR[ 1 ][ 21 ],
   alphaCSR[ 1 ][ 22 ],
   alphaCSR[ 1 ][ 23 ],
   alphaCSR[ 1 ][ 24 ],
   alphaCSR[ 1 ][ 25 ],
   alphaCSR[ 1 ][ 26 ],
   alphaCSR[ 1 ][ 27 ],
   alphaCSR[ 1 ][ 28 ],
   alphaCSR[ 1 ][ 29 ],
   alphaCSR[ 1 ][ 30 ],
   alphaCSR[ 1 ][ 31 ],
   alphaCSR[ 1 ][ 32 ],
   alphaCSR[ 1 ][ 33 ],
   alphaCSR[ 1 ][ 34 ],
   alphaCSR[ 1 ][ 35 ],
   alphaCSR[ 1 ][ 36 ],
   alphaCSR[ 1 ][ 37 ],
   alphaCSR[ 1 ][ 38 ],
   alphaCSR[ 1 ][ 39 ],
   alphaCSR[ 1 ][ 40 ],
   alphaCSR[ 1 ][ 41 ],
   alphaCSR[ 1 ][ 42 ],
   alphaCSR[ 1 ][ 43 ],
   alphaCSR[ 1 ][ 44 ],
   alphaCSR[ 1 ][ 45 ],
   alphaCSR[ 1 ][ 46 ],
   alphaCSR[ 1 ][ 47 ],
   alphaCSR[ 1 ][ 48 ],
   alphaCSR[ 1 ][ 49 ],
   alphaCSR[ 1 ][ 50 ],
   alphaCSR[ 1 ][ 51 ],
   alphaCSR[ 1 ][ 52 ],
   alphaCSR[ 1 ][ 53 ],
   alphaCSR[ 1 ][ 54 ],
   alphaCSR[ 1 ][ 55 ],
   alphaCSR[ 1 ][ 56 ],
   alphaCSR[ 1 ][ 57 ],
   alphaCSR[ 1 ][ 58 ],
   alphaCSR[ 1 ][ 59 ],
   alphaCSR[ 1 ][ 60 ],
   alphaCSR[ 1 ][ 61 ],
   alphaCSR[ 1 ][ 62 ],
   alphaCSR[ 1 ][ 63 ],
   alphaCSR[ 1 ][ 64 ],
   alphaCSR[ 1 ][ 65 ],
   alphaCSR[ 1 ][ 66 ],
   alphaCSR[ 1 ][ 67 ],
   alphaCSR[ 1 ][ 68 ],
   alphaCSR[ 1 ][ 69 ],
   alphaCSR[ 1 ][ 70 ],
   alphaCSR[ 1 ][ 71 ],
   alphaCSR[ 1 ][ 72 ],
   alphaCSR[ 1 ][ 73 ],
   alphaCSR[ 1 ][ 74 ],
   alphaCSR[ 1 ][ 75 ],
   alphaCSR[ 1 ][ 76 ],
   alphaCSR[ 1 ][ 77 ],
   alphaCSR[ 1 ][ 78 ],
   alphaCSR[ 1 ][ 79 ],
   alphaCSR[ 1 ][ 80 ],
   alphaCSR[ 1 ][ 81 ],
   alphaCSR[ 1 ][ 82 ],
   alphaCSR[ 1 ][ 83 ],
   alphaCSR[ 1 ][ 84 ],
   alphaCSR[ 1 ][ 85 ],
   alphaCSR[ 1 ][ 86 ],
   alphaCSR[ 1 ][ 87 ],
   alphaCSR[ 1 ][ 88 ],
   alphaCSR[ 1 ][ 89 ],
   alphaCSR[ 1 ][ 90 ],
   alphaCSR[ 1 ][ 91 ],
   alphaCSR[ 1 ][ 92 ],
   alphaCSR[ 1 ][ 93 ],
   alphaCSR[ 1 ][ 94 ],
   alphaCSR[ 1 ][ 95 ],
   alphaCSR[ 1 ][ 96 ],
   alphaCSR[ 1 ][ 97 ],
   alphaCSR[ 1 ][ 98 ],
   alphaCSR[ 1 ][ 99 ],
   alphaCSR[ 1 ][ 100 ],
   alphaCSR[ 1 ][ 101 ],
   alphaCSR[ 1 ][ 102 ],
   alphaCSR[ 1 ][ 103 ],
   alphaCSR[ 1 ][ 104 ],
   alphaCSR[ 1 ][ 105 ],
   alphaCSR[ 1 ][ 106 ],
   alphaCSR[ 1 ][ 107 ],
   alphaCSR[ 1 ][ 108 ],
   alphaCSR[ 1 ][ 109 ],
   alphaCSR[ 1 ][ 110 ],
   alphaCSR[ 1 ][ 111 ],
   alphaCSR[ 1 ][ 112 ],
   alphaCSR[ 1 ][ 113 ],
   alphaCSR[ 1 ][ 114 ],
   alphaCSR[ 1 ][ 115 ],
   alphaCSR[ 1 ][ 116 ],
   alphaCSR[ 1 ][ 117 ],
   alphaCSR[ 1 ][ 118 ],
   alphaCSR[ 1 ][ 119 ],
   alphaCSR[ 1 ][ 120 ],
   alphaCSR[ 1 ][ 121 ],
   alphaCSR[ 1 ][ 122 ],
   alphaCSR[ 1 ][ 123 ],
   alphaCSR[ 1 ][ 124 ],
   alphaCSR[ 1 ][ 125 ],
   alphaCSR[ 1 ][ 126 ],
   alphaCSR[ 1 ][ 127 ],
   alphaCSR[ 1 ][ 128 ],
   alphaCSR[ 1 ][ 129 ],
   alphaCSR[ 1 ][ 130 ],
   alphaCSR[ 1 ][ 131 ],
   alphaCSR[ 1 ][ 132 ],
   alphaCSR[ 1 ][ 133 ],
   alphaCSR[ 1 ][ 134 ],
   alphaCSR[ 1 ][ 135 ],
   alphaCSR[ 1 ][ 136 ],
   alphaCSR[ 1 ][ 137 ],
   alphaCSR[ 1 ][ 138 ],
   alphaCSR[ 1 ][ 139 ],
   alphaCSR[ 1 ][ 140 ],
   alphaCSR[ 1 ][ 141 ],
   alphaCSR[ 1 ][ 142 ],
   alphaCSR[ 1 ][ 143 ],
   alphaCSR[ 1 ][ 144 ],
   alphaCSR[ 1 ][ 145 ],
   alphaCSR[ 1 ][ 146 ],
   alphaCSR[ 1 ][ 147 ],
   alphaCSR[ 1 ][ 148 ],
   alphaCSR[ 1 ][ 149 ],
   alphaCSR[ 1 ][ 150 ],
   alphaCSR[ 1 ][ 151 ],
   alphaCSR[ 1 ][ 152 ],
   alphaCSR[ 1 ][ 153 ],
   alphaCSR[ 1 ][ 154 ],
   alphaCSR[ 1 ][ 155 ],
   alphaCSR[ 1 ][ 156 ],
   alphaCSR[ 1 ][ 157 ],
   alphaCSR[ 1 ][ 158 ],
   alphaCSR[ 1 ][ 159 ],
   alphaCSR[ 1 ][ 160 ],
   alphaCSR[ 1 ][ 161 ],
   alphaCSR[ 1 ][ 162 ],
   alphaCSR[ 1 ][ 163 ],
   alphaCSR[ 1 ][ 164 ],
   alphaCSR[ 1 ][ 165 ],
   alphaCSR[ 1 ][ 166 ],
   alphaCSR[ 1 ][ 167 ],
   alphaCSR[ 1 ][ 168 ],
   alphaCSR[ 1 ][ 169 ],
   alphaCSR[ 1 ][ 170 ],
   alphaCSR[ 1 ][ 171 ],
   alphaCSR[ 1 ][ 172 ],
   alphaCSR[ 1 ][ 173 ],
   alphaCSR[ 1 ][ 174 ],
   alphaCSR[ 1 ][ 175 ],
   alphaCSR[ 1 ][ 176 ],
   alphaCSR[ 1 ][ 177 ],
   alphaCSR[ 1 ][ 178 ],
   alphaCSR[ 1 ][ 179 ],
   alphaCSR[ 1 ][ 180 ],
   alphaCSR[ 1 ][ 181 ],
   alphaCSR[ 1 ][ 182 ],
   alphaCSR[ 1 ][ 183 ],
   alphaCSR[ 1 ][ 184 ],
   alphaCSR[ 1 ][ 185 ],
   alphaCSR[ 1 ][ 186 ],
   alphaCSR[ 1 ][ 187 ],
   alphaCSR[ 1 ][ 188 ],
   alphaCSR[ 1 ][ 189 ],
   alphaCSR[ 1 ][ 190 ],
   alphaCSR[ 1 ][ 191 ],
   alphaCSR[ 1 ][ 192 ],
   alphaCSR[ 1 ][ 193 ],
   alphaCSR[ 1 ][ 194 ],
   alphaCSR[ 1 ][ 195 ],
   alphaCSR[ 1 ][ 196 ],
   alphaCSR[ 1 ][ 197 ],
   alphaCSR[ 1 ][ 198 ],
   alphaCSR[ 1 ][ 199 ],
   alphaCSR[ 1 ][ 200 ],
   alphaCSR[ 1 ][ 201 ],
   alphaCSR[ 1 ][ 202 ],
   alphaCSR[ 1 ][ 203 ],
   alphaCSR[ 1 ][ 204 ],
   alphaCSR[ 1 ][ 205 ],
   alphaCSR[ 1 ][ 206 ],
   alphaCSR[ 1 ][ 207 ],
   alphaCSR[ 1 ][ 208 ],
   alphaCSR[ 1 ][ 209 ],
   alphaCSR[ 1 ][ 210 ],
   alphaCSR[ 1 ][ 211 ],
   alphaCSR[ 1 ][ 212 ],
   alphaCSR[ 1 ][ 213 ],
   alphaCSR[ 1 ][ 214 ],
   alphaCSR[ 1 ][ 215 ],
   alphaCSR[ 1 ][ 216 ],
   alphaCSR[ 1 ][ 217 ],
   alphaCSR[ 1 ][ 218 ],
   alphaCSR[ 1 ][ 219 ],
   alphaCSR[ 1 ][ 220 ],
   alphaCSR[ 1 ][ 221 ],
   alphaCSR[ 1 ][ 222 ],
   alphaCSR[ 1 ][ 223 ],
   alphaCSR[ 1 ][ 224 ],
   alphaCSR[ 1 ][ 225 ],
   alphaCSR[ 1 ][ 226 ],
   alphaCSR[ 1 ][ 227 ],
   alphaCSR[ 1 ][ 228 ],
   alphaCSR[ 1 ][ 229 ],
   alphaCSR[ 1 ][ 230 ],
   alphaCSR[ 1 ][ 231 ],
   alphaCSR[ 1 ][ 232 ],
   alphaCSR[ 1 ][ 233 ],
   alphaCSR[ 1 ][ 234 ],
   alphaCSR[ 1 ][ 235 ],
   alphaCSR[ 1 ][ 236 ],
   alphaCSR[ 1 ][ 237 ],
   alphaCSR[ 1 ][ 238 ],
   alphaCSR[ 1 ][ 239 ],
   alphaCSR[ 1 ][ 240 ],
   alphaCSR[ 1 ][ 241 ],
   alphaCSR[ 1 ][ 242 ],
   alphaCSR[ 1 ][ 243 ],
   alphaCSR[ 1 ][ 244 ],
   alphaCSR[ 1 ][ 245 ],
   alphaCSR[ 1 ][ 246 ],
   alphaCSR[ 1 ][ 247 ],
   alphaCSR[ 1 ][ 248 ],
   alphaCSR[ 1 ][ 249 ],
   alphaCSR[ 1 ][ 250 ],
   alphaCSR[ 1 ][ 251 ],
   alphaCSR[ 1 ][ 252 ],
   alphaCSR[ 1 ][ 253 ],
   alphaCSR[ 1 ][ 254 ],
   alphaCSR[ 1 ][ 255 ],
   alphaCSR[ 1 ][ 256 ],
   alphaCSR[ 1 ][ 257 ],
   alphaCSR[ 1 ][ 258 ],
   alphaCSR[ 1 ][ 259 ],
   alphaCSR[ 1 ][ 260 ],
   alphaCSR[ 1 ][ 261 ],
   alphaCSR[ 1 ][ 262 ],
   alphaCSR[ 1 ][ 263 ],
   alphaCSR[ 1 ][ 264 ],
   alphaCSR[ 1 ][ 265 ],
   alphaCSR[ 1 ][ 266 ],
   alphaCSR[ 1 ][ 267 ],
   alphaCSR[ 1 ][ 268 ],
   alphaCSR[ 1 ][ 269 ],
   alphaCSR[ 1 ][ 270 ],
   alphaCSR[ 1 ][ 271 ],
   alphaCSR[ 1 ][ 272 ],
   alphaCSR[ 1 ][ 273 ],
   alphaCSR[ 1 ][ 274 ],
   alphaCSR[ 1 ][ 275 ],
   alphaCSR[ 1 ][ 276 ],
   alphaCSR[ 1 ][ 277 ],
   alphaCSR[ 1 ][ 278 ],
   alphaCSR[ 1 ][ 279 ],
   alphaCSR[ 1 ][ 280 ],
   alphaCSR[ 1 ][ 281 ],
   alphaCSR[ 1 ][ 282 ],
   alphaCSR[ 1 ][ 283 ],
   alphaCSR[ 1 ][ 284 ],
   alphaCSR[ 1 ][ 285 ],
   alphaCSR[ 1 ][ 286 ],
   alphaCSR[ 1 ][ 287 ],
   alphaCSR[ 1 ][ 288 ],
   alphaCSR[ 1 ][ 289 ],
   alphaCSR[ 1 ][ 290 ],
   alphaCSR[ 1 ][ 291 ],
   alphaCSR[ 1 ][ 292 ],
   alphaCSR[ 1 ][ 293 ],
   alphaCSR[ 1 ][ 294 ],
   alphaCSR[ 1 ][ 295 ],
   alphaCSR[ 1 ][ 296 ],
   alphaCSR[ 1 ][ 297 ],
   alphaCSR[ 1 ][ 298 ],
   alphaCSR[ 1 ][ 299 ],
   alphaCSR[ 1 ][ 300 ],
   alphaCSR[ 1 ][ 301 ],
   alphaCSR[ 1 ][ 302 ],
   alphaCSR[ 1 ][ 303 ],
   alphaCSR[ 1 ][ 304 ],
   alphaCSR[ 1 ][ 305 ],
   alphaCSR[ 1 ][ 306 ],
   alphaCSR[ 1 ][ 307 ],
   alphaCSR[ 1 ][ 308 ],
   alphaCSR[ 1 ][ 309 ],
   alphaCSR[ 1 ][ 310 ],
   alphaCSR[ 1 ][ 311 ],
   alphaCSR[ 1 ][ 312 ],
   alphaCSR[ 1 ][ 313 ],
   alphaCSR[ 1 ][ 314 ],
   alphaCSR[ 1 ][ 315 ],
   alphaCSR[ 1 ][ 316 ],
   alphaCSR[ 1 ][ 317 ],
   alphaCSR[ 1 ][ 318 ],
   alphaCSR[ 1 ][ 319 ],
   alphaCSR[ 1 ][ 320 ],
   alphaCSR[ 1 ][ 321 ],
   alphaCSR[ 1 ][ 322 ],
   alphaCSR[ 1 ][ 323 ],
   alphaCSR[ 1 ][ 324 ],
   alphaCSR[ 1 ][ 325 ],
   alphaCSR[ 1 ][ 326 ],
   alphaCSR[ 1 ][ 327 ],
   alphaCSR[ 1 ][ 328 ],
   alphaCSR[ 1 ][ 329 ],
   alphaCSR[ 1 ][ 330 ],
   alphaCSR[ 1 ][ 331 ],
   alphaCSR[ 1 ][ 332 ],
   alphaCSR[ 1 ][ 333 ],
   alphaCSR[ 1 ][ 334 ],
   alphaCSR[ 1 ][ 335 ],
   alphaCSR[ 1 ][ 336 ],
   alphaCSR[ 1 ][ 337 ],
   alphaCSR[ 1 ][ 338 ],
   alphaCSR[ 1 ][ 339 ],
   alphaCSR[ 1 ][ 340 ],
   alphaCSR[ 1 ][ 341 ],
   alphaCSR[ 1 ][ 342 ],
   alphaCSR[ 1 ][ 343 ],
   alphaCSR[ 1 ][ 344 ],
   alphaCSR[ 1 ][ 345 ],
   alphaCSR[ 1 ][ 346 ],
   alphaCSR[ 1 ][ 347 ],
   alphaCSR[ 1 ][ 348 ],
   alphaCSR[ 1 ][ 349 ],
   alphaCSR[ 1 ][ 350 ],
   alphaCSR[ 1 ][ 351 ],
   alphaCSR[ 1 ][ 352 ],
   alphaCSR[ 1 ][ 353 ],
   alphaCSR[ 1 ][ 354 ],
   alphaCSR[ 1 ][ 355 ],
   alphaCSR[ 1 ][ 356 ],
   alphaCSR[ 1 ][ 357 ],
   alphaCSR[ 1 ][ 358 ],
   alphaCSR[ 1 ][ 359 ],
   alphaCSR[ 1 ][ 360 ],
   alphaCSR[ 1 ][ 361 ],
   alphaCSR[ 1 ][ 362 ],
   alphaCSR[ 1 ][ 363 ],
   alphaCSR[ 1 ][ 364 ],
   alphaCSR[ 1 ][ 365 ],
   alphaCSR[ 1 ][ 366 ],
   alphaCSR[ 1 ][ 367 ],
   alphaCSR[ 1 ][ 368 ],
   alphaCSR[ 1 ][ 369 ],
   alphaCSR[ 1 ][ 370 ],
   alphaCSR[ 1 ][ 371 ],
   alphaCSR[ 1 ][ 372 ],
   alphaCSR[ 1 ][ 373 ],
   alphaCSR[ 1 ][ 374 ],
   alphaCSR[ 1 ][ 375 ],
   alphaCSR[ 1 ][ 376 ],
   alphaCSR[ 1 ][ 377 ],
   alphaCSR[ 1 ][ 378 ],
   alphaCSR[ 1 ][ 379 ],
   alphaCSR[ 1 ][ 380 ],
   alphaCSR[ 1 ][ 381 ],
   alphaCSR[ 1 ][ 382 ],
   alphaCSR[ 1 ][ 383 ],
   alphaCSR[ 2 ][ 0 ],
   alphaCSR[ 2 ][ 1 ],
   alphaCSR[ 2 ][ 2 ],
   alphaCSR[ 2 ][ 3 ],
   alphaCSR[ 2 ][ 4 ],
   alphaCSR[ 2 ][ 5 ],
   alphaCSR[ 2 ][ 6 ],
   alphaCSR[ 2 ][ 7 ],
   alphaCSR[ 2 ][ 8 ],
   alphaCSR[ 2 ][ 9 ],
   alphaCSR[ 2 ][ 10 ],
   alphaCSR[ 2 ][ 11 ],
   alphaCSR[ 2 ][ 12 ],
   alphaCSR[ 2 ][ 13 ],
   alphaCSR[ 2 ][ 14 ],
   alphaCSR[ 2 ][ 15 ],
   alphaCSR[ 2 ][ 16 ],
   alphaCSR[ 2 ][ 17 ],
   alphaCSR[ 2 ][ 18 ],
   alphaCSR[ 2 ][ 19 ],
   alphaCSR[ 2 ][ 20 ],
   alphaCSR[ 2 ][ 21 ],
   alphaCSR[ 2 ][ 22 ],
   alphaCSR[ 2 ][ 23 ],
   alphaCSR[ 2 ][ 24 ],
   alphaCSR[ 2 ][ 25 ],
   alphaCSR[ 2 ][ 26 ],
   alphaCSR[ 2 ][ 27 ],
   alphaCSR[ 2 ][ 28 ],
   alphaCSR[ 2 ][ 29 ],
   alphaCSR[ 2 ][ 30 ],
   alphaCSR[ 2 ][ 31 ],
   alphaCSR[ 2 ][ 32 ],
   alphaCSR[ 2 ][ 33 ],
   alphaCSR[ 2 ][ 34 ],
   alphaCSR[ 2 ][ 35 ],
   alphaCSR[ 2 ][ 36 ],
   alphaCSR[ 2 ][ 37 ],
   alphaCSR[ 2 ][ 38 ],
   alphaCSR[ 2 ][ 39 ],
   alphaCSR[ 2 ][ 40 ],
   alphaCSR[ 2 ][ 41 ],
   alphaCSR[ 2 ][ 42 ],
   alphaCSR[ 2 ][ 43 ],
   alphaCSR[ 2 ][ 44 ],
   alphaCSR[ 2 ][ 45 ],
   alphaCSR[ 2 ][ 46 ],
   alphaCSR[ 2 ][ 47 ],
   alphaCSR[ 2 ][ 48 ],
   alphaCSR[ 2 ][ 49 ],
   alphaCSR[ 2 ][ 50 ],
   alphaCSR[ 2 ][ 51 ],
   alphaCSR[ 2 ][ 52 ],
   alphaCSR[ 2 ][ 53 ],
   alphaCSR[ 2 ][ 54 ],
   alphaCSR[ 2 ][ 55 ],
   alphaCSR[ 2 ][ 56 ],
   alphaCSR[ 2 ][ 57 ],
   alphaCSR[ 2 ][ 58 ],
   alphaCSR[ 2 ][ 59 ],
   alphaCSR[ 2 ][ 60 ],
   alphaCSR[ 2 ][ 61 ],
   alphaCSR[ 2 ][ 62 ],
   alphaCSR[ 2 ][ 63 ],
   alphaCSR[ 2 ][ 64 ],
   alphaCSR[ 2 ][ 65 ],
   alphaCSR[ 2 ][ 66 ],
   alphaCSR[ 2 ][ 67 ],
   alphaCSR[ 2 ][ 68 ],
   alphaCSR[ 2 ][ 69 ],
   alphaCSR[ 2 ][ 70 ],
   alphaCSR[ 2 ][ 71 ],
   alphaCSR[ 2 ][ 72 ],
   alphaCSR[ 2 ][ 73 ],
   alphaCSR[ 2 ][ 74 ],
   alphaCSR[ 2 ][ 75 ],
   alphaCSR[ 2 ][ 76 ],
   alphaCSR[ 2 ][ 77 ],
   alphaCSR[ 2 ][ 78 ],
   alphaCSR[ 2 ][ 79 ],
   alphaCSR[ 2 ][ 80 ],
   alphaCSR[ 2 ][ 81 ],
   alphaCSR[ 2 ][ 82 ],
   alphaCSR[ 2 ][ 83 ],
   alphaCSR[ 2 ][ 84 ],
   alphaCSR[ 2 ][ 85 ],
   alphaCSR[ 2 ][ 86 ],
   alphaCSR[ 2 ][ 87 ],
   alphaCSR[ 2 ][ 88 ],
   alphaCSR[ 2 ][ 89 ],
   alphaCSR[ 2 ][ 90 ],
   alphaCSR[ 2 ][ 91 ],
   alphaCSR[ 2 ][ 92 ],
   alphaCSR[ 2 ][ 93 ],
   alphaCSR[ 2 ][ 94 ],
   alphaCSR[ 2 ][ 95 ],
   alphaCSR[ 2 ][ 96 ],
   alphaCSR[ 2 ][ 97 ],
   alphaCSR[ 2 ][ 98 ],
   alphaCSR[ 2 ][ 99 ],
   alphaCSR[ 2 ][ 100 ],
   alphaCSR[ 2 ][ 101 ],
   alphaCSR[ 2 ][ 102 ],
   alphaCSR[ 2 ][ 103 ],
   alphaCSR[ 2 ][ 104 ],
   alphaCSR[ 2 ][ 105 ],
   alphaCSR[ 2 ][ 106 ],
   alphaCSR[ 2 ][ 107 ],
   alphaCSR[ 2 ][ 108 ],
   alphaCSR[ 2 ][ 109 ],
   alphaCSR[ 2 ][ 110 ],
   alphaCSR[ 2 ][ 111 ],
   alphaCSR[ 2 ][ 112 ],
   alphaCSR[ 2 ][ 113 ],
   alphaCSR[ 2 ][ 114 ],
   alphaCSR[ 2 ][ 115 ],
   alphaCSR[ 2 ][ 116 ],
   alphaCSR[ 2 ][ 117 ],
   alphaCSR[ 2 ][ 118 ],
   alphaCSR[ 2 ][ 119 ],
   alphaCSR[ 2 ][ 120 ],
   alphaCSR[ 2 ][ 121 ],
   alphaCSR[ 2 ][ 122 ],
   alphaCSR[ 2 ][ 123 ],
   alphaCSR[ 2 ][ 124 ],
   alphaCSR[ 2 ][ 125 ],
   alphaCSR[ 2 ][ 126 ],
   alphaCSR[ 2 ][ 127 ],
   alphaCSR[ 2 ][ 128 ],
   alphaCSR[ 2 ][ 129 ],
   alphaCSR[ 2 ][ 130 ],
   alphaCSR[ 2 ][ 131 ],
   alphaCSR[ 2 ][ 132 ],
   alphaCSR[ 2 ][ 133 ],
   alphaCSR[ 2 ][ 134 ],
   alphaCSR[ 2 ][ 135 ],
   alphaCSR[ 2 ][ 136 ],
   alphaCSR[ 2 ][ 137 ],
   alphaCSR[ 2 ][ 138 ],
   alphaCSR[ 2 ][ 139 ],
   alphaCSR[ 2 ][ 140 ],
   alphaCSR[ 2 ][ 141 ],
   alphaCSR[ 2 ][ 142 ],
   alphaCSR[ 2 ][ 143 ],
   alphaCSR[ 2 ][ 144 ],
   alphaCSR[ 2 ][ 145 ],
   alphaCSR[ 2 ][ 146 ],
   alphaCSR[ 2 ][ 147 ],
   alphaCSR[ 2 ][ 148 ],
   alphaCSR[ 2 ][ 149 ],
   alphaCSR[ 2 ][ 150 ],
   alphaCSR[ 2 ][ 151 ],
   alphaCSR[ 2 ][ 152 ],
   alphaCSR[ 2 ][ 153 ],
   alphaCSR[ 2 ][ 154 ],
   alphaCSR[ 2 ][ 155 ],
   alphaCSR[ 2 ][ 156 ],
   alphaCSR[ 2 ][ 157 ],
   alphaCSR[ 2 ][ 158 ],
   alphaCSR[ 2 ][ 159 ],
   alphaCSR[ 2 ][ 160 ],
   alphaCSR[ 2 ][ 161 ],
   alphaCSR[ 2 ][ 162 ],
   alphaCSR[ 2 ][ 163 ],
   alphaCSR[ 2 ][ 164 ],
   alphaCSR[ 2 ][ 165 ],
   alphaCSR[ 2 ][ 166 ],
   alphaCSR[ 2 ][ 167 ],
   alphaCSR[ 2 ][ 168 ],
   alphaCSR[ 2 ][ 169 ],
   alphaCSR[ 2 ][ 170 ],
   alphaCSR[ 2 ][ 171 ],
   alphaCSR[ 2 ][ 172 ],
   alphaCSR[ 2 ][ 173 ],
   alphaCSR[ 2 ][ 174 ],
   alphaCSR[ 2 ][ 175 ],
   alphaCSR[ 2 ][ 176 ],
   alphaCSR[ 2 ][ 177 ],
   alphaCSR[ 2 ][ 178 ],
   alphaCSR[ 2 ][ 179 ],
   alphaCSR[ 2 ][ 180 ],
   alphaCSR[ 2 ][ 181 ],
   alphaCSR[ 2 ][ 182 ],
   alphaCSR[ 2 ][ 183 ],
   alphaCSR[ 2 ][ 184 ],
   alphaCSR[ 2 ][ 185 ],
   alphaCSR[ 2 ][ 186 ],
   alphaCSR[ 2 ][ 187 ],
   alphaCSR[ 2 ][ 188 ],
   alphaCSR[ 2 ][ 189 ],
   alphaCSR[ 2 ][ 190 ],
   alphaCSR[ 2 ][ 191 ],
   alphaCSR[ 2 ][ 192 ],
   alphaCSR[ 2 ][ 193 ],
   alphaCSR[ 2 ][ 194 ],
   alphaCSR[ 2 ][ 195 ],
   alphaCSR[ 2 ][ 196 ],
   alphaCSR[ 2 ][ 197 ],
   alphaCSR[ 2 ][ 198 ],
   alphaCSR[ 2 ][ 199 ],
   alphaCSR[ 2 ][ 200 ],
   alphaCSR[ 2 ][ 201 ],
   alphaCSR[ 2 ][ 202 ],
   alphaCSR[ 2 ][ 203 ],
   alphaCSR[ 2 ][ 204 ],
   alphaCSR[ 2 ][ 205 ],
   alphaCSR[ 2 ][ 206 ],
   alphaCSR[ 2 ][ 207 ],
   alphaCSR[ 2 ][ 208 ],
   alphaCSR[ 2 ][ 209 ],
   alphaCSR[ 2 ][ 210 ],
   alphaCSR[ 2 ][ 211 ],
   alphaCSR[ 2 ][ 212 ],
   alphaCSR[ 2 ][ 213 ],
   alphaCSR[ 2 ][ 214 ],
   alphaCSR[ 2 ][ 215 ],
   alphaCSR[ 2 ][ 216 ],
   alphaCSR[ 2 ][ 217 ],
   alphaCSR[ 2 ][ 218 ],
   alphaCSR[ 2 ][ 219 ],
   alphaCSR[ 2 ][ 220 ],
   alphaCSR[ 2 ][ 221 ],
   alphaCSR[ 2 ][ 222 ],
   alphaCSR[ 2 ][ 223 ],
   alphaCSR[ 2 ][ 224 ],
   alphaCSR[ 2 ][ 225 ],
   alphaCSR[ 2 ][ 226 ],
   alphaCSR[ 2 ][ 227 ],
   alphaCSR[ 2 ][ 228 ],
   alphaCSR[ 2 ][ 229 ],
   alphaCSR[ 2 ][ 230 ],
   alphaCSR[ 2 ][ 231 ],
   alphaCSR[ 2 ][ 232 ],
   alphaCSR[ 2 ][ 233 ],
   alphaCSR[ 2 ][ 234 ],
   alphaCSR[ 2 ][ 235 ],
   alphaCSR[ 2 ][ 236 ],
   alphaCSR[ 2 ][ 237 ],
   alphaCSR[ 2 ][ 238 ],
   alphaCSR[ 2 ][ 239 ],
   alphaCSR[ 2 ][ 240 ],
   alphaCSR[ 2 ][ 241 ],
   alphaCSR[ 2 ][ 242 ],
   alphaCSR[ 2 ][ 243 ],
   alphaCSR[ 2 ][ 244 ],
   alphaCSR[ 2 ][ 245 ],
   alphaCSR[ 2 ][ 246 ],
   alphaCSR[ 2 ][ 247 ],
   alphaCSR[ 2 ][ 248 ],
   alphaCSR[ 2 ][ 249 ],
   alphaCSR[ 2 ][ 250 ],
   alphaCSR[ 2 ][ 251 ],
   alphaCSR[ 2 ][ 252 ],
   alphaCSR[ 2 ][ 253 ],
   alphaCSR[ 2 ][ 254 ],
   alphaCSR[ 2 ][ 255 ],
   alphaCSR[ 2 ][ 256 ],
   alphaCSR[ 2 ][ 257 ],
   alphaCSR[ 2 ][ 258 ],
   alphaCSR[ 2 ][ 259 ],
   alphaCSR[ 2 ][ 260 ],
   alphaCSR[ 2 ][ 261 ],
   alphaCSR[ 2 ][ 262 ],
   alphaCSR[ 2 ][ 263 ],
   alphaCSR[ 2 ][ 264 ],
   alphaCSR[ 2 ][ 265 ],
   alphaCSR[ 2 ][ 266 ],
   alphaCSR[ 2 ][ 267 ],
   alphaCSR[ 2 ][ 268 ],
   alphaCSR[ 2 ][ 269 ],
   alphaCSR[ 2 ][ 270 ],
   alphaCSR[ 2 ][ 271 ],
   alphaCSR[ 2 ][ 272 ],
   alphaCSR[ 2 ][ 273 ],
   alphaCSR[ 2 ][ 274 ],
   alphaCSR[ 2 ][ 275 ],
   alphaCSR[ 2 ][ 276 ],
   alphaCSR[ 2 ][ 277 ],
   alphaCSR[ 2 ][ 278 ],
   alphaCSR[ 2 ][ 279 ],
   alphaCSR[ 2 ][ 280 ],
   alphaCSR[ 2 ][ 281 ],
   alphaCSR[ 2 ][ 282 ],
   alphaCSR[ 2 ][ 283 ],
   alphaCSR[ 2 ][ 284 ],
   alphaCSR[ 2 ][ 285 ],
   alphaCSR[ 2 ][ 286 ],
   alphaCSR[ 2 ][ 287 ],
   alphaCSR[ 2 ][ 288 ],
   alphaCSR[ 2 ][ 289 ],
   alphaCSR[ 2 ][ 290 ],
   alphaCSR[ 2 ][ 291 ],
   alphaCSR[ 2 ][ 292 ],
   alphaCSR[ 2 ][ 293 ],
   alphaCSR[ 2 ][ 294 ],
   alphaCSR[ 2 ][ 295 ],
   alphaCSR[ 2 ][ 296 ],
   alphaCSR[ 2 ][ 297 ],
   alphaCSR[ 2 ][ 298 ],
   alphaCSR[ 2 ][ 299 ],
   alphaCSR[ 2 ][ 300 ],
   alphaCSR[ 2 ][ 301 ],
   alphaCSR[ 2 ][ 302 ],
   alphaCSR[ 2 ][ 303 ],
   alphaCSR[ 2 ][ 304 ],
   alphaCSR[ 2 ][ 305 ],
   alphaCSR[ 2 ][ 306 ],
   alphaCSR[ 2 ][ 307 ],
   alphaCSR[ 2 ][ 308 ],
   alphaCSR[ 2 ][ 309 ],
   alphaCSR[ 2 ][ 310 ],
   alphaCSR[ 2 ][ 311 ],
   alphaCSR[ 2 ][ 312 ],
   alphaCSR[ 2 ][ 313 ],
   alphaCSR[ 2 ][ 314 ],
   alphaCSR[ 2 ][ 315 ],
   alphaCSR[ 2 ][ 316 ],
   alphaCSR[ 2 ][ 317 ],
   alphaCSR[ 2 ][ 318 ],
   alphaCSR[ 2 ][ 319 ],
   alphaCSR[ 2 ][ 320 ],
   alphaCSR[ 2 ][ 321 ],
   alphaCSR[ 2 ][ 322 ],
   alphaCSR[ 2 ][ 323 ],
   alphaCSR[ 2 ][ 324 ],
   alphaCSR[ 2 ][ 325 ],
   alphaCSR[ 2 ][ 326 ],
   alphaCSR[ 2 ][ 327 ],
   alphaCSR[ 2 ][ 328 ],
   alphaCSR[ 2 ][ 329 ],
   alphaCSR[ 2 ][ 330 ],
   alphaCSR[ 2 ][ 331 ],
   alphaCSR[ 2 ][ 332 ],
   alphaCSR[ 2 ][ 333 ],
   alphaCSR[ 2 ][ 334 ],
   alphaCSR[ 2 ][ 335 ],
   alphaCSR[ 2 ][ 336 ],
   alphaCSR[ 2 ][ 337 ],
   alphaCSR[ 2 ][ 338 ],
   alphaCSR[ 2 ][ 339 ],
   alphaCSR[ 2 ][ 340 ],
   alphaCSR[ 2 ][ 341 ],
   alphaCSR[ 2 ][ 342 ],
   alphaCSR[ 2 ][ 343 ],
   alphaCSR[ 2 ][ 344 ],
   alphaCSR[ 2 ][ 345 ],
   alphaCSR[ 2 ][ 346 ],
   alphaCSR[ 2 ][ 347 ],
   alphaCSR[ 2 ][ 348 ],
   alphaCSR[ 2 ][ 349 ],
   alphaCSR[ 2 ][ 350 ],
   alphaCSR[ 2 ][ 351 ],
   alphaCSR[ 2 ][ 352 ],
   alphaCSR[ 2 ][ 353 ],
   alphaCSR[ 2 ][ 354 ],
   alphaCSR[ 2 ][ 355 ],
   alphaCSR[ 2 ][ 356 ],
   alphaCSR[ 2 ][ 357 ],
   alphaCSR[ 2 ][ 358 ],
   alphaCSR[ 2 ][ 359 ],
   alphaCSR[ 2 ][ 360 ],
   alphaCSR[ 2 ][ 361 ],
   alphaCSR[ 2 ][ 362 ],
   alphaCSR[ 2 ][ 363 ],
   alphaCSR[ 2 ][ 364 ],
   alphaCSR[ 2 ][ 365 ],
   alphaCSR[ 2 ][ 366 ],
   alphaCSR[ 2 ][ 367 ],
   alphaCSR[ 2 ][ 368 ],
   alphaCSR[ 2 ][ 369 ],
   alphaCSR[ 2 ][ 370 ],
   alphaCSR[ 2 ][ 371 ],
   alphaCSR[ 2 ][ 372 ],
   alphaCSR[ 2 ][ 373 ],
   alphaCSR[ 2 ][ 374 ],
   alphaCSR[ 2 ][ 375 ],
   alphaCSR[ 2 ][ 376 ],
   alphaCSR[ 2 ][ 377 ],
   alphaCSR[ 2 ][ 378 ],
   alphaCSR[ 2 ][ 379 ],
   alphaCSR[ 2 ][ 380 ],
   alphaCSR[ 2 ][ 381 ],
   alphaCSR[ 2 ][ 382 ],
   alphaCSR[ 2 ][ 383 ],
   alphaCSR[ 3 ][ 0 ],
   alphaCSR[ 3 ][ 1 ],
   alphaCSR[ 3 ][ 2 ],
   alphaCSR[ 3 ][ 3 ],
   alphaCSR[ 3 ][ 4 ],
   alphaCSR[ 3 ][ 5 ],
   alphaCSR[ 3 ][ 6 ],
   alphaCSR[ 3 ][ 7 ],
   alphaCSR[ 3 ][ 8 ],
   alphaCSR[ 3 ][ 9 ],
   alphaCSR[ 3 ][ 10 ],
   alphaCSR[ 3 ][ 11 ],
   alphaCSR[ 3 ][ 12 ],
   alphaCSR[ 3 ][ 13 ],
   alphaCSR[ 3 ][ 14 ],
   alphaCSR[ 3 ][ 15 ],
   alphaCSR[ 3 ][ 16 ],
   alphaCSR[ 3 ][ 17 ],
   alphaCSR[ 3 ][ 18 ],
   alphaCSR[ 3 ][ 19 ],
   alphaCSR[ 3 ][ 20 ],
   alphaCSR[ 3 ][ 21 ],
   alphaCSR[ 3 ][ 22 ],
   alphaCSR[ 3 ][ 23 ],
   alphaCSR[ 3 ][ 24 ],
   alphaCSR[ 3 ][ 25 ],
   alphaCSR[ 3 ][ 26 ],
   alphaCSR[ 3 ][ 27 ],
   alphaCSR[ 3 ][ 28 ],
   alphaCSR[ 3 ][ 29 ],
   alphaCSR[ 3 ][ 30 ],
   alphaCSR[ 3 ][ 31 ],
   alphaCSR[ 3 ][ 32 ],
   alphaCSR[ 3 ][ 33 ],
   alphaCSR[ 3 ][ 34 ],
   alphaCSR[ 3 ][ 35 ],
   alphaCSR[ 3 ][ 36 ],
   alphaCSR[ 3 ][ 37 ],
   alphaCSR[ 3 ][ 38 ],
   alphaCSR[ 3 ][ 39 ],
   alphaCSR[ 3 ][ 40 ],
   alphaCSR[ 3 ][ 41 ],
   alphaCSR[ 3 ][ 42 ],
   alphaCSR[ 3 ][ 43 ],
   alphaCSR[ 3 ][ 44 ],
   alphaCSR[ 3 ][ 45 ],
   alphaCSR[ 3 ][ 46 ],
   alphaCSR[ 3 ][ 47 ],
   alphaCSR[ 3 ][ 48 ],
   alphaCSR[ 3 ][ 49 ],
   alphaCSR[ 3 ][ 50 ],
   alphaCSR[ 3 ][ 51 ],
   alphaCSR[ 3 ][ 52 ],
   alphaCSR[ 3 ][ 53 ],
   alphaCSR[ 3 ][ 54 ],
   alphaCSR[ 3 ][ 55 ],
   alphaCSR[ 3 ][ 56 ],
   alphaCSR[ 3 ][ 57 ],
   alphaCSR[ 3 ][ 58 ],
   alphaCSR[ 3 ][ 59 ],
   alphaCSR[ 3 ][ 60 ],
   alphaCSR[ 3 ][ 61 ],
   alphaCSR[ 3 ][ 62 ],
   alphaCSR[ 3 ][ 63 ],
   alphaCSR[ 3 ][ 64 ],
   alphaCSR[ 3 ][ 65 ],
   alphaCSR[ 3 ][ 66 ],
   alphaCSR[ 3 ][ 67 ],
   alphaCSR[ 3 ][ 68 ],
   alphaCSR[ 3 ][ 69 ],
   alphaCSR[ 3 ][ 70 ],
   alphaCSR[ 3 ][ 71 ],
   alphaCSR[ 3 ][ 72 ],
   alphaCSR[ 3 ][ 73 ],
   alphaCSR[ 3 ][ 74 ],
   alphaCSR[ 3 ][ 75 ],
   alphaCSR[ 3 ][ 76 ],
   alphaCSR[ 3 ][ 77 ],
   alphaCSR[ 3 ][ 78 ],
   alphaCSR[ 3 ][ 79 ],
   alphaCSR[ 3 ][ 80 ],
   alphaCSR[ 3 ][ 81 ],
   alphaCSR[ 3 ][ 82 ],
   alphaCSR[ 3 ][ 83 ],
   alphaCSR[ 3 ][ 84 ],
   alphaCSR[ 3 ][ 85 ],
   alphaCSR[ 3 ][ 86 ],
   alphaCSR[ 3 ][ 87 ],
   alphaCSR[ 3 ][ 88 ],
   alphaCSR[ 3 ][ 89 ],
   alphaCSR[ 3 ][ 90 ],
   alphaCSR[ 3 ][ 91 ],
   alphaCSR[ 3 ][ 92 ],
   alphaCSR[ 3 ][ 93 ],
   alphaCSR[ 3 ][ 94 ],
   alphaCSR[ 3 ][ 95 ],
   alphaCSR[ 3 ][ 96 ],
   alphaCSR[ 3 ][ 97 ],
   alphaCSR[ 3 ][ 98 ],
   alphaCSR[ 3 ][ 99 ],
   alphaCSR[ 3 ][ 100 ],
   alphaCSR[ 3 ][ 101 ],
   alphaCSR[ 3 ][ 102 ],
   alphaCSR[ 3 ][ 103 ],
   alphaCSR[ 3 ][ 104 ],
   alphaCSR[ 3 ][ 105 ],
   alphaCSR[ 3 ][ 106 ],
   alphaCSR[ 3 ][ 107 ],
   alphaCSR[ 3 ][ 108 ],
   alphaCSR[ 3 ][ 109 ],
   alphaCSR[ 3 ][ 110 ],
   alphaCSR[ 3 ][ 111 ],
   alphaCSR[ 3 ][ 112 ],
   alphaCSR[ 3 ][ 113 ],
   alphaCSR[ 3 ][ 114 ],
   alphaCSR[ 3 ][ 115 ],
   alphaCSR[ 3 ][ 116 ],
   alphaCSR[ 3 ][ 117 ],
   alphaCSR[ 3 ][ 118 ],
   alphaCSR[ 3 ][ 119 ],
   alphaCSR[ 3 ][ 120 ],
   alphaCSR[ 3 ][ 121 ],
   alphaCSR[ 3 ][ 122 ],
   alphaCSR[ 3 ][ 123 ],
   alphaCSR[ 3 ][ 124 ],
   alphaCSR[ 3 ][ 125 ],
   alphaCSR[ 3 ][ 126 ],
   alphaCSR[ 3 ][ 127 ],
   alphaCSR[ 3 ][ 128 ],
   alphaCSR[ 3 ][ 129 ],
   alphaCSR[ 3 ][ 130 ],
   alphaCSR[ 3 ][ 131 ],
   alphaCSR[ 3 ][ 132 ],
   alphaCSR[ 3 ][ 133 ],
   alphaCSR[ 3 ][ 134 ],
   alphaCSR[ 3 ][ 135 ],
   alphaCSR[ 3 ][ 136 ],
   alphaCSR[ 3 ][ 137 ],
   alphaCSR[ 3 ][ 138 ],
   alphaCSR[ 3 ][ 139 ],
   alphaCSR[ 3 ][ 140 ],
   alphaCSR[ 3 ][ 141 ],
   alphaCSR[ 3 ][ 142 ],
   alphaCSR[ 3 ][ 143 ],
   alphaCSR[ 3 ][ 144 ],
   alphaCSR[ 3 ][ 145 ],
   alphaCSR[ 3 ][ 146 ],
   alphaCSR[ 3 ][ 147 ],
   alphaCSR[ 3 ][ 148 ],
   alphaCSR[ 3 ][ 149 ],
   alphaCSR[ 3 ][ 150 ],
   alphaCSR[ 3 ][ 151 ],
   alphaCSR[ 3 ][ 152 ],
   alphaCSR[ 3 ][ 153 ],
   alphaCSR[ 3 ][ 154 ],
   alphaCSR[ 3 ][ 155 ],
   alphaCSR[ 3 ][ 156 ],
   alphaCSR[ 3 ][ 157 ],
   alphaCSR[ 3 ][ 158 ],
   alphaCSR[ 3 ][ 159 ],
   alphaCSR[ 3 ][ 160 ],
   alphaCSR[ 3 ][ 161 ],
   alphaCSR[ 3 ][ 162 ],
   alphaCSR[ 3 ][ 163 ],
   alphaCSR[ 3 ][ 164 ],
   alphaCSR[ 3 ][ 165 ],
   alphaCSR[ 3 ][ 166 ],
   alphaCSR[ 3 ][ 167 ],
   alphaCSR[ 3 ][ 168 ],
   alphaCSR[ 3 ][ 169 ],
   alphaCSR[ 3 ][ 170 ],
   alphaCSR[ 3 ][ 171 ],
   alphaCSR[ 3 ][ 172 ],
   alphaCSR[ 3 ][ 173 ],
   alphaCSR[ 3 ][ 174 ],
   alphaCSR[ 3 ][ 175 ],
   alphaCSR[ 3 ][ 176 ],
   alphaCSR[ 3 ][ 177 ],
   alphaCSR[ 3 ][ 178 ],
   alphaCSR[ 3 ][ 179 ],
   alphaCSR[ 3 ][ 180 ],
   alphaCSR[ 3 ][ 181 ],
   alphaCSR[ 3 ][ 182 ],
   alphaCSR[ 3 ][ 183 ],
   alphaCSR[ 3 ][ 184 ],
   alphaCSR[ 3 ][ 185 ],
   alphaCSR[ 3 ][ 186 ],
   alphaCSR[ 3 ][ 187 ],
   alphaCSR[ 3 ][ 188 ],
   alphaCSR[ 3 ][ 189 ],
   alphaCSR[ 3 ][ 190 ],
   alphaCSR[ 3 ][ 191 ],
   alphaCSR[ 3 ][ 192 ],
   alphaCSR[ 3 ][ 193 ],
   alphaCSR[ 3 ][ 194 ],
   alphaCSR[ 3 ][ 195 ],
   alphaCSR[ 3 ][ 196 ],
   alphaCSR[ 3 ][ 197 ],
   alphaCSR[ 3 ][ 198 ],
   alphaCSR[ 3 ][ 199 ],
   alphaCSR[ 3 ][ 200 ],
   alphaCSR[ 3 ][ 201 ],
   alphaCSR[ 3 ][ 202 ],
   alphaCSR[ 3 ][ 203 ],
   alphaCSR[ 3 ][ 204 ],
   alphaCSR[ 3 ][ 205 ],
   alphaCSR[ 3 ][ 206 ],
   alphaCSR[ 3 ][ 207 ],
   alphaCSR[ 3 ][ 208 ],
   alphaCSR[ 3 ][ 209 ],
   alphaCSR[ 3 ][ 210 ],
   alphaCSR[ 3 ][ 211 ],
   alphaCSR[ 3 ][ 212 ],
   alphaCSR[ 3 ][ 213 ],
   alphaCSR[ 3 ][ 214 ],
   alphaCSR[ 3 ][ 215 ],
   alphaCSR[ 3 ][ 216 ],
   alphaCSR[ 3 ][ 217 ],
   alphaCSR[ 3 ][ 218 ],
   alphaCSR[ 3 ][ 219 ],
   alphaCSR[ 3 ][ 220 ],
   alphaCSR[ 3 ][ 221 ],
   alphaCSR[ 3 ][ 222 ],
   alphaCSR[ 3 ][ 223 ],
   alphaCSR[ 3 ][ 224 ],
   alphaCSR[ 3 ][ 225 ],
   alphaCSR[ 3 ][ 226 ],
   alphaCSR[ 3 ][ 227 ],
   alphaCSR[ 3 ][ 228 ],
   alphaCSR[ 3 ][ 229 ],
   alphaCSR[ 3 ][ 230 ],
   alphaCSR[ 3 ][ 231 ],
   alphaCSR[ 3 ][ 232 ],
   alphaCSR[ 3 ][ 233 ],
   alphaCSR[ 3 ][ 234 ],
   alphaCSR[ 3 ][ 235 ],
   alphaCSR[ 3 ][ 236 ],
   alphaCSR[ 3 ][ 237 ],
   alphaCSR[ 3 ][ 238 ],
   alphaCSR[ 3 ][ 239 ],
   alphaCSR[ 3 ][ 240 ],
   alphaCSR[ 3 ][ 241 ],
   alphaCSR[ 3 ][ 242 ],
   alphaCSR[ 3 ][ 243 ],
   alphaCSR[ 3 ][ 244 ],
   alphaCSR[ 3 ][ 245 ],
   alphaCSR[ 3 ][ 246 ],
   alphaCSR[ 3 ][ 247 ],
   alphaCSR[ 3 ][ 248 ],
   alphaCSR[ 3 ][ 249 ],
   alphaCSR[ 3 ][ 250 ],
   alphaCSR[ 3 ][ 251 ],
   alphaCSR[ 3 ][ 252 ],
   alphaCSR[ 3 ][ 253 ],
   alphaCSR[ 3 ][ 254 ],
   alphaCSR[ 3 ][ 255 ],
   alphaCSR[ 3 ][ 256 ],
   alphaCSR[ 3 ][ 257 ],
   alphaCSR[ 3 ][ 258 ],
   alphaCSR[ 3 ][ 259 ],
   alphaCSR[ 3 ][ 260 ],
   alphaCSR[ 3 ][ 261 ],
   alphaCSR[ 3 ][ 262 ],
   alphaCSR[ 3 ][ 263 ],
   alphaCSR[ 3 ][ 264 ],
   alphaCSR[ 3 ][ 265 ],
   alphaCSR[ 3 ][ 266 ],
   alphaCSR[ 3 ][ 267 ],
   alphaCSR[ 3 ][ 268 ],
   alphaCSR[ 3 ][ 269 ],
   alphaCSR[ 3 ][ 270 ],
   alphaCSR[ 3 ][ 271 ],
   alphaCSR[ 3 ][ 272 ],
   alphaCSR[ 3 ][ 273 ],
   alphaCSR[ 3 ][ 274 ],
   alphaCSR[ 3 ][ 275 ],
   alphaCSR[ 3 ][ 276 ],
   alphaCSR[ 3 ][ 277 ],
   alphaCSR[ 3 ][ 278 ],
   alphaCSR[ 3 ][ 279 ],
   alphaCSR[ 3 ][ 280 ],
   alphaCSR[ 3 ][ 281 ],
   alphaCSR[ 3 ][ 282 ],
   alphaCSR[ 3 ][ 283 ],
   alphaCSR[ 3 ][ 284 ],
   alphaCSR[ 3 ][ 285 ],
   alphaCSR[ 3 ][ 286 ],
   alphaCSR[ 3 ][ 287 ],
   alphaCSR[ 3 ][ 288 ],
   alphaCSR[ 3 ][ 289 ],
   alphaCSR[ 3 ][ 290 ],
   alphaCSR[ 3 ][ 291 ],
   alphaCSR[ 3 ][ 292 ],
   alphaCSR[ 3 ][ 293 ],
   alphaCSR[ 3 ][ 294 ],
   alphaCSR[ 3 ][ 295 ],
   alphaCSR[ 3 ][ 296 ],
   alphaCSR[ 3 ][ 297 ],
   alphaCSR[ 3 ][ 298 ],
   alphaCSR[ 3 ][ 299 ],
   alphaCSR[ 3 ][ 300 ],
   alphaCSR[ 3 ][ 301 ],
   alphaCSR[ 3 ][ 302 ],
   alphaCSR[ 3 ][ 303 ],
   alphaCSR[ 3 ][ 304 ],
   alphaCSR[ 3 ][ 305 ],
   alphaCSR[ 3 ][ 306 ],
   alphaCSR[ 3 ][ 307 ],
   alphaCSR[ 3 ][ 308 ],
   alphaCSR[ 3 ][ 309 ],
   alphaCSR[ 3 ][ 310 ],
   alphaCSR[ 3 ][ 311 ],
   alphaCSR[ 3 ][ 312 ],
   alphaCSR[ 3 ][ 313 ],
   alphaCSR[ 3 ][ 314 ],
   alphaCSR[ 3 ][ 315 ],
   alphaCSR[ 3 ][ 316 ],
   alphaCSR[ 3 ][ 317 ],
   alphaCSR[ 3 ][ 318 ],
   alphaCSR[ 3 ][ 319 ],
   alphaCSR[ 3 ][ 320 ],
   alphaCSR[ 3 ][ 321 ],
   alphaCSR[ 3 ][ 322 ],
   alphaCSR[ 3 ][ 323 ],
   alphaCSR[ 3 ][ 324 ],
   alphaCSR[ 3 ][ 325 ],
   alphaCSR[ 3 ][ 326 ],
   alphaCSR[ 3 ][ 327 ],
   alphaCSR[ 3 ][ 328 ],
   alphaCSR[ 3 ][ 329 ],
   alphaCSR[ 3 ][ 330 ],
   alphaCSR[ 3 ][ 331 ],
   alphaCSR[ 3 ][ 332 ],
   alphaCSR[ 3 ][ 333 ],
   alphaCSR[ 3 ][ 334 ],
   alphaCSR[ 3 ][ 335 ],
   alphaCSR[ 3 ][ 336 ],
   alphaCSR[ 3 ][ 337 ],
   alphaCSR[ 3 ][ 338 ],
   alphaCSR[ 3 ][ 339 ],
   alphaCSR[ 3 ][ 340 ],
   alphaCSR[ 3 ][ 341 ],
   alphaCSR[ 3 ][ 342 ],
   alphaCSR[ 3 ][ 343 ],
   alphaCSR[ 3 ][ 344 ],
   alphaCSR[ 3 ][ 345 ],
   alphaCSR[ 3 ][ 346 ],
   alphaCSR[ 3 ][ 347 ],
   alphaCSR[ 3 ][ 348 ],
   alphaCSR[ 3 ][ 349 ],
   alphaCSR[ 3 ][ 350 ],
   alphaCSR[ 3 ][ 351 ],
   alphaCSR[ 3 ][ 352 ],
   alphaCSR[ 3 ][ 353 ],
   alphaCSR[ 3 ][ 354 ],
   alphaCSR[ 3 ][ 355 ],
   alphaCSR[ 3 ][ 356 ],
   alphaCSR[ 3 ][ 357 ],
   alphaCSR[ 3 ][ 358 ],
   alphaCSR[ 3 ][ 359 ],
   alphaCSR[ 3 ][ 360 ],
   alphaCSR[ 3 ][ 361 ],
   alphaCSR[ 3 ][ 362 ],
   alphaCSR[ 3 ][ 363 ],
   alphaCSR[ 3 ][ 364 ],
   alphaCSR[ 3 ][ 365 ],
   alphaCSR[ 3 ][ 366 ],
   alphaCSR[ 3 ][ 367 ],
   alphaCSR[ 3 ][ 368 ],
   alphaCSR[ 3 ][ 369 ],
   alphaCSR[ 3 ][ 370 ],
   alphaCSR[ 3 ][ 371 ],
   alphaCSR[ 3 ][ 372 ],
   alphaCSR[ 3 ][ 373 ],
   alphaCSR[ 3 ][ 374 ],
   alphaCSR[ 3 ][ 375 ],
   alphaCSR[ 3 ][ 376 ],
   alphaCSR[ 3 ][ 377 ],
   alphaCSR[ 3 ][ 378 ],
   alphaCSR[ 3 ][ 379 ],
   alphaCSR[ 3 ][ 380 ],
   alphaCSR[ 3 ][ 381 ],
   alphaCSR[ 3 ][ 382 ],
   alphaCSR[ 3 ][ 383 ],
   alphaCSR[ 4 ][ 0 ],
   alphaCSR[ 4 ][ 1 ],
   alphaCSR[ 4 ][ 2 ],
   alphaCSR[ 4 ][ 3 ],
   alphaCSR[ 4 ][ 4 ],
   alphaCSR[ 4 ][ 5 ],
   alphaCSR[ 4 ][ 6 ],
   alphaCSR[ 4 ][ 7 ],
   alphaCSR[ 4 ][ 8 ],
   alphaCSR[ 4 ][ 9 ],
   alphaCSR[ 4 ][ 10 ],
   alphaCSR[ 4 ][ 11 ],
   alphaCSR[ 4 ][ 12 ],
   alphaCSR[ 4 ][ 13 ],
   alphaCSR[ 4 ][ 14 ],
   alphaCSR[ 4 ][ 15 ],
   alphaCSR[ 4 ][ 16 ],
   alphaCSR[ 4 ][ 17 ],
   alphaCSR[ 4 ][ 18 ],
   alphaCSR[ 4 ][ 19 ],
   alphaCSR[ 4 ][ 20 ],
   alphaCSR[ 4 ][ 21 ],
   alphaCSR[ 4 ][ 22 ],
   alphaCSR[ 4 ][ 23 ],
   alphaCSR[ 4 ][ 24 ],
   alphaCSR[ 4 ][ 25 ],
   alphaCSR[ 4 ][ 26 ],
   alphaCSR[ 4 ][ 27 ],
   alphaCSR[ 4 ][ 28 ],
   alphaCSR[ 4 ][ 29 ],
   alphaCSR[ 4 ][ 30 ],
   alphaCSR[ 4 ][ 31 ],
   alphaCSR[ 4 ][ 32 ],
   alphaCSR[ 4 ][ 33 ],
   alphaCSR[ 4 ][ 34 ],
   alphaCSR[ 4 ][ 35 ],
   alphaCSR[ 4 ][ 36 ],
   alphaCSR[ 4 ][ 37 ],
   alphaCSR[ 4 ][ 38 ],
   alphaCSR[ 4 ][ 39 ],
   alphaCSR[ 4 ][ 40 ],
   alphaCSR[ 4 ][ 41 ],
   alphaCSR[ 4 ][ 42 ],
   alphaCSR[ 4 ][ 43 ],
   alphaCSR[ 4 ][ 44 ],
   alphaCSR[ 4 ][ 45 ],
   alphaCSR[ 4 ][ 46 ],
   alphaCSR[ 4 ][ 47 ],
   alphaCSR[ 4 ][ 48 ],
   alphaCSR[ 4 ][ 49 ],
   alphaCSR[ 4 ][ 50 ],
   alphaCSR[ 4 ][ 51 ],
   alphaCSR[ 4 ][ 52 ],
   alphaCSR[ 4 ][ 53 ],
   alphaCSR[ 4 ][ 54 ],
   alphaCSR[ 4 ][ 55 ],
   alphaCSR[ 4 ][ 56 ],
   alphaCSR[ 4 ][ 57 ],
   alphaCSR[ 4 ][ 58 ],
   alphaCSR[ 4 ][ 59 ],
   alphaCSR[ 4 ][ 60 ],
   alphaCSR[ 4 ][ 61 ],
   alphaCSR[ 4 ][ 62 ],
   alphaCSR[ 4 ][ 63 ],
   alphaCSR[ 4 ][ 64 ],
   alphaCSR[ 4 ][ 65 ],
   alphaCSR[ 4 ][ 66 ],
   alphaCSR[ 4 ][ 67 ],
   alphaCSR[ 4 ][ 68 ],
   alphaCSR[ 4 ][ 69 ],
   alphaCSR[ 4 ][ 70 ],
   alphaCSR[ 4 ][ 71 ],
   alphaCSR[ 4 ][ 72 ],
   alphaCSR[ 4 ][ 73 ],
   alphaCSR[ 4 ][ 74 ],
   alphaCSR[ 4 ][ 75 ],
   alphaCSR[ 4 ][ 76 ],
   alphaCSR[ 4 ][ 77 ],
   alphaCSR[ 4 ][ 78 ],
   alphaCSR[ 4 ][ 79 ],
   alphaCSR[ 4 ][ 80 ],
   alphaCSR[ 4 ][ 81 ],
   alphaCSR[ 4 ][ 82 ],
   alphaCSR[ 4 ][ 83 ],
   alphaCSR[ 4 ][ 84 ],
   alphaCSR[ 4 ][ 85 ],
   alphaCSR[ 4 ][ 86 ],
   alphaCSR[ 4 ][ 87 ],
   alphaCSR[ 4 ][ 88 ],
   alphaCSR[ 4 ][ 89 ],
   alphaCSR[ 4 ][ 90 ],
   alphaCSR[ 4 ][ 91 ],
   alphaCSR[ 4 ][ 92 ],
   alphaCSR[ 4 ][ 93 ],
   alphaCSR[ 4 ][ 94 ],
   alphaCSR[ 4 ][ 95 ],
   alphaCSR[ 4 ][ 96 ],
   alphaCSR[ 4 ][ 97 ],
   alphaCSR[ 4 ][ 98 ],
   alphaCSR[ 4 ][ 99 ],
   alphaCSR[ 4 ][ 100 ],
   alphaCSR[ 4 ][ 101 ],
   alphaCSR[ 4 ][ 102 ],
   alphaCSR[ 4 ][ 103 ],
   alphaCSR[ 4 ][ 104 ],
   alphaCSR[ 4 ][ 105 ],
   alphaCSR[ 4 ][ 106 ],
   alphaCSR[ 4 ][ 107 ],
   alphaCSR[ 4 ][ 108 ],
   alphaCSR[ 4 ][ 109 ],
   alphaCSR[ 4 ][ 110 ],
   alphaCSR[ 4 ][ 111 ],
   alphaCSR[ 4 ][ 112 ],
   alphaCSR[ 4 ][ 113 ],
   alphaCSR[ 4 ][ 114 ],
   alphaCSR[ 4 ][ 115 ],
   alphaCSR[ 4 ][ 116 ],
   alphaCSR[ 4 ][ 117 ],
   alphaCSR[ 4 ][ 118 ],
   alphaCSR[ 4 ][ 119 ],
   alphaCSR[ 4 ][ 120 ],
   alphaCSR[ 4 ][ 121 ],
   alphaCSR[ 4 ][ 122 ],
   alphaCSR[ 4 ][ 123 ],
   alphaCSR[ 4 ][ 124 ],
   alphaCSR[ 4 ][ 125 ],
   alphaCSR[ 4 ][ 126 ],
   alphaCSR[ 4 ][ 127 ],
   alphaCSR[ 4 ][ 128 ],
   alphaCSR[ 4 ][ 129 ],
   alphaCSR[ 4 ][ 130 ],
   alphaCSR[ 4 ][ 131 ],
   alphaCSR[ 4 ][ 132 ],
   alphaCSR[ 4 ][ 133 ],
   alphaCSR[ 4 ][ 134 ],
   alphaCSR[ 4 ][ 135 ],
   alphaCSR[ 4 ][ 136 ],
   alphaCSR[ 4 ][ 137 ],
   alphaCSR[ 4 ][ 138 ],
   alphaCSR[ 4 ][ 139 ],
   alphaCSR[ 4 ][ 140 ],
   alphaCSR[ 4 ][ 141 ],
   alphaCSR[ 4 ][ 142 ],
   alphaCSR[ 4 ][ 143 ],
   alphaCSR[ 4 ][ 144 ],
   alphaCSR[ 4 ][ 145 ],
   alphaCSR[ 4 ][ 146 ],
   alphaCSR[ 4 ][ 147 ],
   alphaCSR[ 4 ][ 148 ],
   alphaCSR[ 4 ][ 149 ],
   alphaCSR[ 4 ][ 150 ],
   alphaCSR[ 4 ][ 151 ],
   alphaCSR[ 4 ][ 152 ],
   alphaCSR[ 4 ][ 153 ],
   alphaCSR[ 4 ][ 154 ],
   alphaCSR[ 4 ][ 155 ],
   alphaCSR[ 4 ][ 156 ],
   alphaCSR[ 4 ][ 157 ],
   alphaCSR[ 4 ][ 158 ],
   alphaCSR[ 4 ][ 159 ],
   alphaCSR[ 4 ][ 160 ],
   alphaCSR[ 4 ][ 161 ],
   alphaCSR[ 4 ][ 162 ],
   alphaCSR[ 4 ][ 163 ],
   alphaCSR[ 4 ][ 164 ],
   alphaCSR[ 4 ][ 165 ],
   alphaCSR[ 4 ][ 166 ],
   alphaCSR[ 4 ][ 167 ],
   alphaCSR[ 4 ][ 168 ],
   alphaCSR[ 4 ][ 169 ],
   alphaCSR[ 4 ][ 170 ],
   alphaCSR[ 4 ][ 171 ],
   alphaCSR[ 4 ][ 172 ],
   alphaCSR[ 4 ][ 173 ],
   alphaCSR[ 4 ][ 174 ],
   alphaCSR[ 4 ][ 175 ],
   alphaCSR[ 4 ][ 176 ],
   alphaCSR[ 4 ][ 177 ],
   alphaCSR[ 4 ][ 178 ],
   alphaCSR[ 4 ][ 179 ],
   alphaCSR[ 4 ][ 180 ],
   alphaCSR[ 4 ][ 181 ],
   alphaCSR[ 4 ][ 182 ],
   alphaCSR[ 4 ][ 183 ],
   alphaCSR[ 4 ][ 184 ],
   alphaCSR[ 4 ][ 185 ],
   alphaCSR[ 4 ][ 186 ],
   alphaCSR[ 4 ][ 187 ],
   alphaCSR[ 4 ][ 188 ],
   alphaCSR[ 4 ][ 189 ],
   alphaCSR[ 4 ][ 190 ],
   alphaCSR[ 4 ][ 191 ],
   alphaCSR[ 4 ][ 192 ],
   alphaCSR[ 4 ][ 193 ],
   alphaCSR[ 4 ][ 194 ],
   alphaCSR[ 4 ][ 195 ],
   alphaCSR[ 4 ][ 196 ],
   alphaCSR[ 4 ][ 197 ],
   alphaCSR[ 4 ][ 198 ],
   alphaCSR[ 4 ][ 199 ],
   alphaCSR[ 4 ][ 200 ],
   alphaCSR[ 4 ][ 201 ],
   alphaCSR[ 4 ][ 202 ],
   alphaCSR[ 4 ][ 203 ],
   alphaCSR[ 4 ][ 204 ],
   alphaCSR[ 4 ][ 205 ],
   alphaCSR[ 4 ][ 206 ],
   alphaCSR[ 4 ][ 207 ],
   alphaCSR[ 4 ][ 208 ],
   alphaCSR[ 4 ][ 209 ],
   alphaCSR[ 4 ][ 210 ],
   alphaCSR[ 4 ][ 211 ],
   alphaCSR[ 4 ][ 212 ],
   alphaCSR[ 4 ][ 213 ],
   alphaCSR[ 4 ][ 214 ],
   alphaCSR[ 4 ][ 215 ],
   alphaCSR[ 4 ][ 216 ],
   alphaCSR[ 4 ][ 217 ],
   alphaCSR[ 4 ][ 218 ],
   alphaCSR[ 4 ][ 219 ],
   alphaCSR[ 4 ][ 220 ],
   alphaCSR[ 4 ][ 221 ],
   alphaCSR[ 4 ][ 222 ],
   alphaCSR[ 4 ][ 223 ],
   alphaCSR[ 4 ][ 224 ],
   alphaCSR[ 4 ][ 225 ],
   alphaCSR[ 4 ][ 226 ],
   alphaCSR[ 4 ][ 227 ],
   alphaCSR[ 4 ][ 228 ],
   alphaCSR[ 4 ][ 229 ],
   alphaCSR[ 4 ][ 230 ],
   alphaCSR[ 4 ][ 231 ],
   alphaCSR[ 4 ][ 232 ],
   alphaCSR[ 4 ][ 233 ],
   alphaCSR[ 4 ][ 234 ],
   alphaCSR[ 4 ][ 235 ],
   alphaCSR[ 4 ][ 236 ],
   alphaCSR[ 4 ][ 237 ],
   alphaCSR[ 4 ][ 238 ],
   alphaCSR[ 4 ][ 239 ],
   alphaCSR[ 4 ][ 240 ],
   alphaCSR[ 4 ][ 241 ],
   alphaCSR[ 4 ][ 242 ],
   alphaCSR[ 4 ][ 243 ],
   alphaCSR[ 4 ][ 244 ],
   alphaCSR[ 4 ][ 245 ],
   alphaCSR[ 4 ][ 246 ],
   alphaCSR[ 4 ][ 247 ],
   alphaCSR[ 4 ][ 248 ],
   alphaCSR[ 4 ][ 249 ],
   alphaCSR[ 4 ][ 250 ],
   alphaCSR[ 4 ][ 251 ],
   alphaCSR[ 4 ][ 252 ],
   alphaCSR[ 4 ][ 253 ],
   alphaCSR[ 4 ][ 254 ],
   alphaCSR[ 4 ][ 255 ],
   alphaCSR[ 4 ][ 256 ],
   alphaCSR[ 4 ][ 257 ],
   alphaCSR[ 4 ][ 258 ],
   alphaCSR[ 4 ][ 259 ],
   alphaCSR[ 4 ][ 260 ],
   alphaCSR[ 4 ][ 261 ],
   alphaCSR[ 4 ][ 262 ],
   alphaCSR[ 4 ][ 263 ],
   alphaCSR[ 4 ][ 264 ],
   alphaCSR[ 4 ][ 265 ],
   alphaCSR[ 4 ][ 266 ],
   alphaCSR[ 4 ][ 267 ],
   alphaCSR[ 4 ][ 268 ],
   alphaCSR[ 4 ][ 269 ],
   alphaCSR[ 4 ][ 270 ],
   alphaCSR[ 4 ][ 271 ],
   alphaCSR[ 4 ][ 272 ],
   alphaCSR[ 4 ][ 273 ],
   alphaCSR[ 4 ][ 274 ],
   alphaCSR[ 4 ][ 275 ],
   alphaCSR[ 4 ][ 276 ],
   alphaCSR[ 4 ][ 277 ],
   alphaCSR[ 4 ][ 278 ],
   alphaCSR[ 4 ][ 279 ],
   alphaCSR[ 4 ][ 280 ],
   alphaCSR[ 4 ][ 281 ],
   alphaCSR[ 4 ][ 282 ],
   alphaCSR[ 4 ][ 283 ],
   alphaCSR[ 4 ][ 284 ],
   alphaCSR[ 4 ][ 285 ],
   alphaCSR[ 4 ][ 286 ],
   alphaCSR[ 4 ][ 287 ],
   alphaCSR[ 4 ][ 288 ],
   alphaCSR[ 4 ][ 289 ],
   alphaCSR[ 4 ][ 290 ],
   alphaCSR[ 4 ][ 291 ],
   alphaCSR[ 4 ][ 292 ],
   alphaCSR[ 4 ][ 293 ],
   alphaCSR[ 4 ][ 294 ],
   alphaCSR[ 4 ][ 295 ],
   alphaCSR[ 4 ][ 296 ],
   alphaCSR[ 4 ][ 297 ],
   alphaCSR[ 4 ][ 298 ],
   alphaCSR[ 4 ][ 299 ],
   alphaCSR[ 4 ][ 300 ],
   alphaCSR[ 4 ][ 301 ],
   alphaCSR[ 4 ][ 302 ],
   alphaCSR[ 4 ][ 303 ],
   alphaCSR[ 4 ][ 304 ],
   alphaCSR[ 4 ][ 305 ],
   alphaCSR[ 4 ][ 306 ],
   alphaCSR[ 4 ][ 307 ],
   alphaCSR[ 4 ][ 308 ],
   alphaCSR[ 4 ][ 309 ],
   alphaCSR[ 4 ][ 310 ],
   alphaCSR[ 4 ][ 311 ],
   alphaCSR[ 4 ][ 312 ],
   alphaCSR[ 4 ][ 313 ],
   alphaCSR[ 4 ][ 314 ],
   alphaCSR[ 4 ][ 315 ],
   alphaCSR[ 4 ][ 316 ],
   alphaCSR[ 4 ][ 317 ],
   alphaCSR[ 4 ][ 318 ],
   alphaCSR[ 4 ][ 319 ],
   alphaCSR[ 4 ][ 320 ],
   alphaCSR[ 4 ][ 321 ],
   alphaCSR[ 4 ][ 322 ],
   alphaCSR[ 4 ][ 323 ],
   alphaCSR[ 4 ][ 324 ],
   alphaCSR[ 4 ][ 325 ],
   alphaCSR[ 4 ][ 326 ],
   alphaCSR[ 4 ][ 327 ],
   alphaCSR[ 4 ][ 328 ],
   alphaCSR[ 4 ][ 329 ],
   alphaCSR[ 4 ][ 330 ],
   alphaCSR[ 4 ][ 331 ],
   alphaCSR[ 4 ][ 332 ],
   alphaCSR[ 4 ][ 333 ],
   alphaCSR[ 4 ][ 334 ],
   alphaCSR[ 4 ][ 335 ],
   alphaCSR[ 4 ][ 336 ],
   alphaCSR[ 4 ][ 337 ],
   alphaCSR[ 4 ][ 338 ],
   alphaCSR[ 4 ][ 339 ],
   alphaCSR[ 4 ][ 340 ],
   alphaCSR[ 4 ][ 341 ],
   alphaCSR[ 4 ][ 342 ],
   alphaCSR[ 4 ][ 343 ],
   alphaCSR[ 4 ][ 344 ],
   alphaCSR[ 4 ][ 345 ],
   alphaCSR[ 4 ][ 346 ],
   alphaCSR[ 4 ][ 347 ],
   alphaCSR[ 4 ][ 348 ],
   alphaCSR[ 4 ][ 349 ],
   alphaCSR[ 4 ][ 350 ],
   alphaCSR[ 4 ][ 351 ],
   alphaCSR[ 4 ][ 352 ],
   alphaCSR[ 4 ][ 353 ],
   alphaCSR[ 4 ][ 354 ],
   alphaCSR[ 4 ][ 355 ],
   alphaCSR[ 4 ][ 356 ],
   alphaCSR[ 4 ][ 357 ],
   alphaCSR[ 4 ][ 358 ],
   alphaCSR[ 4 ][ 359 ],
   alphaCSR[ 4 ][ 360 ],
   alphaCSR[ 4 ][ 361 ],
   alphaCSR[ 4 ][ 362 ],
   alphaCSR[ 4 ][ 363 ],
   alphaCSR[ 4 ][ 364 ],
   alphaCSR[ 4 ][ 365 ],
   alphaCSR[ 4 ][ 366 ],
   alphaCSR[ 4 ][ 367 ],
   alphaCSR[ 4 ][ 368 ],
   alphaCSR[ 4 ][ 369 ],
   alphaCSR[ 4 ][ 370 ],
   alphaCSR[ 4 ][ 371 ],
   alphaCSR[ 4 ][ 372 ],
   alphaCSR[ 4 ][ 373 ],
   alphaCSR[ 4 ][ 374 ],
   alphaCSR[ 4 ][ 375 ],
   alphaCSR[ 4 ][ 376 ],
   alphaCSR[ 4 ][ 377 ],
   alphaCSR[ 4 ][ 378 ],
   alphaCSR[ 4 ][ 379 ],
   alphaCSR[ 4 ][ 380 ],
   alphaCSR[ 4 ][ 381 ],
   alphaCSR[ 4 ][ 382 ],
   alphaCSR[ 4 ][ 383 ],
   alphaCSR[ 5 ][ 0 ],
   alphaCSR[ 5 ][ 1 ],
   alphaCSR[ 5 ][ 2 ],
   alphaCSR[ 5 ][ 3 ],
   alphaCSR[ 5 ][ 4 ],
   alphaCSR[ 5 ][ 5 ],
   alphaCSR[ 5 ][ 6 ],
   alphaCSR[ 5 ][ 7 ],
   alphaCSR[ 5 ][ 8 ],
   alphaCSR[ 5 ][ 9 ],
   alphaCSR[ 5 ][ 10 ],
   alphaCSR[ 5 ][ 11 ],
   alphaCSR[ 5 ][ 12 ],
   alphaCSR[ 5 ][ 13 ],
   alphaCSR[ 5 ][ 14 ],
   alphaCSR[ 5 ][ 15 ],
   alphaCSR[ 5 ][ 16 ],
   alphaCSR[ 5 ][ 17 ],
   alphaCSR[ 5 ][ 18 ],
   alphaCSR[ 5 ][ 19 ],
   alphaCSR[ 5 ][ 20 ],
   alphaCSR[ 5 ][ 21 ],
   alphaCSR[ 5 ][ 22 ],
   alphaCSR[ 5 ][ 23 ],
   alphaCSR[ 5 ][ 24 ],
   alphaCSR[ 5 ][ 25 ],
   alphaCSR[ 5 ][ 26 ],
   alphaCSR[ 5 ][ 27 ],
   alphaCSR[ 5 ][ 28 ],
   alphaCSR[ 5 ][ 29 ],
   alphaCSR[ 5 ][ 30 ],
   alphaCSR[ 5 ][ 31 ],
   alphaCSR[ 5 ][ 32 ],
   alphaCSR[ 5 ][ 33 ],
   alphaCSR[ 5 ][ 34 ],
   alphaCSR[ 5 ][ 35 ],
   alphaCSR[ 5 ][ 36 ],
   alphaCSR[ 5 ][ 37 ],
   alphaCSR[ 5 ][ 38 ],
   alphaCSR[ 5 ][ 39 ],
   alphaCSR[ 5 ][ 40 ],
   alphaCSR[ 5 ][ 41 ],
   alphaCSR[ 5 ][ 42 ],
   alphaCSR[ 5 ][ 43 ],
   alphaCSR[ 5 ][ 44 ],
   alphaCSR[ 5 ][ 45 ],
   alphaCSR[ 5 ][ 46 ],
   alphaCSR[ 5 ][ 47 ],
   alphaCSR[ 5 ][ 48 ],
   alphaCSR[ 5 ][ 49 ],
   alphaCSR[ 5 ][ 50 ],
   alphaCSR[ 5 ][ 51 ],
   alphaCSR[ 5 ][ 52 ],
   alphaCSR[ 5 ][ 53 ],
   alphaCSR[ 5 ][ 54 ],
   alphaCSR[ 5 ][ 55 ],
   alphaCSR[ 5 ][ 56 ],
   alphaCSR[ 5 ][ 57 ],
   alphaCSR[ 5 ][ 58 ],
   alphaCSR[ 5 ][ 59 ],
   alphaCSR[ 5 ][ 60 ],
   alphaCSR[ 5 ][ 61 ],
   alphaCSR[ 5 ][ 62 ],
   alphaCSR[ 5 ][ 63 ],
   alphaCSR[ 5 ][ 64 ],
   alphaCSR[ 5 ][ 65 ],
   alphaCSR[ 5 ][ 66 ],
   alphaCSR[ 5 ][ 67 ],
   alphaCSR[ 5 ][ 68 ],
   alphaCSR[ 5 ][ 69 ],
   alphaCSR[ 5 ][ 70 ],
   alphaCSR[ 5 ][ 71 ],
   alphaCSR[ 5 ][ 72 ],
   alphaCSR[ 5 ][ 73 ],
   alphaCSR[ 5 ][ 74 ],
   alphaCSR[ 5 ][ 75 ],
   alphaCSR[ 5 ][ 76 ],
   alphaCSR[ 5 ][ 77 ],
   alphaCSR[ 5 ][ 78 ],
   alphaCSR[ 5 ][ 79 ],
   alphaCSR[ 5 ][ 80 ],
   alphaCSR[ 5 ][ 81 ],
   alphaCSR[ 5 ][ 82 ],
   alphaCSR[ 5 ][ 83 ],
   alphaCSR[ 5 ][ 84 ],
   alphaCSR[ 5 ][ 85 ],
   alphaCSR[ 5 ][ 86 ],
   alphaCSR[ 5 ][ 87 ],
   alphaCSR[ 5 ][ 88 ],
   alphaCSR[ 5 ][ 89 ],
   alphaCSR[ 5 ][ 90 ],
   alphaCSR[ 5 ][ 91 ],
   alphaCSR[ 5 ][ 92 ],
   alphaCSR[ 5 ][ 93 ],
   alphaCSR[ 5 ][ 94 ],
   alphaCSR[ 5 ][ 95 ],
   alphaCSR[ 5 ][ 96 ],
   alphaCSR[ 5 ][ 97 ],
   alphaCSR[ 5 ][ 98 ],
   alphaCSR[ 5 ][ 99 ],
   alphaCSR[ 5 ][ 100 ],
   alphaCSR[ 5 ][ 101 ],
   alphaCSR[ 5 ][ 102 ],
   alphaCSR[ 5 ][ 103 ],
   alphaCSR[ 5 ][ 104 ],
   alphaCSR[ 5 ][ 105 ],
   alphaCSR[ 5 ][ 106 ],
   alphaCSR[ 5 ][ 107 ],
   alphaCSR[ 5 ][ 108 ],
   alphaCSR[ 5 ][ 109 ],
   alphaCSR[ 5 ][ 110 ],
   alphaCSR[ 5 ][ 111 ],
   alphaCSR[ 5 ][ 112 ],
   alphaCSR[ 5 ][ 113 ],
   alphaCSR[ 5 ][ 114 ],
   alphaCSR[ 5 ][ 115 ],
   alphaCSR[ 5 ][ 116 ],
   alphaCSR[ 5 ][ 117 ],
   alphaCSR[ 5 ][ 118 ],
   alphaCSR[ 5 ][ 119 ],
   alphaCSR[ 5 ][ 120 ],
   alphaCSR[ 5 ][ 121 ],
   alphaCSR[ 5 ][ 122 ],
   alphaCSR[ 5 ][ 123 ],
   alphaCSR[ 5 ][ 124 ],
   alphaCSR[ 5 ][ 125 ],
   alphaCSR[ 5 ][ 126 ],
   alphaCSR[ 5 ][ 127 ],
   alphaCSR[ 5 ][ 128 ],
   alphaCSR[ 5 ][ 129 ],
   alphaCSR[ 5 ][ 130 ],
   alphaCSR[ 5 ][ 131 ],
   alphaCSR[ 5 ][ 132 ],
   alphaCSR[ 5 ][ 133 ],
   alphaCSR[ 5 ][ 134 ],
   alphaCSR[ 5 ][ 135 ],
   alphaCSR[ 5 ][ 136 ],
   alphaCSR[ 5 ][ 137 ],
   alphaCSR[ 5 ][ 138 ],
   alphaCSR[ 5 ][ 139 ],
   alphaCSR[ 5 ][ 140 ],
   alphaCSR[ 5 ][ 141 ],
   alphaCSR[ 5 ][ 142 ],
   alphaCSR[ 5 ][ 143 ],
   alphaCSR[ 5 ][ 144 ],
   alphaCSR[ 5 ][ 145 ],
   alphaCSR[ 5 ][ 146 ],
   alphaCSR[ 5 ][ 147 ],
   alphaCSR[ 5 ][ 148 ],
   alphaCSR[ 5 ][ 149 ],
   alphaCSR[ 5 ][ 150 ],
   alphaCSR[ 5 ][ 151 ],
   alphaCSR[ 5 ][ 152 ],
   alphaCSR[ 5 ][ 153 ],
   alphaCSR[ 5 ][ 154 ],
   alphaCSR[ 5 ][ 155 ],
   alphaCSR[ 5 ][ 156 ],
   alphaCSR[ 5 ][ 157 ],
   alphaCSR[ 5 ][ 158 ],
   alphaCSR[ 5 ][ 159 ],
   alphaCSR[ 5 ][ 160 ],
   alphaCSR[ 5 ][ 161 ],
   alphaCSR[ 5 ][ 162 ],
   alphaCSR[ 5 ][ 163 ],
   alphaCSR[ 5 ][ 164 ],
   alphaCSR[ 5 ][ 165 ],
   alphaCSR[ 5 ][ 166 ],
   alphaCSR[ 5 ][ 167 ],
   alphaCSR[ 5 ][ 168 ],
   alphaCSR[ 5 ][ 169 ],
   alphaCSR[ 5 ][ 170 ],
   alphaCSR[ 5 ][ 171 ],
   alphaCSR[ 5 ][ 172 ],
   alphaCSR[ 5 ][ 173 ],
   alphaCSR[ 5 ][ 174 ],
   alphaCSR[ 5 ][ 175 ],
   alphaCSR[ 5 ][ 176 ],
   alphaCSR[ 5 ][ 177 ],
   alphaCSR[ 5 ][ 178 ],
   alphaCSR[ 5 ][ 179 ],
   alphaCSR[ 5 ][ 180 ],
   alphaCSR[ 5 ][ 181 ],
   alphaCSR[ 5 ][ 182 ],
   alphaCSR[ 5 ][ 183 ],
   alphaCSR[ 5 ][ 184 ],
   alphaCSR[ 5 ][ 185 ],
   alphaCSR[ 5 ][ 186 ],
   alphaCSR[ 5 ][ 187 ],
   alphaCSR[ 5 ][ 188 ],
   alphaCSR[ 5 ][ 189 ],
   alphaCSR[ 5 ][ 190 ],
   alphaCSR[ 5 ][ 191 ],
   alphaCSR[ 5 ][ 192 ],
   alphaCSR[ 5 ][ 193 ],
   alphaCSR[ 5 ][ 194 ],
   alphaCSR[ 5 ][ 195 ],
   alphaCSR[ 5 ][ 196 ],
   alphaCSR[ 5 ][ 197 ],
   alphaCSR[ 5 ][ 198 ],
   alphaCSR[ 5 ][ 199 ],
   alphaCSR[ 5 ][ 200 ],
   alphaCSR[ 5 ][ 201 ],
   alphaCSR[ 5 ][ 202 ],
   alphaCSR[ 5 ][ 203 ],
   alphaCSR[ 5 ][ 204 ],
   alphaCSR[ 5 ][ 205 ],
   alphaCSR[ 5 ][ 206 ],
   alphaCSR[ 5 ][ 207 ],
   alphaCSR[ 5 ][ 208 ],
   alphaCSR[ 5 ][ 209 ],
   alphaCSR[ 5 ][ 210 ],
   alphaCSR[ 5 ][ 211 ],
   alphaCSR[ 5 ][ 212 ],
   alphaCSR[ 5 ][ 213 ],
   alphaCSR[ 5 ][ 214 ],
   alphaCSR[ 5 ][ 215 ],
   alphaCSR[ 5 ][ 216 ],
   alphaCSR[ 5 ][ 217 ],
   alphaCSR[ 5 ][ 218 ],
   alphaCSR[ 5 ][ 219 ],
   alphaCSR[ 5 ][ 220 ],
   alphaCSR[ 5 ][ 221 ],
   alphaCSR[ 5 ][ 222 ],
   alphaCSR[ 5 ][ 223 ],
   alphaCSR[ 5 ][ 224 ],
   alphaCSR[ 5 ][ 225 ],
   alphaCSR[ 5 ][ 226 ],
   alphaCSR[ 5 ][ 227 ],
   alphaCSR[ 5 ][ 228 ],
   alphaCSR[ 5 ][ 229 ],
   alphaCSR[ 5 ][ 230 ],
   alphaCSR[ 5 ][ 231 ],
   alphaCSR[ 5 ][ 232 ],
   alphaCSR[ 5 ][ 233 ],
   alphaCSR[ 5 ][ 234 ],
   alphaCSR[ 5 ][ 235 ],
   alphaCSR[ 5 ][ 236 ],
   alphaCSR[ 5 ][ 237 ],
   alphaCSR[ 5 ][ 238 ],
   alphaCSR[ 5 ][ 239 ],
   alphaCSR[ 5 ][ 240 ],
   alphaCSR[ 5 ][ 241 ],
   alphaCSR[ 5 ][ 242 ],
   alphaCSR[ 5 ][ 243 ],
   alphaCSR[ 5 ][ 244 ],
   alphaCSR[ 5 ][ 245 ],
   alphaCSR[ 5 ][ 246 ],
   alphaCSR[ 5 ][ 247 ],
   alphaCSR[ 5 ][ 248 ],
   alphaCSR[ 5 ][ 249 ],
   alphaCSR[ 5 ][ 250 ],
   alphaCSR[ 5 ][ 251 ],
   alphaCSR[ 5 ][ 252 ],
   alphaCSR[ 5 ][ 253 ],
   alphaCSR[ 5 ][ 254 ],
   alphaCSR[ 5 ][ 255 ],
   alphaCSR[ 5 ][ 256 ],
   alphaCSR[ 5 ][ 257 ],
   alphaCSR[ 5 ][ 258 ],
   alphaCSR[ 5 ][ 259 ],
   alphaCSR[ 5 ][ 260 ],
   alphaCSR[ 5 ][ 261 ],
   alphaCSR[ 5 ][ 262 ],
   alphaCSR[ 5 ][ 263 ],
   alphaCSR[ 5 ][ 264 ],
   alphaCSR[ 5 ][ 265 ],
   alphaCSR[ 5 ][ 266 ],
   alphaCSR[ 5 ][ 267 ],
   alphaCSR[ 5 ][ 268 ],
   alphaCSR[ 5 ][ 269 ],
   alphaCSR[ 5 ][ 270 ],
   alphaCSR[ 5 ][ 271 ],
   alphaCSR[ 5 ][ 272 ],
   alphaCSR[ 5 ][ 273 ],
   alphaCSR[ 5 ][ 274 ],
   alphaCSR[ 5 ][ 275 ],
   alphaCSR[ 5 ][ 276 ],
   alphaCSR[ 5 ][ 277 ],
   alphaCSR[ 5 ][ 278 ],
   alphaCSR[ 5 ][ 279 ],
   alphaCSR[ 5 ][ 280 ],
   alphaCSR[ 5 ][ 281 ],
   alphaCSR[ 5 ][ 282 ],
   alphaCSR[ 5 ][ 283 ],
   alphaCSR[ 5 ][ 284 ],
   alphaCSR[ 5 ][ 285 ],
   alphaCSR[ 5 ][ 286 ],
   alphaCSR[ 5 ][ 287 ],
   alphaCSR[ 5 ][ 288 ],
   alphaCSR[ 5 ][ 289 ],
   alphaCSR[ 5 ][ 290 ],
   alphaCSR[ 5 ][ 291 ],
   alphaCSR[ 5 ][ 292 ],
   alphaCSR[ 5 ][ 293 ],
   alphaCSR[ 5 ][ 294 ],
   alphaCSR[ 5 ][ 295 ],
   alphaCSR[ 5 ][ 296 ],
   alphaCSR[ 5 ][ 297 ],
   alphaCSR[ 5 ][ 298 ],
   alphaCSR[ 5 ][ 299 ],
   alphaCSR[ 5 ][ 300 ],
   alphaCSR[ 5 ][ 301 ],
   alphaCSR[ 5 ][ 302 ],
   alphaCSR[ 5 ][ 303 ],
   alphaCSR[ 5 ][ 304 ],
   alphaCSR[ 5 ][ 305 ],
   alphaCSR[ 5 ][ 306 ],
   alphaCSR[ 5 ][ 307 ],
   alphaCSR[ 5 ][ 308 ],
   alphaCSR[ 5 ][ 309 ],
   alphaCSR[ 5 ][ 310 ],
   alphaCSR[ 5 ][ 311 ],
   alphaCSR[ 5 ][ 312 ],
   alphaCSR[ 5 ][ 313 ],
   alphaCSR[ 5 ][ 314 ],
   alphaCSR[ 5 ][ 315 ],
   alphaCSR[ 5 ][ 316 ],
   alphaCSR[ 5 ][ 317 ],
   alphaCSR[ 5 ][ 318 ],
   alphaCSR[ 5 ][ 319 ],
   alphaCSR[ 5 ][ 320 ],
   alphaCSR[ 5 ][ 321 ],
   alphaCSR[ 5 ][ 322 ],
   alphaCSR[ 5 ][ 323 ],
   alphaCSR[ 5 ][ 324 ],
   alphaCSR[ 5 ][ 325 ],
   alphaCSR[ 5 ][ 326 ],
   alphaCSR[ 5 ][ 327 ],
   alphaCSR[ 5 ][ 328 ],
   alphaCSR[ 5 ][ 329 ],
   alphaCSR[ 5 ][ 330 ],
   alphaCSR[ 5 ][ 331 ],
   alphaCSR[ 5 ][ 332 ],
   alphaCSR[ 5 ][ 333 ],
   alphaCSR[ 5 ][ 334 ],
   alphaCSR[ 5 ][ 335 ],
   alphaCSR[ 5 ][ 336 ],
   alphaCSR[ 5 ][ 337 ],
   alphaCSR[ 5 ][ 338 ],
   alphaCSR[ 5 ][ 339 ],
   alphaCSR[ 5 ][ 340 ],
   alphaCSR[ 5 ][ 341 ],
   alphaCSR[ 5 ][ 342 ],
   alphaCSR[ 5 ][ 343 ],
   alphaCSR[ 5 ][ 344 ],
   alphaCSR[ 5 ][ 345 ],
   alphaCSR[ 5 ][ 346 ],
   alphaCSR[ 5 ][ 347 ],
   alphaCSR[ 5 ][ 348 ],
   alphaCSR[ 5 ][ 349 ],
   alphaCSR[ 5 ][ 350 ],
   alphaCSR[ 5 ][ 351 ],
   alphaCSR[ 5 ][ 352 ],
   alphaCSR[ 5 ][ 353 ],
   alphaCSR[ 5 ][ 354 ],
   alphaCSR[ 5 ][ 355 ],
   alphaCSR[ 5 ][ 356 ],
   alphaCSR[ 5 ][ 357 ],
   alphaCSR[ 5 ][ 358 ],
   alphaCSR[ 5 ][ 359 ],
   alphaCSR[ 5 ][ 360 ],
   alphaCSR[ 5 ][ 361 ],
   alphaCSR[ 5 ][ 362 ],
   alphaCSR[ 5 ][ 363 ],
   alphaCSR[ 5 ][ 364 ],
   alphaCSR[ 5 ][ 365 ],
   alphaCSR[ 5 ][ 366 ],
   alphaCSR[ 5 ][ 367 ],
   alphaCSR[ 5 ][ 368 ],
   alphaCSR[ 5 ][ 369 ],
   alphaCSR[ 5 ][ 370 ],
   alphaCSR[ 5 ][ 371 ],
   alphaCSR[ 5 ][ 372 ],
   alphaCSR[ 5 ][ 373 ],
   alphaCSR[ 5 ][ 374 ],
   alphaCSR[ 5 ][ 375 ],
   alphaCSR[ 5 ][ 376 ],
   alphaCSR[ 5 ][ 377 ],
   alphaCSR[ 5 ][ 378 ],
   alphaCSR[ 5 ][ 379 ],
   alphaCSR[ 5 ][ 380 ],
   alphaCSR[ 5 ][ 381 ],
   alphaCSR[ 5 ][ 382 ],
   alphaCSR[ 5 ][ 383 ],
   alphaCSR[ 6 ][ 0 ],
   alphaCSR[ 6 ][ 1 ],
   alphaCSR[ 6 ][ 2 ],
   alphaCSR[ 6 ][ 3 ],
   alphaCSR[ 6 ][ 4 ],
   alphaCSR[ 6 ][ 5 ],
   alphaCSR[ 6 ][ 6 ],
   alphaCSR[ 6 ][ 7 ],
   alphaCSR[ 6 ][ 8 ],
   alphaCSR[ 6 ][ 9 ],
   alphaCSR[ 6 ][ 10 ],
   alphaCSR[ 6 ][ 11 ],
   alphaCSR[ 6 ][ 12 ],
   alphaCSR[ 6 ][ 13 ],
   alphaCSR[ 6 ][ 14 ],
   alphaCSR[ 6 ][ 15 ],
   alphaCSR[ 6 ][ 16 ],
   alphaCSR[ 6 ][ 17 ],
   alphaCSR[ 6 ][ 18 ],
   alphaCSR[ 6 ][ 19 ],
   alphaCSR[ 6 ][ 20 ],
   alphaCSR[ 6 ][ 21 ],
   alphaCSR[ 6 ][ 22 ],
   alphaCSR[ 6 ][ 23 ],
   alphaCSR[ 6 ][ 24 ],
   alphaCSR[ 6 ][ 25 ],
   alphaCSR[ 6 ][ 26 ],
   alphaCSR[ 6 ][ 27 ],
   alphaCSR[ 6 ][ 28 ],
   alphaCSR[ 6 ][ 29 ],
   alphaCSR[ 6 ][ 30 ],
   alphaCSR[ 6 ][ 31 ],
   alphaCSR[ 6 ][ 32 ],
   alphaCSR[ 6 ][ 33 ],
   alphaCSR[ 6 ][ 34 ],
   alphaCSR[ 6 ][ 35 ],
   alphaCSR[ 6 ][ 36 ],
   alphaCSR[ 6 ][ 37 ],
   alphaCSR[ 6 ][ 38 ],
   alphaCSR[ 6 ][ 39 ],
   alphaCSR[ 6 ][ 40 ],
   alphaCSR[ 6 ][ 41 ],
   alphaCSR[ 6 ][ 42 ],
   alphaCSR[ 6 ][ 43 ],
   alphaCSR[ 6 ][ 44 ],
   alphaCSR[ 6 ][ 45 ],
   alphaCSR[ 6 ][ 46 ],
   alphaCSR[ 6 ][ 47 ],
   alphaCSR[ 6 ][ 48 ],
   alphaCSR[ 6 ][ 49 ],
   alphaCSR[ 6 ][ 50 ],
   alphaCSR[ 6 ][ 51 ],
   alphaCSR[ 6 ][ 52 ],
   alphaCSR[ 6 ][ 53 ],
   alphaCSR[ 6 ][ 54 ],
   alphaCSR[ 6 ][ 55 ],
   alphaCSR[ 6 ][ 56 ],
   alphaCSR[ 6 ][ 57 ],
   alphaCSR[ 6 ][ 58 ],
   alphaCSR[ 6 ][ 59 ],
   alphaCSR[ 6 ][ 60 ],
   alphaCSR[ 6 ][ 61 ],
   alphaCSR[ 6 ][ 62 ],
   alphaCSR[ 6 ][ 63 ],
   alphaCSR[ 6 ][ 64 ],
   alphaCSR[ 6 ][ 65 ],
   alphaCSR[ 6 ][ 66 ],
   alphaCSR[ 6 ][ 67 ],
   alphaCSR[ 6 ][ 68 ],
   alphaCSR[ 6 ][ 69 ],
   alphaCSR[ 6 ][ 70 ],
   alphaCSR[ 6 ][ 71 ],
   alphaCSR[ 6 ][ 72 ],
   alphaCSR[ 6 ][ 73 ],
   alphaCSR[ 6 ][ 74 ],
   alphaCSR[ 6 ][ 75 ],
   alphaCSR[ 6 ][ 76 ],
   alphaCSR[ 6 ][ 77 ],
   alphaCSR[ 6 ][ 78 ],
   alphaCSR[ 6 ][ 79 ],
   alphaCSR[ 6 ][ 80 ],
   alphaCSR[ 6 ][ 81 ],
   alphaCSR[ 6 ][ 82 ],
   alphaCSR[ 6 ][ 83 ],
   alphaCSR[ 6 ][ 84 ],
   alphaCSR[ 6 ][ 85 ],
   alphaCSR[ 6 ][ 86 ],
   alphaCSR[ 6 ][ 87 ],
   alphaCSR[ 6 ][ 88 ],
   alphaCSR[ 6 ][ 89 ],
   alphaCSR[ 6 ][ 90 ],
   alphaCSR[ 6 ][ 91 ],
   alphaCSR[ 6 ][ 92 ],
   alphaCSR[ 6 ][ 93 ],
   alphaCSR[ 6 ][ 94 ],
   alphaCSR[ 6 ][ 95 ],
   alphaCSR[ 6 ][ 96 ],
   alphaCSR[ 6 ][ 97 ],
   alphaCSR[ 6 ][ 98 ],
   alphaCSR[ 6 ][ 99 ],
   alphaCSR[ 6 ][ 100 ],
   alphaCSR[ 6 ][ 101 ],
   alphaCSR[ 6 ][ 102 ],
   alphaCSR[ 6 ][ 103 ],
   alphaCSR[ 6 ][ 104 ],
   alphaCSR[ 6 ][ 105 ],
   alphaCSR[ 6 ][ 106 ],
   alphaCSR[ 6 ][ 107 ],
   alphaCSR[ 6 ][ 108 ],
   alphaCSR[ 6 ][ 109 ],
   alphaCSR[ 6 ][ 110 ],
   alphaCSR[ 6 ][ 111 ],
   alphaCSR[ 6 ][ 112 ],
   alphaCSR[ 6 ][ 113 ],
   alphaCSR[ 6 ][ 114 ],
   alphaCSR[ 6 ][ 115 ],
   alphaCSR[ 6 ][ 116 ],
   alphaCSR[ 6 ][ 117 ],
   alphaCSR[ 6 ][ 118 ],
   alphaCSR[ 6 ][ 119 ],
   alphaCSR[ 6 ][ 120 ],
   alphaCSR[ 6 ][ 121 ],
   alphaCSR[ 6 ][ 122 ],
   alphaCSR[ 6 ][ 123 ],
   alphaCSR[ 6 ][ 124 ],
   alphaCSR[ 6 ][ 125 ],
   alphaCSR[ 6 ][ 126 ],
   alphaCSR[ 6 ][ 127 ],
   alphaCSR[ 6 ][ 128 ],
   alphaCSR[ 6 ][ 129 ],
   alphaCSR[ 6 ][ 130 ],
   alphaCSR[ 6 ][ 131 ],
   alphaCSR[ 6 ][ 132 ],
   alphaCSR[ 6 ][ 133 ],
   alphaCSR[ 6 ][ 134 ],
   alphaCSR[ 6 ][ 135 ],
   alphaCSR[ 6 ][ 136 ],
   alphaCSR[ 6 ][ 137 ],
   alphaCSR[ 6 ][ 138 ],
   alphaCSR[ 6 ][ 139 ],
   alphaCSR[ 6 ][ 140 ],
   alphaCSR[ 6 ][ 141 ],
   alphaCSR[ 6 ][ 142 ],
   alphaCSR[ 6 ][ 143 ],
   alphaCSR[ 6 ][ 144 ],
   alphaCSR[ 6 ][ 145 ],
   alphaCSR[ 6 ][ 146 ],
   alphaCSR[ 6 ][ 147 ],
   alphaCSR[ 6 ][ 148 ],
   alphaCSR[ 6 ][ 149 ],
   alphaCSR[ 6 ][ 150 ],
   alphaCSR[ 6 ][ 151 ],
   alphaCSR[ 6 ][ 152 ],
   alphaCSR[ 6 ][ 153 ],
   alphaCSR[ 6 ][ 154 ],
   alphaCSR[ 6 ][ 155 ],
   alphaCSR[ 6 ][ 156 ],
   alphaCSR[ 6 ][ 157 ],
   alphaCSR[ 6 ][ 158 ],
   alphaCSR[ 6 ][ 159 ],
   alphaCSR[ 6 ][ 160 ],
   alphaCSR[ 6 ][ 161 ],
   alphaCSR[ 6 ][ 162 ],
   alphaCSR[ 6 ][ 163 ],
   alphaCSR[ 6 ][ 164 ],
   alphaCSR[ 6 ][ 165 ],
   alphaCSR[ 6 ][ 166 ],
   alphaCSR[ 6 ][ 167 ],
   alphaCSR[ 6 ][ 168 ],
   alphaCSR[ 6 ][ 169 ],
   alphaCSR[ 6 ][ 170 ],
   alphaCSR[ 6 ][ 171 ],
   alphaCSR[ 6 ][ 172 ],
   alphaCSR[ 6 ][ 173 ],
   alphaCSR[ 6 ][ 174 ],
   alphaCSR[ 6 ][ 175 ],
   alphaCSR[ 6 ][ 176 ],
   alphaCSR[ 6 ][ 177 ],
   alphaCSR[ 6 ][ 178 ],
   alphaCSR[ 6 ][ 179 ],
   alphaCSR[ 6 ][ 180 ],
   alphaCSR[ 6 ][ 181 ],
   alphaCSR[ 6 ][ 182 ],
   alphaCSR[ 6 ][ 183 ],
   alphaCSR[ 6 ][ 184 ],
   alphaCSR[ 6 ][ 185 ],
   alphaCSR[ 6 ][ 186 ],
   alphaCSR[ 6 ][ 187 ],
   alphaCSR[ 6 ][ 188 ],
   alphaCSR[ 6 ][ 189 ],
   alphaCSR[ 6 ][ 190 ],
   alphaCSR[ 6 ][ 191 ],
   alphaCSR[ 6 ][ 192 ],
   alphaCSR[ 6 ][ 193 ],
   alphaCSR[ 6 ][ 194 ],
   alphaCSR[ 6 ][ 195 ],
   alphaCSR[ 6 ][ 196 ],
   alphaCSR[ 6 ][ 197 ],
   alphaCSR[ 6 ][ 198 ],
   alphaCSR[ 6 ][ 199 ],
   alphaCSR[ 6 ][ 200 ],
   alphaCSR[ 6 ][ 201 ],
   alphaCSR[ 6 ][ 202 ],
   alphaCSR[ 6 ][ 203 ],
   alphaCSR[ 6 ][ 204 ],
   alphaCSR[ 6 ][ 205 ],
   alphaCSR[ 6 ][ 206 ],
   alphaCSR[ 6 ][ 207 ],
   alphaCSR[ 6 ][ 208 ],
   alphaCSR[ 6 ][ 209 ],
   alphaCSR[ 6 ][ 210 ],
   alphaCSR[ 6 ][ 211 ],
   alphaCSR[ 6 ][ 212 ],
   alphaCSR[ 6 ][ 213 ],
   alphaCSR[ 6 ][ 214 ],
   alphaCSR[ 6 ][ 215 ],
   alphaCSR[ 6 ][ 216 ],
   alphaCSR[ 6 ][ 217 ],
   alphaCSR[ 6 ][ 218 ],
   alphaCSR[ 6 ][ 219 ],
   alphaCSR[ 6 ][ 220 ],
   alphaCSR[ 6 ][ 221 ],
   alphaCSR[ 6 ][ 222 ],
   alphaCSR[ 6 ][ 223 ],
   alphaCSR[ 6 ][ 224 ],
   alphaCSR[ 6 ][ 225 ],
   alphaCSR[ 6 ][ 226 ],
   alphaCSR[ 6 ][ 227 ],
   alphaCSR[ 6 ][ 228 ],
   alphaCSR[ 6 ][ 229 ],
   alphaCSR[ 6 ][ 230 ],
   alphaCSR[ 6 ][ 231 ],
   alphaCSR[ 6 ][ 232 ],
   alphaCSR[ 6 ][ 233 ],
   alphaCSR[ 6 ][ 234 ],
   alphaCSR[ 6 ][ 235 ],
   alphaCSR[ 6 ][ 236 ],
   alphaCSR[ 6 ][ 237 ],
   alphaCSR[ 6 ][ 238 ],
   alphaCSR[ 6 ][ 239 ],
   alphaCSR[ 6 ][ 240 ],
   alphaCSR[ 6 ][ 241 ],
   alphaCSR[ 6 ][ 242 ],
   alphaCSR[ 6 ][ 243 ],
   alphaCSR[ 6 ][ 244 ],
   alphaCSR[ 6 ][ 245 ],
   alphaCSR[ 6 ][ 246 ],
   alphaCSR[ 6 ][ 247 ],
   alphaCSR[ 6 ][ 248 ],
   alphaCSR[ 6 ][ 249 ],
   alphaCSR[ 6 ][ 250 ],
   alphaCSR[ 6 ][ 251 ],
   alphaCSR[ 6 ][ 252 ],
   alphaCSR[ 6 ][ 253 ],
   alphaCSR[ 6 ][ 254 ],
   alphaCSR[ 6 ][ 255 ],
   alphaCSR[ 6 ][ 256 ],
   alphaCSR[ 6 ][ 257 ],
   alphaCSR[ 6 ][ 258 ],
   alphaCSR[ 6 ][ 259 ],
   alphaCSR[ 6 ][ 260 ],
   alphaCSR[ 6 ][ 261 ],
   alphaCSR[ 6 ][ 262 ],
   alphaCSR[ 6 ][ 263 ],
   alphaCSR[ 6 ][ 264 ],
   alphaCSR[ 6 ][ 265 ],
   alphaCSR[ 6 ][ 266 ],
   alphaCSR[ 6 ][ 267 ],
   alphaCSR[ 6 ][ 268 ],
   alphaCSR[ 6 ][ 269 ],
   alphaCSR[ 6 ][ 270 ],
   alphaCSR[ 6 ][ 271 ],
   alphaCSR[ 6 ][ 272 ],
   alphaCSR[ 6 ][ 273 ],
   alphaCSR[ 6 ][ 274 ],
   alphaCSR[ 6 ][ 275 ],
   alphaCSR[ 6 ][ 276 ],
   alphaCSR[ 6 ][ 277 ],
   alphaCSR[ 6 ][ 278 ],
   alphaCSR[ 6 ][ 279 ],
   alphaCSR[ 6 ][ 280 ],
   alphaCSR[ 6 ][ 281 ],
   alphaCSR[ 6 ][ 282 ],
   alphaCSR[ 6 ][ 283 ],
   alphaCSR[ 6 ][ 284 ],
   alphaCSR[ 6 ][ 285 ],
   alphaCSR[ 6 ][ 286 ],
   alphaCSR[ 6 ][ 287 ],
   alphaCSR[ 6 ][ 288 ],
   alphaCSR[ 6 ][ 289 ],
   alphaCSR[ 6 ][ 290 ],
   alphaCSR[ 6 ][ 291 ],
   alphaCSR[ 6 ][ 292 ],
   alphaCSR[ 6 ][ 293 ],
   alphaCSR[ 6 ][ 294 ],
   alphaCSR[ 6 ][ 295 ],
   alphaCSR[ 6 ][ 296 ],
   alphaCSR[ 6 ][ 297 ],
   alphaCSR[ 6 ][ 298 ],
   alphaCSR[ 6 ][ 299 ],
   alphaCSR[ 6 ][ 300 ],
   alphaCSR[ 6 ][ 301 ],
   alphaCSR[ 6 ][ 302 ],
   alphaCSR[ 6 ][ 303 ],
   alphaCSR[ 6 ][ 304 ],
   alphaCSR[ 6 ][ 305 ],
   alphaCSR[ 6 ][ 306 ],
   alphaCSR[ 6 ][ 307 ],
   alphaCSR[ 6 ][ 308 ],
   alphaCSR[ 6 ][ 309 ],
   alphaCSR[ 6 ][ 310 ],
   alphaCSR[ 6 ][ 311 ],
   alphaCSR[ 6 ][ 312 ],
   alphaCSR[ 6 ][ 313 ],
   alphaCSR[ 6 ][ 314 ],
   alphaCSR[ 6 ][ 315 ],
   alphaCSR[ 6 ][ 316 ],
   alphaCSR[ 6 ][ 317 ],
   alphaCSR[ 6 ][ 318 ],
   alphaCSR[ 6 ][ 319 ],
   alphaCSR[ 6 ][ 320 ],
   alphaCSR[ 6 ][ 321 ],
   alphaCSR[ 6 ][ 322 ],
   alphaCSR[ 6 ][ 323 ],
   alphaCSR[ 6 ][ 324 ],
   alphaCSR[ 6 ][ 325 ],
   alphaCSR[ 6 ][ 326 ],
   alphaCSR[ 6 ][ 327 ],
   alphaCSR[ 6 ][ 328 ],
   alphaCSR[ 6 ][ 329 ],
   alphaCSR[ 6 ][ 330 ],
   alphaCSR[ 6 ][ 331 ],
   alphaCSR[ 6 ][ 332 ],
   alphaCSR[ 6 ][ 333 ],
   alphaCSR[ 6 ][ 334 ],
   alphaCSR[ 6 ][ 335 ],
   alphaCSR[ 6 ][ 336 ],
   alphaCSR[ 6 ][ 337 ],
   alphaCSR[ 6 ][ 338 ],
   alphaCSR[ 6 ][ 339 ],
   alphaCSR[ 6 ][ 340 ],
   alphaCSR[ 6 ][ 341 ],
   alphaCSR[ 6 ][ 342 ],
   alphaCSR[ 6 ][ 343 ],
   alphaCSR[ 6 ][ 344 ],
   alphaCSR[ 6 ][ 345 ],
   alphaCSR[ 6 ][ 346 ],
   alphaCSR[ 6 ][ 347 ],
   alphaCSR[ 6 ][ 348 ],
   alphaCSR[ 6 ][ 349 ],
   alphaCSR[ 6 ][ 350 ],
   alphaCSR[ 6 ][ 351 ],
   alphaCSR[ 6 ][ 352 ],
   alphaCSR[ 6 ][ 353 ],
   alphaCSR[ 6 ][ 354 ],
   alphaCSR[ 6 ][ 355 ],
   alphaCSR[ 6 ][ 356 ],
   alphaCSR[ 6 ][ 357 ],
   alphaCSR[ 6 ][ 358 ],
   alphaCSR[ 6 ][ 359 ],
   alphaCSR[ 6 ][ 360 ],
   alphaCSR[ 6 ][ 361 ],
   alphaCSR[ 6 ][ 362 ],
   alphaCSR[ 6 ][ 363 ],
   alphaCSR[ 6 ][ 364 ],
   alphaCSR[ 6 ][ 365 ],
   alphaCSR[ 6 ][ 366 ],
   alphaCSR[ 6 ][ 367 ],
   alphaCSR[ 6 ][ 368 ],
   alphaCSR[ 6 ][ 369 ],
   alphaCSR[ 6 ][ 370 ],
   alphaCSR[ 6 ][ 371 ],
   alphaCSR[ 6 ][ 372 ],
   alphaCSR[ 6 ][ 373 ],
   alphaCSR[ 6 ][ 374 ],
   alphaCSR[ 6 ][ 375 ],
   alphaCSR[ 6 ][ 376 ],
   alphaCSR[ 6 ][ 377 ],
   alphaCSR[ 6 ][ 378 ],
   alphaCSR[ 6 ][ 379 ],
   alphaCSR[ 6 ][ 380 ],
   alphaCSR[ 6 ][ 381 ],
   alphaCSR[ 6 ][ 382 ],
   alphaCSR[ 6 ][ 383 ],
   alphaCSR[ 7 ][ 0 ],
   alphaCSR[ 7 ][ 1 ],
   alphaCSR[ 7 ][ 2 ],
   alphaCSR[ 7 ][ 3 ],
   alphaCSR[ 7 ][ 4 ],
   alphaCSR[ 7 ][ 5 ],
   alphaCSR[ 7 ][ 6 ],
   alphaCSR[ 7 ][ 7 ],
   alphaCSR[ 7 ][ 8 ],
   alphaCSR[ 7 ][ 9 ],
   alphaCSR[ 7 ][ 10 ],
   alphaCSR[ 7 ][ 11 ],
   alphaCSR[ 7 ][ 12 ],
   alphaCSR[ 7 ][ 13 ],
   alphaCSR[ 7 ][ 14 ],
   alphaCSR[ 7 ][ 15 ],
   alphaCSR[ 7 ][ 16 ],
   alphaCSR[ 7 ][ 17 ],
   alphaCSR[ 7 ][ 18 ],
   alphaCSR[ 7 ][ 19 ],
   alphaCSR[ 7 ][ 20 ],
   alphaCSR[ 7 ][ 21 ],
   alphaCSR[ 7 ][ 22 ],
   alphaCSR[ 7 ][ 23 ],
   alphaCSR[ 7 ][ 24 ],
   alphaCSR[ 7 ][ 25 ],
   alphaCSR[ 7 ][ 26 ],
   alphaCSR[ 7 ][ 27 ],
   alphaCSR[ 7 ][ 28 ],
   alphaCSR[ 7 ][ 29 ],
   alphaCSR[ 7 ][ 30 ],
   alphaCSR[ 7 ][ 31 ],
   alphaCSR[ 7 ][ 32 ],
   alphaCSR[ 7 ][ 33 ],
   alphaCSR[ 7 ][ 34 ],
   alphaCSR[ 7 ][ 35 ],
   alphaCSR[ 7 ][ 36 ],
   alphaCSR[ 7 ][ 37 ],
   alphaCSR[ 7 ][ 38 ],
   alphaCSR[ 7 ][ 39 ],
   alphaCSR[ 7 ][ 40 ],
   alphaCSR[ 7 ][ 41 ],
   alphaCSR[ 7 ][ 42 ],
   alphaCSR[ 7 ][ 43 ],
   alphaCSR[ 7 ][ 44 ],
   alphaCSR[ 7 ][ 45 ],
   alphaCSR[ 7 ][ 46 ],
   alphaCSR[ 7 ][ 47 ],
   alphaCSR[ 7 ][ 48 ],
   alphaCSR[ 7 ][ 49 ],
   alphaCSR[ 7 ][ 50 ],
   alphaCSR[ 7 ][ 51 ],
   alphaCSR[ 7 ][ 52 ],
   alphaCSR[ 7 ][ 53 ],
   alphaCSR[ 7 ][ 54 ],
   alphaCSR[ 7 ][ 55 ],
   alphaCSR[ 7 ][ 56 ],
   alphaCSR[ 7 ][ 57 ],
   alphaCSR[ 7 ][ 58 ],
   alphaCSR[ 7 ][ 59 ],
   alphaCSR[ 7 ][ 60 ],
   alphaCSR[ 7 ][ 61 ],
   alphaCSR[ 7 ][ 62 ],
   alphaCSR[ 7 ][ 63 ],
   alphaCSR[ 7 ][ 64 ],
   alphaCSR[ 7 ][ 65 ],
   alphaCSR[ 7 ][ 66 ],
   alphaCSR[ 7 ][ 67 ],
   alphaCSR[ 7 ][ 68 ],
   alphaCSR[ 7 ][ 69 ],
   alphaCSR[ 7 ][ 70 ],
   alphaCSR[ 7 ][ 71 ],
   alphaCSR[ 7 ][ 72 ],
   alphaCSR[ 7 ][ 73 ],
   alphaCSR[ 7 ][ 74 ],
   alphaCSR[ 7 ][ 75 ],
   alphaCSR[ 7 ][ 76 ],
   alphaCSR[ 7 ][ 77 ],
   alphaCSR[ 7 ][ 78 ],
   alphaCSR[ 7 ][ 79 ],
   alphaCSR[ 7 ][ 80 ],
   alphaCSR[ 7 ][ 81 ],
   alphaCSR[ 7 ][ 82 ],
   alphaCSR[ 7 ][ 83 ],
   alphaCSR[ 7 ][ 84 ],
   alphaCSR[ 7 ][ 85 ],
   alphaCSR[ 7 ][ 86 ],
   alphaCSR[ 7 ][ 87 ],
   alphaCSR[ 7 ][ 88 ],
   alphaCSR[ 7 ][ 89 ],
   alphaCSR[ 7 ][ 90 ],
   alphaCSR[ 7 ][ 91 ],
   alphaCSR[ 7 ][ 92 ],
   alphaCSR[ 7 ][ 93 ],
   alphaCSR[ 7 ][ 94 ],
   alphaCSR[ 7 ][ 95 ],
   alphaCSR[ 7 ][ 96 ],
   alphaCSR[ 7 ][ 97 ],
   alphaCSR[ 7 ][ 98 ],
   alphaCSR[ 7 ][ 99 ],
   alphaCSR[ 7 ][ 100 ],
   alphaCSR[ 7 ][ 101 ],
   alphaCSR[ 7 ][ 102 ],
   alphaCSR[ 7 ][ 103 ],
   alphaCSR[ 7 ][ 104 ],
   alphaCSR[ 7 ][ 105 ],
   alphaCSR[ 7 ][ 106 ],
   alphaCSR[ 7 ][ 107 ],
   alphaCSR[ 7 ][ 108 ],
   alphaCSR[ 7 ][ 109 ],
   alphaCSR[ 7 ][ 110 ],
   alphaCSR[ 7 ][ 111 ],
   alphaCSR[ 7 ][ 112 ],
   alphaCSR[ 7 ][ 113 ],
   alphaCSR[ 7 ][ 114 ],
   alphaCSR[ 7 ][ 115 ],
   alphaCSR[ 7 ][ 116 ],
   alphaCSR[ 7 ][ 117 ],
   alphaCSR[ 7 ][ 118 ],
   alphaCSR[ 7 ][ 119 ],
   alphaCSR[ 7 ][ 120 ],
   alphaCSR[ 7 ][ 121 ],
   alphaCSR[ 7 ][ 122 ],
   alphaCSR[ 7 ][ 123 ],
   alphaCSR[ 7 ][ 124 ],
   alphaCSR[ 7 ][ 125 ],
   alphaCSR[ 7 ][ 126 ],
   alphaCSR[ 7 ][ 127 ],
   alphaCSR[ 7 ][ 128 ],
   alphaCSR[ 7 ][ 129 ],
   alphaCSR[ 7 ][ 130 ],
   alphaCSR[ 7 ][ 131 ],
   alphaCSR[ 7 ][ 132 ],
   alphaCSR[ 7 ][ 133 ],
   alphaCSR[ 7 ][ 134 ],
   alphaCSR[ 7 ][ 135 ],
   alphaCSR[ 7 ][ 136 ],
   alphaCSR[ 7 ][ 137 ],
   alphaCSR[ 7 ][ 138 ],
   alphaCSR[ 7 ][ 139 ],
   alphaCSR[ 7 ][ 140 ],
   alphaCSR[ 7 ][ 141 ],
   alphaCSR[ 7 ][ 142 ],
   alphaCSR[ 7 ][ 143 ],
   alphaCSR[ 7 ][ 144 ],
   alphaCSR[ 7 ][ 145 ],
   alphaCSR[ 7 ][ 146 ],
   alphaCSR[ 7 ][ 147 ],
   alphaCSR[ 7 ][ 148 ],
   alphaCSR[ 7 ][ 149 ],
   alphaCSR[ 7 ][ 150 ],
   alphaCSR[ 7 ][ 151 ],
   alphaCSR[ 7 ][ 152 ],
   alphaCSR[ 7 ][ 153 ],
   alphaCSR[ 7 ][ 154 ],
   alphaCSR[ 7 ][ 155 ],
   alphaCSR[ 7 ][ 156 ],
   alphaCSR[ 7 ][ 157 ],
   alphaCSR[ 7 ][ 158 ],
   alphaCSR[ 7 ][ 159 ],
   alphaCSR[ 7 ][ 160 ],
   alphaCSR[ 7 ][ 161 ],
   alphaCSR[ 7 ][ 162 ],
   alphaCSR[ 7 ][ 163 ],
   alphaCSR[ 7 ][ 164 ],
   alphaCSR[ 7 ][ 165 ],
   alphaCSR[ 7 ][ 166 ],
   alphaCSR[ 7 ][ 167 ],
   alphaCSR[ 7 ][ 168 ],
   alphaCSR[ 7 ][ 169 ],
   alphaCSR[ 7 ][ 170 ],
   alphaCSR[ 7 ][ 171 ],
   alphaCSR[ 7 ][ 172 ],
   alphaCSR[ 7 ][ 173 ],
   alphaCSR[ 7 ][ 174 ],
   alphaCSR[ 7 ][ 175 ],
   alphaCSR[ 7 ][ 176 ],
   alphaCSR[ 7 ][ 177 ],
   alphaCSR[ 7 ][ 178 ],
   alphaCSR[ 7 ][ 179 ],
   alphaCSR[ 7 ][ 180 ],
   alphaCSR[ 7 ][ 181 ],
   alphaCSR[ 7 ][ 182 ],
   alphaCSR[ 7 ][ 183 ],
   alphaCSR[ 7 ][ 184 ],
   alphaCSR[ 7 ][ 185 ],
   alphaCSR[ 7 ][ 186 ],
   alphaCSR[ 7 ][ 187 ],
   alphaCSR[ 7 ][ 188 ],
   alphaCSR[ 7 ][ 189 ],
   alphaCSR[ 7 ][ 190 ],
   alphaCSR[ 7 ][ 191 ],
   alphaCSR[ 7 ][ 192 ],
   alphaCSR[ 7 ][ 193 ],
   alphaCSR[ 7 ][ 194 ],
   alphaCSR[ 7 ][ 195 ],
   alphaCSR[ 7 ][ 196 ],
   alphaCSR[ 7 ][ 197 ],
   alphaCSR[ 7 ][ 198 ],
   alphaCSR[ 7 ][ 199 ],
   alphaCSR[ 7 ][ 200 ],
   alphaCSR[ 7 ][ 201 ],
   alphaCSR[ 7 ][ 202 ],
   alphaCSR[ 7 ][ 203 ],
   alphaCSR[ 7 ][ 204 ],
   alphaCSR[ 7 ][ 205 ],
   alphaCSR[ 7 ][ 206 ],
   alphaCSR[ 7 ][ 207 ],
   alphaCSR[ 7 ][ 208 ],
   alphaCSR[ 7 ][ 209 ],
   alphaCSR[ 7 ][ 210 ],
   alphaCSR[ 7 ][ 211 ],
   alphaCSR[ 7 ][ 212 ],
   alphaCSR[ 7 ][ 213 ],
   alphaCSR[ 7 ][ 214 ],
   alphaCSR[ 7 ][ 215 ],
   alphaCSR[ 7 ][ 216 ],
   alphaCSR[ 7 ][ 217 ],
   alphaCSR[ 7 ][ 218 ],
   alphaCSR[ 7 ][ 219 ],
   alphaCSR[ 7 ][ 220 ],
   alphaCSR[ 7 ][ 221 ],
   alphaCSR[ 7 ][ 222 ],
   alphaCSR[ 7 ][ 223 ],
   alphaCSR[ 7 ][ 224 ],
   alphaCSR[ 7 ][ 225 ],
   alphaCSR[ 7 ][ 226 ],
   alphaCSR[ 7 ][ 227 ],
   alphaCSR[ 7 ][ 228 ],
   alphaCSR[ 7 ][ 229 ],
   alphaCSR[ 7 ][ 230 ],
   alphaCSR[ 7 ][ 231 ],
   alphaCSR[ 7 ][ 232 ],
   alphaCSR[ 7 ][ 233 ],
   alphaCSR[ 7 ][ 234 ],
   alphaCSR[ 7 ][ 235 ],
   alphaCSR[ 7 ][ 236 ],
   alphaCSR[ 7 ][ 237 ],
   alphaCSR[ 7 ][ 238 ],
   alphaCSR[ 7 ][ 239 ],
   alphaCSR[ 7 ][ 240 ],
   alphaCSR[ 7 ][ 241 ],
   alphaCSR[ 7 ][ 242 ],
   alphaCSR[ 7 ][ 243 ],
   alphaCSR[ 7 ][ 244 ],
   alphaCSR[ 7 ][ 245 ],
   alphaCSR[ 7 ][ 246 ],
   alphaCSR[ 7 ][ 247 ],
   alphaCSR[ 7 ][ 248 ],
   alphaCSR[ 7 ][ 249 ],
   alphaCSR[ 7 ][ 250 ],
   alphaCSR[ 7 ][ 251 ],
   alphaCSR[ 7 ][ 252 ],
   alphaCSR[ 7 ][ 253 ],
   alphaCSR[ 7 ][ 254 ],
   alphaCSR[ 7 ][ 255 ],
   alphaCSR[ 7 ][ 256 ],
   alphaCSR[ 7 ][ 257 ],
   alphaCSR[ 7 ][ 258 ],
   alphaCSR[ 7 ][ 259 ],
   alphaCSR[ 7 ][ 260 ],
   alphaCSR[ 7 ][ 261 ],
   alphaCSR[ 7 ][ 262 ],
   alphaCSR[ 7 ][ 263 ],
   alphaCSR[ 7 ][ 264 ],
   alphaCSR[ 7 ][ 265 ],
   alphaCSR[ 7 ][ 266 ],
   alphaCSR[ 7 ][ 267 ],
   alphaCSR[ 7 ][ 268 ],
   alphaCSR[ 7 ][ 269 ],
   alphaCSR[ 7 ][ 270 ],
   alphaCSR[ 7 ][ 271 ],
   alphaCSR[ 7 ][ 272 ],
   alphaCSR[ 7 ][ 273 ],
   alphaCSR[ 7 ][ 274 ],
   alphaCSR[ 7 ][ 275 ],
   alphaCSR[ 7 ][ 276 ],
   alphaCSR[ 7 ][ 277 ],
   alphaCSR[ 7 ][ 278 ],
   alphaCSR[ 7 ][ 279 ],
   alphaCSR[ 7 ][ 280 ],
   alphaCSR[ 7 ][ 281 ],
   alphaCSR[ 7 ][ 282 ],
   alphaCSR[ 7 ][ 283 ],
   alphaCSR[ 7 ][ 284 ],
   alphaCSR[ 7 ][ 285 ],
   alphaCSR[ 7 ][ 286 ],
   alphaCSR[ 7 ][ 287 ],
   alphaCSR[ 7 ][ 288 ],
   alphaCSR[ 7 ][ 289 ],
   alphaCSR[ 7 ][ 290 ],
   alphaCSR[ 7 ][ 291 ],
   alphaCSR[ 7 ][ 292 ],
   alphaCSR[ 7 ][ 293 ],
   alphaCSR[ 7 ][ 294 ],
   alphaCSR[ 7 ][ 295 ],
   alphaCSR[ 7 ][ 296 ],
   alphaCSR[ 7 ][ 297 ],
   alphaCSR[ 7 ][ 298 ],
   alphaCSR[ 7 ][ 299 ],
   alphaCSR[ 7 ][ 300 ],
   alphaCSR[ 7 ][ 301 ],
   alphaCSR[ 7 ][ 302 ],
   alphaCSR[ 7 ][ 303 ],
   alphaCSR[ 7 ][ 304 ],
   alphaCSR[ 7 ][ 305 ],
   alphaCSR[ 7 ][ 306 ],
   alphaCSR[ 7 ][ 307 ],
   alphaCSR[ 7 ][ 308 ],
   alphaCSR[ 7 ][ 309 ],
   alphaCSR[ 7 ][ 310 ],
   alphaCSR[ 7 ][ 311 ],
   alphaCSR[ 7 ][ 312 ],
   alphaCSR[ 7 ][ 313 ],
   alphaCSR[ 7 ][ 314 ],
   alphaCSR[ 7 ][ 315 ],
   alphaCSR[ 7 ][ 316 ],
   alphaCSR[ 7 ][ 317 ],
   alphaCSR[ 7 ][ 318 ],
   alphaCSR[ 7 ][ 319 ],
   alphaCSR[ 7 ][ 320 ],
   alphaCSR[ 7 ][ 321 ],
   alphaCSR[ 7 ][ 322 ],
   alphaCSR[ 7 ][ 323 ],
   alphaCSR[ 7 ][ 324 ],
   alphaCSR[ 7 ][ 325 ],
   alphaCSR[ 7 ][ 326 ],
   alphaCSR[ 7 ][ 327 ],
   alphaCSR[ 7 ][ 328 ],
   alphaCSR[ 7 ][ 329 ],
   alphaCSR[ 7 ][ 330 ],
   alphaCSR[ 7 ][ 331 ],
   alphaCSR[ 7 ][ 332 ],
   alphaCSR[ 7 ][ 333 ],
   alphaCSR[ 7 ][ 334 ],
   alphaCSR[ 7 ][ 335 ],
   alphaCSR[ 7 ][ 336 ],
   alphaCSR[ 7 ][ 337 ],
   alphaCSR[ 7 ][ 338 ],
   alphaCSR[ 7 ][ 339 ],
   alphaCSR[ 7 ][ 340 ],
   alphaCSR[ 7 ][ 341 ],
   alphaCSR[ 7 ][ 342 ],
   alphaCSR[ 7 ][ 343 ],
   alphaCSR[ 7 ][ 344 ],
   alphaCSR[ 7 ][ 345 ],
   alphaCSR[ 7 ][ 346 ],
   alphaCSR[ 7 ][ 347 ],
   alphaCSR[ 7 ][ 348 ],
   alphaCSR[ 7 ][ 349 ],
   alphaCSR[ 7 ][ 350 ],
   alphaCSR[ 7 ][ 351 ],
   alphaCSR[ 7 ][ 352 ],
   alphaCSR[ 7 ][ 353 ],
   alphaCSR[ 7 ][ 354 ],
   alphaCSR[ 7 ][ 355 ],
   alphaCSR[ 7 ][ 356 ],
   alphaCSR[ 7 ][ 357 ],
   alphaCSR[ 7 ][ 358 ],
   alphaCSR[ 7 ][ 359 ],
   alphaCSR[ 7 ][ 360 ],
   alphaCSR[ 7 ][ 361 ],
   alphaCSR[ 7 ][ 362 ],
   alphaCSR[ 7 ][ 363 ],
   alphaCSR[ 7 ][ 364 ],
   alphaCSR[ 7 ][ 365 ],
   alphaCSR[ 7 ][ 366 ],
   alphaCSR[ 7 ][ 367 ],
   alphaCSR[ 7 ][ 368 ],
   alphaCSR[ 7 ][ 369 ],
   alphaCSR[ 7 ][ 370 ],
   alphaCSR[ 7 ][ 371 ],
   alphaCSR[ 7 ][ 372 ],
   alphaCSR[ 7 ][ 373 ],
   alphaCSR[ 7 ][ 374 ],
   alphaCSR[ 7 ][ 375 ],
   alphaCSR[ 7 ][ 376 ],
   alphaCSR[ 7 ][ 377 ],
   alphaCSR[ 7 ][ 378 ],
   alphaCSR[ 7 ][ 379 ],
   alphaCSR[ 7 ][ 380 ],
   alphaCSR[ 7 ][ 381 ],
   alphaCSR[ 7 ][ 382 ],
   alphaCSR[ 7 ][ 383 ],
   alphaCSR[ 8 ][ 0 ],
   alphaCSR[ 8 ][ 1 ],
   alphaCSR[ 8 ][ 2 ],
   alphaCSR[ 8 ][ 3 ],
   alphaCSR[ 8 ][ 4 ],
   alphaCSR[ 8 ][ 5 ],
   alphaCSR[ 8 ][ 6 ],
   alphaCSR[ 8 ][ 7 ],
   alphaCSR[ 8 ][ 8 ],
   alphaCSR[ 8 ][ 9 ],
   alphaCSR[ 8 ][ 10 ],
   alphaCSR[ 8 ][ 11 ],
   alphaCSR[ 8 ][ 12 ],
   alphaCSR[ 8 ][ 13 ],
   alphaCSR[ 8 ][ 14 ],
   alphaCSR[ 8 ][ 15 ],
   alphaCSR[ 8 ][ 16 ],
   alphaCSR[ 8 ][ 17 ],
   alphaCSR[ 8 ][ 18 ],
   alphaCSR[ 8 ][ 19 ],
   alphaCSR[ 8 ][ 20 ],
   alphaCSR[ 8 ][ 21 ],
   alphaCSR[ 8 ][ 22 ],
   alphaCSR[ 8 ][ 23 ],
   alphaCSR[ 8 ][ 24 ],
   alphaCSR[ 8 ][ 25 ],
   alphaCSR[ 8 ][ 26 ],
   alphaCSR[ 8 ][ 27 ],
   alphaCSR[ 8 ][ 28 ],
   alphaCSR[ 8 ][ 29 ],
   alphaCSR[ 8 ][ 30 ],
   alphaCSR[ 8 ][ 31 ],
   alphaCSR[ 8 ][ 32 ],
   alphaCSR[ 8 ][ 33 ],
   alphaCSR[ 8 ][ 34 ],
   alphaCSR[ 8 ][ 35 ],
   alphaCSR[ 8 ][ 36 ],
   alphaCSR[ 8 ][ 37 ],
   alphaCSR[ 8 ][ 38 ],
   alphaCSR[ 8 ][ 39 ],
   alphaCSR[ 8 ][ 40 ],
   alphaCSR[ 8 ][ 41 ],
   alphaCSR[ 8 ][ 42 ],
   alphaCSR[ 8 ][ 43 ],
   alphaCSR[ 8 ][ 44 ],
   alphaCSR[ 8 ][ 45 ],
   alphaCSR[ 8 ][ 46 ],
   alphaCSR[ 8 ][ 47 ],
   alphaCSR[ 8 ][ 48 ],
   alphaCSR[ 8 ][ 49 ],
   alphaCSR[ 8 ][ 50 ],
   alphaCSR[ 8 ][ 51 ],
   alphaCSR[ 8 ][ 52 ],
   alphaCSR[ 8 ][ 53 ],
   alphaCSR[ 8 ][ 54 ],
   alphaCSR[ 8 ][ 55 ],
   alphaCSR[ 8 ][ 56 ],
   alphaCSR[ 8 ][ 57 ],
   alphaCSR[ 8 ][ 58 ],
   alphaCSR[ 8 ][ 59 ],
   alphaCSR[ 8 ][ 60 ],
   alphaCSR[ 8 ][ 61 ],
   alphaCSR[ 8 ][ 62 ],
   alphaCSR[ 8 ][ 63 ],
   alphaCSR[ 8 ][ 64 ],
   alphaCSR[ 8 ][ 65 ],
   alphaCSR[ 8 ][ 66 ],
   alphaCSR[ 8 ][ 67 ],
   alphaCSR[ 8 ][ 68 ],
   alphaCSR[ 8 ][ 69 ],
   alphaCSR[ 8 ][ 70 ],
   alphaCSR[ 8 ][ 71 ],
   alphaCSR[ 8 ][ 72 ],
   alphaCSR[ 8 ][ 73 ],
   alphaCSR[ 8 ][ 74 ],
   alphaCSR[ 8 ][ 75 ],
   alphaCSR[ 8 ][ 76 ],
   alphaCSR[ 8 ][ 77 ],
   alphaCSR[ 8 ][ 78 ],
   alphaCSR[ 8 ][ 79 ],
   alphaCSR[ 8 ][ 80 ],
   alphaCSR[ 8 ][ 81 ],
   alphaCSR[ 8 ][ 82 ],
   alphaCSR[ 8 ][ 83 ],
   alphaCSR[ 8 ][ 84 ],
   alphaCSR[ 8 ][ 85 ],
   alphaCSR[ 8 ][ 86 ],
   alphaCSR[ 8 ][ 87 ],
   alphaCSR[ 8 ][ 88 ],
   alphaCSR[ 8 ][ 89 ],
   alphaCSR[ 8 ][ 90 ],
   alphaCSR[ 8 ][ 91 ],
   alphaCSR[ 8 ][ 92 ],
   alphaCSR[ 8 ][ 93 ],
   alphaCSR[ 8 ][ 94 ],
   alphaCSR[ 8 ][ 95 ],
   alphaCSR[ 8 ][ 96 ],
   alphaCSR[ 8 ][ 97 ],
   alphaCSR[ 8 ][ 98 ],
   alphaCSR[ 8 ][ 99 ],
   alphaCSR[ 8 ][ 100 ],
   alphaCSR[ 8 ][ 101 ],
   alphaCSR[ 8 ][ 102 ],
   alphaCSR[ 8 ][ 103 ],
   alphaCSR[ 8 ][ 104 ],
   alphaCSR[ 8 ][ 105 ],
   alphaCSR[ 8 ][ 106 ],
   alphaCSR[ 8 ][ 107 ],
   alphaCSR[ 8 ][ 108 ],
   alphaCSR[ 8 ][ 109 ],
   alphaCSR[ 8 ][ 110 ],
   alphaCSR[ 8 ][ 111 ],
   alphaCSR[ 8 ][ 112 ],
   alphaCSR[ 8 ][ 113 ],
   alphaCSR[ 8 ][ 114 ],
   alphaCSR[ 8 ][ 115 ],
   alphaCSR[ 8 ][ 116 ],
   alphaCSR[ 8 ][ 117 ],
   alphaCSR[ 8 ][ 118 ],
   alphaCSR[ 8 ][ 119 ],
   alphaCSR[ 8 ][ 120 ],
   alphaCSR[ 8 ][ 121 ],
   alphaCSR[ 8 ][ 122 ],
   alphaCSR[ 8 ][ 123 ],
   alphaCSR[ 8 ][ 124 ],
   alphaCSR[ 8 ][ 125 ],
   alphaCSR[ 8 ][ 126 ],
   alphaCSR[ 8 ][ 127 ],
   alphaCSR[ 8 ][ 128 ],
   alphaCSR[ 8 ][ 129 ],
   alphaCSR[ 8 ][ 130 ],
   alphaCSR[ 8 ][ 131 ],
   alphaCSR[ 8 ][ 132 ],
   alphaCSR[ 8 ][ 133 ],
   alphaCSR[ 8 ][ 134 ],
   alphaCSR[ 8 ][ 135 ],
   alphaCSR[ 8 ][ 136 ],
   alphaCSR[ 8 ][ 137 ],
   alphaCSR[ 8 ][ 138 ],
   alphaCSR[ 8 ][ 139 ],
   alphaCSR[ 8 ][ 140 ],
   alphaCSR[ 8 ][ 141 ],
   alphaCSR[ 8 ][ 142 ],
   alphaCSR[ 8 ][ 143 ],
   alphaCSR[ 8 ][ 144 ],
   alphaCSR[ 8 ][ 145 ],
   alphaCSR[ 8 ][ 146 ],
   alphaCSR[ 8 ][ 147 ],
   alphaCSR[ 8 ][ 148 ],
   alphaCSR[ 8 ][ 149 ],
   alphaCSR[ 8 ][ 150 ],
   alphaCSR[ 8 ][ 151 ],
   alphaCSR[ 8 ][ 152 ],
   alphaCSR[ 8 ][ 153 ],
   alphaCSR[ 8 ][ 154 ],
   alphaCSR[ 8 ][ 155 ],
   alphaCSR[ 8 ][ 156 ],
   alphaCSR[ 8 ][ 157 ],
   alphaCSR[ 8 ][ 158 ],
   alphaCSR[ 8 ][ 159 ],
   alphaCSR[ 8 ][ 160 ],
   alphaCSR[ 8 ][ 161 ],
   alphaCSR[ 8 ][ 162 ],
   alphaCSR[ 8 ][ 163 ],
   alphaCSR[ 8 ][ 164 ],
   alphaCSR[ 8 ][ 165 ],
   alphaCSR[ 8 ][ 166 ],
   alphaCSR[ 8 ][ 167 ],
   alphaCSR[ 8 ][ 168 ],
   alphaCSR[ 8 ][ 169 ],
   alphaCSR[ 8 ][ 170 ],
   alphaCSR[ 8 ][ 171 ],
   alphaCSR[ 8 ][ 172 ],
   alphaCSR[ 8 ][ 173 ],
   alphaCSR[ 8 ][ 174 ],
   alphaCSR[ 8 ][ 175 ],
   alphaCSR[ 8 ][ 176 ],
   alphaCSR[ 8 ][ 177 ],
   alphaCSR[ 8 ][ 178 ],
   alphaCSR[ 8 ][ 179 ],
   alphaCSR[ 8 ][ 180 ],
   alphaCSR[ 8 ][ 181 ],
   alphaCSR[ 8 ][ 182 ],
   alphaCSR[ 8 ][ 183 ],
   alphaCSR[ 8 ][ 184 ],
   alphaCSR[ 8 ][ 185 ],
   alphaCSR[ 8 ][ 186 ],
   alphaCSR[ 8 ][ 187 ],
   alphaCSR[ 8 ][ 188 ],
   alphaCSR[ 8 ][ 189 ],
   alphaCSR[ 8 ][ 190 ],
   alphaCSR[ 8 ][ 191 ],
   alphaCSR[ 8 ][ 192 ],
   alphaCSR[ 8 ][ 193 ],
   alphaCSR[ 8 ][ 194 ],
   alphaCSR[ 8 ][ 195 ],
   alphaCSR[ 8 ][ 196 ],
   alphaCSR[ 8 ][ 197 ],
   alphaCSR[ 8 ][ 198 ],
   alphaCSR[ 8 ][ 199 ],
   alphaCSR[ 8 ][ 200 ],
   alphaCSR[ 8 ][ 201 ],
   alphaCSR[ 8 ][ 202 ],
   alphaCSR[ 8 ][ 203 ],
   alphaCSR[ 8 ][ 204 ],
   alphaCSR[ 8 ][ 205 ],
   alphaCSR[ 8 ][ 206 ],
   alphaCSR[ 8 ][ 207 ],
   alphaCSR[ 8 ][ 208 ],
   alphaCSR[ 8 ][ 209 ],
   alphaCSR[ 8 ][ 210 ],
   alphaCSR[ 8 ][ 211 ],
   alphaCSR[ 8 ][ 212 ],
   alphaCSR[ 8 ][ 213 ],
   alphaCSR[ 8 ][ 214 ],
   alphaCSR[ 8 ][ 215 ],
   alphaCSR[ 8 ][ 216 ],
   alphaCSR[ 8 ][ 217 ],
   alphaCSR[ 8 ][ 218 ],
   alphaCSR[ 8 ][ 219 ],
   alphaCSR[ 8 ][ 220 ],
   alphaCSR[ 8 ][ 221 ],
   alphaCSR[ 8 ][ 222 ],
   alphaCSR[ 8 ][ 223 ],
   alphaCSR[ 8 ][ 224 ],
   alphaCSR[ 8 ][ 225 ],
   alphaCSR[ 8 ][ 226 ],
   alphaCSR[ 8 ][ 227 ],
   alphaCSR[ 8 ][ 228 ],
   alphaCSR[ 8 ][ 229 ],
   alphaCSR[ 8 ][ 230 ],
   alphaCSR[ 8 ][ 231 ],
   alphaCSR[ 8 ][ 232 ],
   alphaCSR[ 8 ][ 233 ],
   alphaCSR[ 8 ][ 234 ],
   alphaCSR[ 8 ][ 235 ],
   alphaCSR[ 8 ][ 236 ],
   alphaCSR[ 8 ][ 237 ],
   alphaCSR[ 8 ][ 238 ],
   alphaCSR[ 8 ][ 239 ],
   alphaCSR[ 8 ][ 240 ],
   alphaCSR[ 8 ][ 241 ],
   alphaCSR[ 8 ][ 242 ],
   alphaCSR[ 8 ][ 243 ],
   alphaCSR[ 8 ][ 244 ],
   alphaCSR[ 8 ][ 245 ],
   alphaCSR[ 8 ][ 246 ],
   alphaCSR[ 8 ][ 247 ],
   alphaCSR[ 8 ][ 248 ],
   alphaCSR[ 8 ][ 249 ],
   alphaCSR[ 8 ][ 250 ],
   alphaCSR[ 8 ][ 251 ],
   alphaCSR[ 8 ][ 252 ],
   alphaCSR[ 8 ][ 253 ],
   alphaCSR[ 8 ][ 254 ],
   alphaCSR[ 8 ][ 255 ],
   alphaCSR[ 8 ][ 256 ],
   alphaCSR[ 8 ][ 257 ],
   alphaCSR[ 8 ][ 258 ],
   alphaCSR[ 8 ][ 259 ],
   alphaCSR[ 8 ][ 260 ],
   alphaCSR[ 8 ][ 261 ],
   alphaCSR[ 8 ][ 262 ],
   alphaCSR[ 8 ][ 263 ],
   alphaCSR[ 8 ][ 264 ],
   alphaCSR[ 8 ][ 265 ],
   alphaCSR[ 8 ][ 266 ],
   alphaCSR[ 8 ][ 267 ],
   alphaCSR[ 8 ][ 268 ],
   alphaCSR[ 8 ][ 269 ],
   alphaCSR[ 8 ][ 270 ],
   alphaCSR[ 8 ][ 271 ],
   alphaCSR[ 8 ][ 272 ],
   alphaCSR[ 8 ][ 273 ],
   alphaCSR[ 8 ][ 274 ],
   alphaCSR[ 8 ][ 275 ],
   alphaCSR[ 8 ][ 276 ],
   alphaCSR[ 8 ][ 277 ],
   alphaCSR[ 8 ][ 278 ],
   alphaCSR[ 8 ][ 279 ],
   alphaCSR[ 8 ][ 280 ],
   alphaCSR[ 8 ][ 281 ],
   alphaCSR[ 8 ][ 282 ],
   alphaCSR[ 8 ][ 283 ],
   alphaCSR[ 8 ][ 284 ],
   alphaCSR[ 8 ][ 285 ],
   alphaCSR[ 8 ][ 286 ],
   alphaCSR[ 8 ][ 287 ],
   alphaCSR[ 8 ][ 288 ],
   alphaCSR[ 8 ][ 289 ],
   alphaCSR[ 8 ][ 290 ],
   alphaCSR[ 8 ][ 291 ],
   alphaCSR[ 8 ][ 292 ],
   alphaCSR[ 8 ][ 293 ],
   alphaCSR[ 8 ][ 294 ],
   alphaCSR[ 8 ][ 295 ],
   alphaCSR[ 8 ][ 296 ],
   alphaCSR[ 8 ][ 297 ],
   alphaCSR[ 8 ][ 298 ],
   alphaCSR[ 8 ][ 299 ],
   alphaCSR[ 8 ][ 300 ],
   alphaCSR[ 8 ][ 301 ],
   alphaCSR[ 8 ][ 302 ],
   alphaCSR[ 8 ][ 303 ],
   alphaCSR[ 8 ][ 304 ],
   alphaCSR[ 8 ][ 305 ],
   alphaCSR[ 8 ][ 306 ],
   alphaCSR[ 8 ][ 307 ],
   alphaCSR[ 8 ][ 308 ],
   alphaCSR[ 8 ][ 309 ],
   alphaCSR[ 8 ][ 310 ],
   alphaCSR[ 8 ][ 311 ],
   alphaCSR[ 8 ][ 312 ],
   alphaCSR[ 8 ][ 313 ],
   alphaCSR[ 8 ][ 314 ],
   alphaCSR[ 8 ][ 315 ],
   alphaCSR[ 8 ][ 316 ],
   alphaCSR[ 8 ][ 317 ],
   alphaCSR[ 8 ][ 318 ],
   alphaCSR[ 8 ][ 319 ],
   alphaCSR[ 8 ][ 320 ],
   alphaCSR[ 8 ][ 321 ],
   alphaCSR[ 8 ][ 322 ],
   alphaCSR[ 8 ][ 323 ],
   alphaCSR[ 8 ][ 324 ],
   alphaCSR[ 8 ][ 325 ],
   alphaCSR[ 8 ][ 326 ],
   alphaCSR[ 8 ][ 327 ],
   alphaCSR[ 8 ][ 328 ],
   alphaCSR[ 8 ][ 329 ],
   alphaCSR[ 8 ][ 330 ],
   alphaCSR[ 8 ][ 331 ],
   alphaCSR[ 8 ][ 332 ],
   alphaCSR[ 8 ][ 333 ],
   alphaCSR[ 8 ][ 334 ],
   alphaCSR[ 8 ][ 335 ],
   alphaCSR[ 8 ][ 336 ],
   alphaCSR[ 8 ][ 337 ],
   alphaCSR[ 8 ][ 338 ],
   alphaCSR[ 8 ][ 339 ],
   alphaCSR[ 8 ][ 340 ],
   alphaCSR[ 8 ][ 341 ],
   alphaCSR[ 8 ][ 342 ],
   alphaCSR[ 8 ][ 343 ],
   alphaCSR[ 8 ][ 344 ],
   alphaCSR[ 8 ][ 345 ],
   alphaCSR[ 8 ][ 346 ],
   alphaCSR[ 8 ][ 347 ],
   alphaCSR[ 8 ][ 348 ],
   alphaCSR[ 8 ][ 349 ],
   alphaCSR[ 8 ][ 350 ],
   alphaCSR[ 8 ][ 351 ],
   alphaCSR[ 8 ][ 352 ],
   alphaCSR[ 8 ][ 353 ],
   alphaCSR[ 8 ][ 354 ],
   alphaCSR[ 8 ][ 355 ],
   alphaCSR[ 8 ][ 356 ],
   alphaCSR[ 8 ][ 357 ],
   alphaCSR[ 8 ][ 358 ],
   alphaCSR[ 8 ][ 359 ],
   alphaCSR[ 8 ][ 360 ],
   alphaCSR[ 8 ][ 361 ],
   alphaCSR[ 8 ][ 362 ],
   alphaCSR[ 8 ][ 363 ],
   alphaCSR[ 8 ][ 364 ],
   alphaCSR[ 8 ][ 365 ],
   alphaCSR[ 8 ][ 366 ],
   alphaCSR[ 8 ][ 367 ],
   alphaCSR[ 8 ][ 368 ],
   alphaCSR[ 8 ][ 369 ],
   alphaCSR[ 8 ][ 370 ],
   alphaCSR[ 8 ][ 371 ],
   alphaCSR[ 8 ][ 372 ],
   alphaCSR[ 8 ][ 373 ],
   alphaCSR[ 8 ][ 374 ],
   alphaCSR[ 8 ][ 375 ],
   alphaCSR[ 8 ][ 376 ],
   alphaCSR[ 8 ][ 377 ],
   alphaCSR[ 8 ][ 378 ],
   alphaCSR[ 8 ][ 379 ],
   alphaCSR[ 8 ][ 380 ],
   alphaCSR[ 8 ][ 381 ],
   alphaCSR[ 8 ][ 382 ],
   alphaCSR[ 8 ][ 383 ],
   alphaCSR[ 9 ][ 0 ],
   alphaCSR[ 9 ][ 1 ],
   alphaCSR[ 9 ][ 2 ],
   alphaCSR[ 9 ][ 3 ],
   alphaCSR[ 9 ][ 4 ],
   alphaCSR[ 9 ][ 5 ],
   alphaCSR[ 9 ][ 6 ],
   alphaCSR[ 9 ][ 7 ],
   alphaCSR[ 9 ][ 8 ],
   alphaCSR[ 9 ][ 9 ],
   alphaCSR[ 9 ][ 10 ],
   alphaCSR[ 9 ][ 11 ],
   alphaCSR[ 9 ][ 12 ],
   alphaCSR[ 9 ][ 13 ],
   alphaCSR[ 9 ][ 14 ],
   alphaCSR[ 9 ][ 15 ],
   alphaCSR[ 9 ][ 16 ],
   alphaCSR[ 9 ][ 17 ],
   alphaCSR[ 9 ][ 18 ],
   alphaCSR[ 9 ][ 19 ],
   alphaCSR[ 9 ][ 20 ],
   alphaCSR[ 9 ][ 21 ],
   alphaCSR[ 9 ][ 22 ],
   alphaCSR[ 9 ][ 23 ],
   alphaCSR[ 9 ][ 24 ],
   alphaCSR[ 9 ][ 25 ],
   alphaCSR[ 9 ][ 26 ],
   alphaCSR[ 9 ][ 27 ],
   alphaCSR[ 9 ][ 28 ],
   alphaCSR[ 9 ][ 29 ],
   alphaCSR[ 9 ][ 30 ],
   alphaCSR[ 9 ][ 31 ],
   alphaCSR[ 9 ][ 32 ],
   alphaCSR[ 9 ][ 33 ],
   alphaCSR[ 9 ][ 34 ],
   alphaCSR[ 9 ][ 35 ],
   alphaCSR[ 9 ][ 36 ],
   alphaCSR[ 9 ][ 37 ],
   alphaCSR[ 9 ][ 38 ],
   alphaCSR[ 9 ][ 39 ],
   alphaCSR[ 9 ][ 40 ],
   alphaCSR[ 9 ][ 41 ],
   alphaCSR[ 9 ][ 42 ],
   alphaCSR[ 9 ][ 43 ],
   alphaCSR[ 9 ][ 44 ],
   alphaCSR[ 9 ][ 45 ],
   alphaCSR[ 9 ][ 46 ],
   alphaCSR[ 9 ][ 47 ],
   alphaCSR[ 9 ][ 48 ],
   alphaCSR[ 9 ][ 49 ],
   alphaCSR[ 9 ][ 50 ],
   alphaCSR[ 9 ][ 51 ],
   alphaCSR[ 9 ][ 52 ],
   alphaCSR[ 9 ][ 53 ],
   alphaCSR[ 9 ][ 54 ],
   alphaCSR[ 9 ][ 55 ],
   alphaCSR[ 9 ][ 56 ],
   alphaCSR[ 9 ][ 57 ],
   alphaCSR[ 9 ][ 58 ],
   alphaCSR[ 9 ][ 59 ],
   alphaCSR[ 9 ][ 60 ],
   alphaCSR[ 9 ][ 61 ],
   alphaCSR[ 9 ][ 62 ],
   alphaCSR[ 9 ][ 63 ],
   alphaCSR[ 9 ][ 64 ],
   alphaCSR[ 9 ][ 65 ],
   alphaCSR[ 9 ][ 66 ],
   alphaCSR[ 9 ][ 67 ],
   alphaCSR[ 9 ][ 68 ],
   alphaCSR[ 9 ][ 69 ],
   alphaCSR[ 9 ][ 70 ],
   alphaCSR[ 9 ][ 71 ],
   alphaCSR[ 9 ][ 72 ],
   alphaCSR[ 9 ][ 73 ],
   alphaCSR[ 9 ][ 74 ],
   alphaCSR[ 9 ][ 75 ],
   alphaCSR[ 9 ][ 76 ],
   alphaCSR[ 9 ][ 77 ],
   alphaCSR[ 9 ][ 78 ],
   alphaCSR[ 9 ][ 79 ],
   alphaCSR[ 9 ][ 80 ],
   alphaCSR[ 9 ][ 81 ],
   alphaCSR[ 9 ][ 82 ],
   alphaCSR[ 9 ][ 83 ],
   alphaCSR[ 9 ][ 84 ],
   alphaCSR[ 9 ][ 85 ],
   alphaCSR[ 9 ][ 86 ],
   alphaCSR[ 9 ][ 87 ],
   alphaCSR[ 9 ][ 88 ],
   alphaCSR[ 9 ][ 89 ],
   alphaCSR[ 9 ][ 90 ],
   alphaCSR[ 9 ][ 91 ],
   alphaCSR[ 9 ][ 92 ],
   alphaCSR[ 9 ][ 93 ],
   alphaCSR[ 9 ][ 94 ],
   alphaCSR[ 9 ][ 95 ],
   alphaCSR[ 9 ][ 96 ],
   alphaCSR[ 9 ][ 97 ],
   alphaCSR[ 9 ][ 98 ],
   alphaCSR[ 9 ][ 99 ],
   alphaCSR[ 9 ][ 100 ],
   alphaCSR[ 9 ][ 101 ],
   alphaCSR[ 9 ][ 102 ],
   alphaCSR[ 9 ][ 103 ],
   alphaCSR[ 9 ][ 104 ],
   alphaCSR[ 9 ][ 105 ],
   alphaCSR[ 9 ][ 106 ],
   alphaCSR[ 9 ][ 107 ],
   alphaCSR[ 9 ][ 108 ],
   alphaCSR[ 9 ][ 109 ],
   alphaCSR[ 9 ][ 110 ],
   alphaCSR[ 9 ][ 111 ],
   alphaCSR[ 9 ][ 112 ],
   alphaCSR[ 9 ][ 113 ],
   alphaCSR[ 9 ][ 114 ],
   alphaCSR[ 9 ][ 115 ],
   alphaCSR[ 9 ][ 116 ],
   alphaCSR[ 9 ][ 117 ],
   alphaCSR[ 9 ][ 118 ],
   alphaCSR[ 9 ][ 119 ],
   alphaCSR[ 9 ][ 120 ],
   alphaCSR[ 9 ][ 121 ],
   alphaCSR[ 9 ][ 122 ],
   alphaCSR[ 9 ][ 123 ],
   alphaCSR[ 9 ][ 124 ],
   alphaCSR[ 9 ][ 125 ],
   alphaCSR[ 9 ][ 126 ],
   alphaCSR[ 9 ][ 127 ],
   alphaCSR[ 9 ][ 128 ],
   alphaCSR[ 9 ][ 129 ],
   alphaCSR[ 9 ][ 130 ],
   alphaCSR[ 9 ][ 131 ],
   alphaCSR[ 9 ][ 132 ],
   alphaCSR[ 9 ][ 133 ],
   alphaCSR[ 9 ][ 134 ],
   alphaCSR[ 9 ][ 135 ],
   alphaCSR[ 9 ][ 136 ],
   alphaCSR[ 9 ][ 137 ],
   alphaCSR[ 9 ][ 138 ],
   alphaCSR[ 9 ][ 139 ],
   alphaCSR[ 9 ][ 140 ],
   alphaCSR[ 9 ][ 141 ],
   alphaCSR[ 9 ][ 142 ],
   alphaCSR[ 9 ][ 143 ],
   alphaCSR[ 9 ][ 144 ],
   alphaCSR[ 9 ][ 145 ],
   alphaCSR[ 9 ][ 146 ],
   alphaCSR[ 9 ][ 147 ],
   alphaCSR[ 9 ][ 148 ],
   alphaCSR[ 9 ][ 149 ],
   alphaCSR[ 9 ][ 150 ],
   alphaCSR[ 9 ][ 151 ],
   alphaCSR[ 9 ][ 152 ],
   alphaCSR[ 9 ][ 153 ],
   alphaCSR[ 9 ][ 154 ],
   alphaCSR[ 9 ][ 155 ],
   alphaCSR[ 9 ][ 156 ],
   alphaCSR[ 9 ][ 157 ],
   alphaCSR[ 9 ][ 158 ],
   alphaCSR[ 9 ][ 159 ],
   alphaCSR[ 9 ][ 160 ],
   alphaCSR[ 9 ][ 161 ],
   alphaCSR[ 9 ][ 162 ],
   alphaCSR[ 9 ][ 163 ],
   alphaCSR[ 9 ][ 164 ],
   alphaCSR[ 9 ][ 165 ],
   alphaCSR[ 9 ][ 166 ],
   alphaCSR[ 9 ][ 167 ],
   alphaCSR[ 9 ][ 168 ],
   alphaCSR[ 9 ][ 169 ],
   alphaCSR[ 9 ][ 170 ],
   alphaCSR[ 9 ][ 171 ],
   alphaCSR[ 9 ][ 172 ],
   alphaCSR[ 9 ][ 173 ],
   alphaCSR[ 9 ][ 174 ],
   alphaCSR[ 9 ][ 175 ],
   alphaCSR[ 9 ][ 176 ],
   alphaCSR[ 9 ][ 177 ],
   alphaCSR[ 9 ][ 178 ],
   alphaCSR[ 9 ][ 179 ],
   alphaCSR[ 9 ][ 180 ],
   alphaCSR[ 9 ][ 181 ],
   alphaCSR[ 9 ][ 182 ],
   alphaCSR[ 9 ][ 183 ],
   alphaCSR[ 9 ][ 184 ],
   alphaCSR[ 9 ][ 185 ],
   alphaCSR[ 9 ][ 186 ],
   alphaCSR[ 9 ][ 187 ],
   alphaCSR[ 9 ][ 188 ],
   alphaCSR[ 9 ][ 189 ],
   alphaCSR[ 9 ][ 190 ],
   alphaCSR[ 9 ][ 191 ],
   alphaCSR[ 9 ][ 192 ],
   alphaCSR[ 9 ][ 193 ],
   alphaCSR[ 9 ][ 194 ],
   alphaCSR[ 9 ][ 195 ],
   alphaCSR[ 9 ][ 196 ],
   alphaCSR[ 9 ][ 197 ],
   alphaCSR[ 9 ][ 198 ],
   alphaCSR[ 9 ][ 199 ],
   alphaCSR[ 9 ][ 200 ],
   alphaCSR[ 9 ][ 201 ],
   alphaCSR[ 9 ][ 202 ],
   alphaCSR[ 9 ][ 203 ],
   alphaCSR[ 9 ][ 204 ],
   alphaCSR[ 9 ][ 205 ],
   alphaCSR[ 9 ][ 206 ],
   alphaCSR[ 9 ][ 207 ],
   alphaCSR[ 9 ][ 208 ],
   alphaCSR[ 9 ][ 209 ],
   alphaCSR[ 9 ][ 210 ],
   alphaCSR[ 9 ][ 211 ],
   alphaCSR[ 9 ][ 212 ],
   alphaCSR[ 9 ][ 213 ],
   alphaCSR[ 9 ][ 214 ],
   alphaCSR[ 9 ][ 215 ],
   alphaCSR[ 9 ][ 216 ],
   alphaCSR[ 9 ][ 217 ],
   alphaCSR[ 9 ][ 218 ],
   alphaCSR[ 9 ][ 219 ],
   alphaCSR[ 9 ][ 220 ],
   alphaCSR[ 9 ][ 221 ],
   alphaCSR[ 9 ][ 222 ],
   alphaCSR[ 9 ][ 223 ],
   alphaCSR[ 9 ][ 224 ],
   alphaCSR[ 9 ][ 225 ],
   alphaCSR[ 9 ][ 226 ],
   alphaCSR[ 9 ][ 227 ],
   alphaCSR[ 9 ][ 228 ],
   alphaCSR[ 9 ][ 229 ],
   alphaCSR[ 9 ][ 230 ],
   alphaCSR[ 9 ][ 231 ],
   alphaCSR[ 9 ][ 232 ],
   alphaCSR[ 9 ][ 233 ],
   alphaCSR[ 9 ][ 234 ],
   alphaCSR[ 9 ][ 235 ],
   alphaCSR[ 9 ][ 236 ],
   alphaCSR[ 9 ][ 237 ],
   alphaCSR[ 9 ][ 238 ],
   alphaCSR[ 9 ][ 239 ],
   alphaCSR[ 9 ][ 240 ],
   alphaCSR[ 9 ][ 241 ],
   alphaCSR[ 9 ][ 242 ],
   alphaCSR[ 9 ][ 243 ],
   alphaCSR[ 9 ][ 244 ],
   alphaCSR[ 9 ][ 245 ],
   alphaCSR[ 9 ][ 246 ],
   alphaCSR[ 9 ][ 247 ],
   alphaCSR[ 9 ][ 248 ],
   alphaCSR[ 9 ][ 249 ],
   alphaCSR[ 9 ][ 250 ],
   alphaCSR[ 9 ][ 251 ],
   alphaCSR[ 9 ][ 252 ],
   alphaCSR[ 9 ][ 253 ],
   alphaCSR[ 9 ][ 254 ],
   alphaCSR[ 9 ][ 255 ],
   alphaCSR[ 9 ][ 256 ],
   alphaCSR[ 9 ][ 257 ],
   alphaCSR[ 9 ][ 258 ],
   alphaCSR[ 9 ][ 259 ],
   alphaCSR[ 9 ][ 260 ],
   alphaCSR[ 9 ][ 261 ],
   alphaCSR[ 9 ][ 262 ],
   alphaCSR[ 9 ][ 263 ],
   alphaCSR[ 9 ][ 264 ],
   alphaCSR[ 9 ][ 265 ],
   alphaCSR[ 9 ][ 266 ],
   alphaCSR[ 9 ][ 267 ],
   alphaCSR[ 9 ][ 268 ],
   alphaCSR[ 9 ][ 269 ],
   alphaCSR[ 9 ][ 270 ],
   alphaCSR[ 9 ][ 271 ],
   alphaCSR[ 9 ][ 272 ],
   alphaCSR[ 9 ][ 273 ],
   alphaCSR[ 9 ][ 274 ],
   alphaCSR[ 9 ][ 275 ],
   alphaCSR[ 9 ][ 276 ],
   alphaCSR[ 9 ][ 277 ],
   alphaCSR[ 9 ][ 278 ],
   alphaCSR[ 9 ][ 279 ],
   alphaCSR[ 9 ][ 280 ],
   alphaCSR[ 9 ][ 281 ],
   alphaCSR[ 9 ][ 282 ],
   alphaCSR[ 9 ][ 283 ],
   alphaCSR[ 9 ][ 284 ],
   alphaCSR[ 9 ][ 285 ],
   alphaCSR[ 9 ][ 286 ],
   alphaCSR[ 9 ][ 287 ],
   alphaCSR[ 9 ][ 288 ],
   alphaCSR[ 9 ][ 289 ],
   alphaCSR[ 9 ][ 290 ],
   alphaCSR[ 9 ][ 291 ],
   alphaCSR[ 9 ][ 292 ],
   alphaCSR[ 9 ][ 293 ],
   alphaCSR[ 9 ][ 294 ],
   alphaCSR[ 9 ][ 295 ],
   alphaCSR[ 9 ][ 296 ],
   alphaCSR[ 9 ][ 297 ],
   alphaCSR[ 9 ][ 298 ],
   alphaCSR[ 9 ][ 299 ],
   alphaCSR[ 9 ][ 300 ],
   alphaCSR[ 9 ][ 301 ],
   alphaCSR[ 9 ][ 302 ],
   alphaCSR[ 9 ][ 303 ],
   alphaCSR[ 9 ][ 304 ],
   alphaCSR[ 9 ][ 305 ],
   alphaCSR[ 9 ][ 306 ],
   alphaCSR[ 9 ][ 307 ],
   alphaCSR[ 9 ][ 308 ],
   alphaCSR[ 9 ][ 309 ],
   alphaCSR[ 9 ][ 310 ],
   alphaCSR[ 9 ][ 311 ],
   alphaCSR[ 9 ][ 312 ],
   alphaCSR[ 9 ][ 313 ],
   alphaCSR[ 9 ][ 314 ],
   alphaCSR[ 9 ][ 315 ],
   alphaCSR[ 9 ][ 316 ],
   alphaCSR[ 9 ][ 317 ],
   alphaCSR[ 9 ][ 318 ],
   alphaCSR[ 9 ][ 319 ],
   alphaCSR[ 9 ][ 320 ],
   alphaCSR[ 9 ][ 321 ],
   alphaCSR[ 9 ][ 322 ],
   alphaCSR[ 9 ][ 323 ],
   alphaCSR[ 9 ][ 324 ],
   alphaCSR[ 9 ][ 325 ],
   alphaCSR[ 9 ][ 326 ],
   alphaCSR[ 9 ][ 327 ],
   alphaCSR[ 9 ][ 328 ],
   alphaCSR[ 9 ][ 329 ],
   alphaCSR[ 9 ][ 330 ],
   alphaCSR[ 9 ][ 331 ],
   alphaCSR[ 9 ][ 332 ],
   alphaCSR[ 9 ][ 333 ],
   alphaCSR[ 9 ][ 334 ],
   alphaCSR[ 9 ][ 335 ],
   alphaCSR[ 9 ][ 336 ],
   alphaCSR[ 9 ][ 337 ],
   alphaCSR[ 9 ][ 338 ],
   alphaCSR[ 9 ][ 339 ],
   alphaCSR[ 9 ][ 340 ],
   alphaCSR[ 9 ][ 341 ],
   alphaCSR[ 9 ][ 342 ],
   alphaCSR[ 9 ][ 343 ],
   alphaCSR[ 9 ][ 344 ],
   alphaCSR[ 9 ][ 345 ],
   alphaCSR[ 9 ][ 346 ],
   alphaCSR[ 9 ][ 347 ],
   alphaCSR[ 9 ][ 348 ],
   alphaCSR[ 9 ][ 349 ],
   alphaCSR[ 9 ][ 350 ],
   alphaCSR[ 9 ][ 351 ],
   alphaCSR[ 9 ][ 352 ],
   alphaCSR[ 9 ][ 353 ],
   alphaCSR[ 9 ][ 354 ],
   alphaCSR[ 9 ][ 355 ],
   alphaCSR[ 9 ][ 356 ],
   alphaCSR[ 9 ][ 357 ],
   alphaCSR[ 9 ][ 358 ],
   alphaCSR[ 9 ][ 359 ],
   alphaCSR[ 9 ][ 360 ],
   alphaCSR[ 9 ][ 361 ],
   alphaCSR[ 9 ][ 362 ],
   alphaCSR[ 9 ][ 363 ],
   alphaCSR[ 9 ][ 364 ],
   alphaCSR[ 9 ][ 365 ],
   alphaCSR[ 9 ][ 366 ],
   alphaCSR[ 9 ][ 367 ],
   alphaCSR[ 9 ][ 368 ],
   alphaCSR[ 9 ][ 369 ],
   alphaCSR[ 9 ][ 370 ],
   alphaCSR[ 9 ][ 371 ],
   alphaCSR[ 9 ][ 372 ],
   alphaCSR[ 9 ][ 373 ],
   alphaCSR[ 9 ][ 374 ],
   alphaCSR[ 9 ][ 375 ],
   alphaCSR[ 9 ][ 376 ],
   alphaCSR[ 9 ][ 377 ],
   alphaCSR[ 9 ][ 378 ],
   alphaCSR[ 9 ][ 379 ],
   alphaCSR[ 9 ][ 380 ],
   alphaCSR[ 9 ][ 381 ],
   alphaCSR[ 9 ][ 382 ],
   alphaCSR[ 9 ][ 383 ],
   alphaCSR[ 10 ][ 0 ],
   alphaCSR[ 10 ][ 1 ],
   alphaCSR[ 10 ][ 2 ],
   alphaCSR[ 10 ][ 3 ],
   alphaCSR[ 10 ][ 4 ],
   alphaCSR[ 10 ][ 5 ],
   alphaCSR[ 10 ][ 6 ],
   alphaCSR[ 10 ][ 7 ],
   alphaCSR[ 10 ][ 8 ],
   alphaCSR[ 10 ][ 9 ],
   alphaCSR[ 10 ][ 10 ],
   alphaCSR[ 10 ][ 11 ],
   alphaCSR[ 10 ][ 12 ],
   alphaCSR[ 10 ][ 13 ],
   alphaCSR[ 10 ][ 14 ],
   alphaCSR[ 10 ][ 15 ],
   alphaCSR[ 10 ][ 16 ],
   alphaCSR[ 10 ][ 17 ],
   alphaCSR[ 10 ][ 18 ],
   alphaCSR[ 10 ][ 19 ],
   alphaCSR[ 10 ][ 20 ],
   alphaCSR[ 10 ][ 21 ],
   alphaCSR[ 10 ][ 22 ],
   alphaCSR[ 10 ][ 23 ],
   alphaCSR[ 10 ][ 24 ],
   alphaCSR[ 10 ][ 25 ],
   alphaCSR[ 10 ][ 26 ],
   alphaCSR[ 10 ][ 27 ],
   alphaCSR[ 10 ][ 28 ],
   alphaCSR[ 10 ][ 29 ],
   alphaCSR[ 10 ][ 30 ],
   alphaCSR[ 10 ][ 31 ],
   alphaCSR[ 10 ][ 32 ],
   alphaCSR[ 10 ][ 33 ],
   alphaCSR[ 10 ][ 34 ],
   alphaCSR[ 10 ][ 35 ],
   alphaCSR[ 10 ][ 36 ],
   alphaCSR[ 10 ][ 37 ],
   alphaCSR[ 10 ][ 38 ],
   alphaCSR[ 10 ][ 39 ],
   alphaCSR[ 10 ][ 40 ],
   alphaCSR[ 10 ][ 41 ],
   alphaCSR[ 10 ][ 42 ],
   alphaCSR[ 10 ][ 43 ],
   alphaCSR[ 10 ][ 44 ],
   alphaCSR[ 10 ][ 45 ],
   alphaCSR[ 10 ][ 46 ],
   alphaCSR[ 10 ][ 47 ],
   alphaCSR[ 10 ][ 48 ],
   alphaCSR[ 10 ][ 49 ],
   alphaCSR[ 10 ][ 50 ],
   alphaCSR[ 10 ][ 51 ],
   alphaCSR[ 10 ][ 52 ],
   alphaCSR[ 10 ][ 53 ],
   alphaCSR[ 10 ][ 54 ],
   alphaCSR[ 10 ][ 55 ],
   alphaCSR[ 10 ][ 56 ],
   alphaCSR[ 10 ][ 57 ],
   alphaCSR[ 10 ][ 58 ],
   alphaCSR[ 10 ][ 59 ],
   alphaCSR[ 10 ][ 60 ],
   alphaCSR[ 10 ][ 61 ],
   alphaCSR[ 10 ][ 62 ],
   alphaCSR[ 10 ][ 63 ],
   alphaCSR[ 10 ][ 64 ],
   alphaCSR[ 10 ][ 65 ],
   alphaCSR[ 10 ][ 66 ],
   alphaCSR[ 10 ][ 67 ],
   alphaCSR[ 10 ][ 68 ],
   alphaCSR[ 10 ][ 69 ],
   alphaCSR[ 10 ][ 70 ],
   alphaCSR[ 10 ][ 71 ],
   alphaCSR[ 10 ][ 72 ],
   alphaCSR[ 10 ][ 73 ],
   alphaCSR[ 10 ][ 74 ],
   alphaCSR[ 10 ][ 75 ],
   alphaCSR[ 10 ][ 76 ],
   alphaCSR[ 10 ][ 77 ],
   alphaCSR[ 10 ][ 78 ],
   alphaCSR[ 10 ][ 79 ],
   alphaCSR[ 10 ][ 80 ],
   alphaCSR[ 10 ][ 81 ],
   alphaCSR[ 10 ][ 82 ],
   alphaCSR[ 10 ][ 83 ],
   alphaCSR[ 10 ][ 84 ],
   alphaCSR[ 10 ][ 85 ],
   alphaCSR[ 10 ][ 86 ],
   alphaCSR[ 10 ][ 87 ],
   alphaCSR[ 10 ][ 88 ],
   alphaCSR[ 10 ][ 89 ],
   alphaCSR[ 10 ][ 90 ],
   alphaCSR[ 10 ][ 91 ],
   alphaCSR[ 10 ][ 92 ],
   alphaCSR[ 10 ][ 93 ],
   alphaCSR[ 10 ][ 94 ],
   alphaCSR[ 10 ][ 95 ],
   alphaCSR[ 10 ][ 96 ],
   alphaCSR[ 10 ][ 97 ],
   alphaCSR[ 10 ][ 98 ],
   alphaCSR[ 10 ][ 99 ],
   alphaCSR[ 10 ][ 100 ],
   alphaCSR[ 10 ][ 101 ],
   alphaCSR[ 10 ][ 102 ],
   alphaCSR[ 10 ][ 103 ],
   alphaCSR[ 10 ][ 104 ],
   alphaCSR[ 10 ][ 105 ],
   alphaCSR[ 10 ][ 106 ],
   alphaCSR[ 10 ][ 107 ],
   alphaCSR[ 10 ][ 108 ],
   alphaCSR[ 10 ][ 109 ],
   alphaCSR[ 10 ][ 110 ],
   alphaCSR[ 10 ][ 111 ],
   alphaCSR[ 10 ][ 112 ],
   alphaCSR[ 10 ][ 113 ],
   alphaCSR[ 10 ][ 114 ],
   alphaCSR[ 10 ][ 115 ],
   alphaCSR[ 10 ][ 116 ],
   alphaCSR[ 10 ][ 117 ],
   alphaCSR[ 10 ][ 118 ],
   alphaCSR[ 10 ][ 119 ],
   alphaCSR[ 10 ][ 120 ],
   alphaCSR[ 10 ][ 121 ],
   alphaCSR[ 10 ][ 122 ],
   alphaCSR[ 10 ][ 123 ],
   alphaCSR[ 10 ][ 124 ],
   alphaCSR[ 10 ][ 125 ],
   alphaCSR[ 10 ][ 126 ],
   alphaCSR[ 10 ][ 127 ],
   alphaCSR[ 10 ][ 128 ],
   alphaCSR[ 10 ][ 129 ],
   alphaCSR[ 10 ][ 130 ],
   alphaCSR[ 10 ][ 131 ],
   alphaCSR[ 10 ][ 132 ],
   alphaCSR[ 10 ][ 133 ],
   alphaCSR[ 10 ][ 134 ],
   alphaCSR[ 10 ][ 135 ],
   alphaCSR[ 10 ][ 136 ],
   alphaCSR[ 10 ][ 137 ],
   alphaCSR[ 10 ][ 138 ],
   alphaCSR[ 10 ][ 139 ],
   alphaCSR[ 10 ][ 140 ],
   alphaCSR[ 10 ][ 141 ],
   alphaCSR[ 10 ][ 142 ],
   alphaCSR[ 10 ][ 143 ],
   alphaCSR[ 10 ][ 144 ],
   alphaCSR[ 10 ][ 145 ],
   alphaCSR[ 10 ][ 146 ],
   alphaCSR[ 10 ][ 147 ],
   alphaCSR[ 10 ][ 148 ],
   alphaCSR[ 10 ][ 149 ],
   alphaCSR[ 10 ][ 150 ],
   alphaCSR[ 10 ][ 151 ],
   alphaCSR[ 10 ][ 152 ],
   alphaCSR[ 10 ][ 153 ],
   alphaCSR[ 10 ][ 154 ],
   alphaCSR[ 10 ][ 155 ],
   alphaCSR[ 10 ][ 156 ],
   alphaCSR[ 10 ][ 157 ],
   alphaCSR[ 10 ][ 158 ],
   alphaCSR[ 10 ][ 159 ],
   alphaCSR[ 10 ][ 160 ],
   alphaCSR[ 10 ][ 161 ],
   alphaCSR[ 10 ][ 162 ],
   alphaCSR[ 10 ][ 163 ],
   alphaCSR[ 10 ][ 164 ],
   alphaCSR[ 10 ][ 165 ],
   alphaCSR[ 10 ][ 166 ],
   alphaCSR[ 10 ][ 167 ],
   alphaCSR[ 10 ][ 168 ],
   alphaCSR[ 10 ][ 169 ],
   alphaCSR[ 10 ][ 170 ],
   alphaCSR[ 10 ][ 171 ],
   alphaCSR[ 10 ][ 172 ],
   alphaCSR[ 10 ][ 173 ],
   alphaCSR[ 10 ][ 174 ],
   alphaCSR[ 10 ][ 175 ],
   alphaCSR[ 10 ][ 176 ],
   alphaCSR[ 10 ][ 177 ],
   alphaCSR[ 10 ][ 178 ],
   alphaCSR[ 10 ][ 179 ],
   alphaCSR[ 10 ][ 180 ],
   alphaCSR[ 10 ][ 181 ],
   alphaCSR[ 10 ][ 182 ],
   alphaCSR[ 10 ][ 183 ],
   alphaCSR[ 10 ][ 184 ],
   alphaCSR[ 10 ][ 185 ],
   alphaCSR[ 10 ][ 186 ],
   alphaCSR[ 10 ][ 187 ],
   alphaCSR[ 10 ][ 188 ],
   alphaCSR[ 10 ][ 189 ],
   alphaCSR[ 10 ][ 190 ],
   alphaCSR[ 10 ][ 191 ],
   alphaCSR[ 10 ][ 192 ],
   alphaCSR[ 10 ][ 193 ],
   alphaCSR[ 10 ][ 194 ],
   alphaCSR[ 10 ][ 195 ],
   alphaCSR[ 10 ][ 196 ],
   alphaCSR[ 10 ][ 197 ],
   alphaCSR[ 10 ][ 198 ],
   alphaCSR[ 10 ][ 199 ],
   alphaCSR[ 10 ][ 200 ],
   alphaCSR[ 10 ][ 201 ],
   alphaCSR[ 10 ][ 202 ],
   alphaCSR[ 10 ][ 203 ],
   alphaCSR[ 10 ][ 204 ],
   alphaCSR[ 10 ][ 205 ],
   alphaCSR[ 10 ][ 206 ],
   alphaCSR[ 10 ][ 207 ],
   alphaCSR[ 10 ][ 208 ],
   alphaCSR[ 10 ][ 209 ],
   alphaCSR[ 10 ][ 210 ],
   alphaCSR[ 10 ][ 211 ],
   alphaCSR[ 10 ][ 212 ],
   alphaCSR[ 10 ][ 213 ],
   alphaCSR[ 10 ][ 214 ],
   alphaCSR[ 10 ][ 215 ],
   alphaCSR[ 10 ][ 216 ],
   alphaCSR[ 10 ][ 217 ],
   alphaCSR[ 10 ][ 218 ],
   alphaCSR[ 10 ][ 219 ],
   alphaCSR[ 10 ][ 220 ],
   alphaCSR[ 10 ][ 221 ],
   alphaCSR[ 10 ][ 222 ],
   alphaCSR[ 10 ][ 223 ],
   alphaCSR[ 10 ][ 224 ],
   alphaCSR[ 10 ][ 225 ],
   alphaCSR[ 10 ][ 226 ],
   alphaCSR[ 10 ][ 227 ],
   alphaCSR[ 10 ][ 228 ],
   alphaCSR[ 10 ][ 229 ],
   alphaCSR[ 10 ][ 230 ],
   alphaCSR[ 10 ][ 231 ],
   alphaCSR[ 10 ][ 232 ],
   alphaCSR[ 10 ][ 233 ],
   alphaCSR[ 10 ][ 234 ],
   alphaCSR[ 10 ][ 235 ],
   alphaCSR[ 10 ][ 236 ],
   alphaCSR[ 10 ][ 237 ],
   alphaCSR[ 10 ][ 238 ],
   alphaCSR[ 10 ][ 239 ],
   alphaCSR[ 10 ][ 240 ],
   alphaCSR[ 10 ][ 241 ],
   alphaCSR[ 10 ][ 242 ],
   alphaCSR[ 10 ][ 243 ],
   alphaCSR[ 10 ][ 244 ],
   alphaCSR[ 10 ][ 245 ],
   alphaCSR[ 10 ][ 246 ],
   alphaCSR[ 10 ][ 247 ],
   alphaCSR[ 10 ][ 248 ],
   alphaCSR[ 10 ][ 249 ],
   alphaCSR[ 10 ][ 250 ],
   alphaCSR[ 10 ][ 251 ],
   alphaCSR[ 10 ][ 252 ],
   alphaCSR[ 10 ][ 253 ],
   alphaCSR[ 10 ][ 254 ],
   alphaCSR[ 10 ][ 255 ],
   alphaCSR[ 10 ][ 256 ],
   alphaCSR[ 10 ][ 257 ],
   alphaCSR[ 10 ][ 258 ],
   alphaCSR[ 10 ][ 259 ],
   alphaCSR[ 10 ][ 260 ],
   alphaCSR[ 10 ][ 261 ],
   alphaCSR[ 10 ][ 262 ],
   alphaCSR[ 10 ][ 263 ],
   alphaCSR[ 10 ][ 264 ],
   alphaCSR[ 10 ][ 265 ],
   alphaCSR[ 10 ][ 266 ],
   alphaCSR[ 10 ][ 267 ],
   alphaCSR[ 10 ][ 268 ],
   alphaCSR[ 10 ][ 269 ],
   alphaCSR[ 10 ][ 270 ],
   alphaCSR[ 10 ][ 271 ],
   alphaCSR[ 10 ][ 272 ],
   alphaCSR[ 10 ][ 273 ],
   alphaCSR[ 10 ][ 274 ],
   alphaCSR[ 10 ][ 275 ],
   alphaCSR[ 10 ][ 276 ],
   alphaCSR[ 10 ][ 277 ],
   alphaCSR[ 10 ][ 278 ],
   alphaCSR[ 10 ][ 279 ],
   alphaCSR[ 10 ][ 280 ],
   alphaCSR[ 10 ][ 281 ],
   alphaCSR[ 10 ][ 282 ],
   alphaCSR[ 10 ][ 283 ],
   alphaCSR[ 10 ][ 284 ],
   alphaCSR[ 10 ][ 285 ],
   alphaCSR[ 10 ][ 286 ],
   alphaCSR[ 10 ][ 287 ],
   alphaCSR[ 10 ][ 288 ],
   alphaCSR[ 10 ][ 289 ],
   alphaCSR[ 10 ][ 290 ],
   alphaCSR[ 10 ][ 291 ],
   alphaCSR[ 10 ][ 292 ],
   alphaCSR[ 10 ][ 293 ],
   alphaCSR[ 10 ][ 294 ],
   alphaCSR[ 10 ][ 295 ],
   alphaCSR[ 10 ][ 296 ],
   alphaCSR[ 10 ][ 297 ],
   alphaCSR[ 10 ][ 298 ],
   alphaCSR[ 10 ][ 299 ],
   alphaCSR[ 10 ][ 300 ],
   alphaCSR[ 10 ][ 301 ],
   alphaCSR[ 10 ][ 302 ],
   alphaCSR[ 10 ][ 303 ],
   alphaCSR[ 10 ][ 304 ],
   alphaCSR[ 10 ][ 305 ],
   alphaCSR[ 10 ][ 306 ],
   alphaCSR[ 10 ][ 307 ],
   alphaCSR[ 10 ][ 308 ],
   alphaCSR[ 10 ][ 309 ],
   alphaCSR[ 10 ][ 310 ],
   alphaCSR[ 10 ][ 311 ],
   alphaCSR[ 10 ][ 312 ],
   alphaCSR[ 10 ][ 313 ],
   alphaCSR[ 10 ][ 314 ],
   alphaCSR[ 10 ][ 315 ],
   alphaCSR[ 10 ][ 316 ],
   alphaCSR[ 10 ][ 317 ],
   alphaCSR[ 10 ][ 318 ],
   alphaCSR[ 10 ][ 319 ],
   alphaCSR[ 10 ][ 320 ],
   alphaCSR[ 10 ][ 321 ],
   alphaCSR[ 10 ][ 322 ],
   alphaCSR[ 10 ][ 323 ],
   alphaCSR[ 10 ][ 324 ],
   alphaCSR[ 10 ][ 325 ],
   alphaCSR[ 10 ][ 326 ],
   alphaCSR[ 10 ][ 327 ],
   alphaCSR[ 10 ][ 328 ],
   alphaCSR[ 10 ][ 329 ],
   alphaCSR[ 10 ][ 330 ],
   alphaCSR[ 10 ][ 331 ],
   alphaCSR[ 10 ][ 332 ],
   alphaCSR[ 10 ][ 333 ],
   alphaCSR[ 10 ][ 334 ],
   alphaCSR[ 10 ][ 335 ],
   alphaCSR[ 10 ][ 336 ],
   alphaCSR[ 10 ][ 337 ],
   alphaCSR[ 10 ][ 338 ],
   alphaCSR[ 10 ][ 339 ],
   alphaCSR[ 10 ][ 340 ],
   alphaCSR[ 10 ][ 341 ],
   alphaCSR[ 10 ][ 342 ],
   alphaCSR[ 10 ][ 343 ],
   alphaCSR[ 10 ][ 344 ],
   alphaCSR[ 10 ][ 345 ],
   alphaCSR[ 10 ][ 346 ],
   alphaCSR[ 10 ][ 347 ],
   alphaCSR[ 10 ][ 348 ],
   alphaCSR[ 10 ][ 349 ],
   alphaCSR[ 10 ][ 350 ],
   alphaCSR[ 10 ][ 351 ],
   alphaCSR[ 10 ][ 352 ],
   alphaCSR[ 10 ][ 353 ],
   alphaCSR[ 10 ][ 354 ],
   alphaCSR[ 10 ][ 355 ],
   alphaCSR[ 10 ][ 356 ],
   alphaCSR[ 10 ][ 357 ],
   alphaCSR[ 10 ][ 358 ],
   alphaCSR[ 10 ][ 359 ],
   alphaCSR[ 10 ][ 360 ],
   alphaCSR[ 10 ][ 361 ],
   alphaCSR[ 10 ][ 362 ],
   alphaCSR[ 10 ][ 363 ],
   alphaCSR[ 10 ][ 364 ],
   alphaCSR[ 10 ][ 365 ],
   alphaCSR[ 10 ][ 366 ],
   alphaCSR[ 10 ][ 367 ],
   alphaCSR[ 10 ][ 368 ],
   alphaCSR[ 10 ][ 369 ],
   alphaCSR[ 10 ][ 370 ],
   alphaCSR[ 10 ][ 371 ],
   alphaCSR[ 10 ][ 372 ],
   alphaCSR[ 10 ][ 373 ],
   alphaCSR[ 10 ][ 374 ],
   alphaCSR[ 10 ][ 375 ],
   alphaCSR[ 10 ][ 376 ],
   alphaCSR[ 10 ][ 377 ],
   alphaCSR[ 10 ][ 378 ],
   alphaCSR[ 10 ][ 379 ],
   alphaCSR[ 10 ][ 380 ],
   alphaCSR[ 10 ][ 381 ],
   alphaCSR[ 10 ][ 382 ],
   alphaCSR[ 10 ][ 383 ],
   alphaCSR[ 11 ][ 0 ],
   alphaCSR[ 11 ][ 1 ],
   alphaCSR[ 11 ][ 2 ],
   alphaCSR[ 11 ][ 3 ],
   alphaCSR[ 11 ][ 4 ],
   alphaCSR[ 11 ][ 5 ],
   alphaCSR[ 11 ][ 6 ],
   alphaCSR[ 11 ][ 7 ],
   alphaCSR[ 11 ][ 8 ],
   alphaCSR[ 11 ][ 9 ],
   alphaCSR[ 11 ][ 10 ],
   alphaCSR[ 11 ][ 11 ],
   alphaCSR[ 11 ][ 12 ],
   alphaCSR[ 11 ][ 13 ],
   alphaCSR[ 11 ][ 14 ],
   alphaCSR[ 11 ][ 15 ],
   alphaCSR[ 11 ][ 16 ],
   alphaCSR[ 11 ][ 17 ],
   alphaCSR[ 11 ][ 18 ],
   alphaCSR[ 11 ][ 19 ],
   alphaCSR[ 11 ][ 20 ],
   alphaCSR[ 11 ][ 21 ],
   alphaCSR[ 11 ][ 22 ],
   alphaCSR[ 11 ][ 23 ],
   alphaCSR[ 11 ][ 24 ],
   alphaCSR[ 11 ][ 25 ],
   alphaCSR[ 11 ][ 26 ],
   alphaCSR[ 11 ][ 27 ],
   alphaCSR[ 11 ][ 28 ],
   alphaCSR[ 11 ][ 29 ],
   alphaCSR[ 11 ][ 30 ],
   alphaCSR[ 11 ][ 31 ],
   alphaCSR[ 11 ][ 32 ],
   alphaCSR[ 11 ][ 33 ],
   alphaCSR[ 11 ][ 34 ],
   alphaCSR[ 11 ][ 35 ],
   alphaCSR[ 11 ][ 36 ],
   alphaCSR[ 11 ][ 37 ],
   alphaCSR[ 11 ][ 38 ],
   alphaCSR[ 11 ][ 39 ],
   alphaCSR[ 11 ][ 40 ],
   alphaCSR[ 11 ][ 41 ],
   alphaCSR[ 11 ][ 42 ],
   alphaCSR[ 11 ][ 43 ],
   alphaCSR[ 11 ][ 44 ],
   alphaCSR[ 11 ][ 45 ],
   alphaCSR[ 11 ][ 46 ],
   alphaCSR[ 11 ][ 47 ],
   alphaCSR[ 11 ][ 48 ],
   alphaCSR[ 11 ][ 49 ],
   alphaCSR[ 11 ][ 50 ],
   alphaCSR[ 11 ][ 51 ],
   alphaCSR[ 11 ][ 52 ],
   alphaCSR[ 11 ][ 53 ],
   alphaCSR[ 11 ][ 54 ],
   alphaCSR[ 11 ][ 55 ],
   alphaCSR[ 11 ][ 56 ],
   alphaCSR[ 11 ][ 57 ],
   alphaCSR[ 11 ][ 58 ],
   alphaCSR[ 11 ][ 59 ],
   alphaCSR[ 11 ][ 60 ],
   alphaCSR[ 11 ][ 61 ],
   alphaCSR[ 11 ][ 62 ],
   alphaCSR[ 11 ][ 63 ],
   alphaCSR[ 11 ][ 64 ],
   alphaCSR[ 11 ][ 65 ],
   alphaCSR[ 11 ][ 66 ],
   alphaCSR[ 11 ][ 67 ],
   alphaCSR[ 11 ][ 68 ],
   alphaCSR[ 11 ][ 69 ],
   alphaCSR[ 11 ][ 70 ],
   alphaCSR[ 11 ][ 71 ],
   alphaCSR[ 11 ][ 72 ],
   alphaCSR[ 11 ][ 73 ],
   alphaCSR[ 11 ][ 74 ],
   alphaCSR[ 11 ][ 75 ],
   alphaCSR[ 11 ][ 76 ],
   alphaCSR[ 11 ][ 77 ],
   alphaCSR[ 11 ][ 78 ],
   alphaCSR[ 11 ][ 79 ],
   alphaCSR[ 11 ][ 80 ],
   alphaCSR[ 11 ][ 81 ],
   alphaCSR[ 11 ][ 82 ],
   alphaCSR[ 11 ][ 83 ],
   alphaCSR[ 11 ][ 84 ],
   alphaCSR[ 11 ][ 85 ],
   alphaCSR[ 11 ][ 86 ],
   alphaCSR[ 11 ][ 87 ],
   alphaCSR[ 11 ][ 88 ],
   alphaCSR[ 11 ][ 89 ],
   alphaCSR[ 11 ][ 90 ],
   alphaCSR[ 11 ][ 91 ],
   alphaCSR[ 11 ][ 92 ],
   alphaCSR[ 11 ][ 93 ],
   alphaCSR[ 11 ][ 94 ],
   alphaCSR[ 11 ][ 95 ],
   alphaCSR[ 11 ][ 96 ],
   alphaCSR[ 11 ][ 97 ],
   alphaCSR[ 11 ][ 98 ],
   alphaCSR[ 11 ][ 99 ],
   alphaCSR[ 11 ][ 100 ],
   alphaCSR[ 11 ][ 101 ],
   alphaCSR[ 11 ][ 102 ],
   alphaCSR[ 11 ][ 103 ],
   alphaCSR[ 11 ][ 104 ],
   alphaCSR[ 11 ][ 105 ],
   alphaCSR[ 11 ][ 106 ],
   alphaCSR[ 11 ][ 107 ],
   alphaCSR[ 11 ][ 108 ],
   alphaCSR[ 11 ][ 109 ],
   alphaCSR[ 11 ][ 110 ],
   alphaCSR[ 11 ][ 111 ],
   alphaCSR[ 11 ][ 112 ],
   alphaCSR[ 11 ][ 113 ],
   alphaCSR[ 11 ][ 114 ],
   alphaCSR[ 11 ][ 115 ],
   alphaCSR[ 11 ][ 116 ],
   alphaCSR[ 11 ][ 117 ],
   alphaCSR[ 11 ][ 118 ],
   alphaCSR[ 11 ][ 119 ],
   alphaCSR[ 11 ][ 120 ],
   alphaCSR[ 11 ][ 121 ],
   alphaCSR[ 11 ][ 122 ],
   alphaCSR[ 11 ][ 123 ],
   alphaCSR[ 11 ][ 124 ],
   alphaCSR[ 11 ][ 125 ],
   alphaCSR[ 11 ][ 126 ],
   alphaCSR[ 11 ][ 127 ],
   alphaCSR[ 11 ][ 128 ],
   alphaCSR[ 11 ][ 129 ],
   alphaCSR[ 11 ][ 130 ],
   alphaCSR[ 11 ][ 131 ],
   alphaCSR[ 11 ][ 132 ],
   alphaCSR[ 11 ][ 133 ],
   alphaCSR[ 11 ][ 134 ],
   alphaCSR[ 11 ][ 135 ],
   alphaCSR[ 11 ][ 136 ],
   alphaCSR[ 11 ][ 137 ],
   alphaCSR[ 11 ][ 138 ],
   alphaCSR[ 11 ][ 139 ],
   alphaCSR[ 11 ][ 140 ],
   alphaCSR[ 11 ][ 141 ],
   alphaCSR[ 11 ][ 142 ],
   alphaCSR[ 11 ][ 143 ],
   alphaCSR[ 11 ][ 144 ],
   alphaCSR[ 11 ][ 145 ],
   alphaCSR[ 11 ][ 146 ],
   alphaCSR[ 11 ][ 147 ],
   alphaCSR[ 11 ][ 148 ],
   alphaCSR[ 11 ][ 149 ],
   alphaCSR[ 11 ][ 150 ],
   alphaCSR[ 11 ][ 151 ],
   alphaCSR[ 11 ][ 152 ],
   alphaCSR[ 11 ][ 153 ],
   alphaCSR[ 11 ][ 154 ],
   alphaCSR[ 11 ][ 155 ],
   alphaCSR[ 11 ][ 156 ],
   alphaCSR[ 11 ][ 157 ],
   alphaCSR[ 11 ][ 158 ],
   alphaCSR[ 11 ][ 159 ],
   alphaCSR[ 11 ][ 160 ],
   alphaCSR[ 11 ][ 161 ],
   alphaCSR[ 11 ][ 162 ],
   alphaCSR[ 11 ][ 163 ],
   alphaCSR[ 11 ][ 164 ],
   alphaCSR[ 11 ][ 165 ],
   alphaCSR[ 11 ][ 166 ],
   alphaCSR[ 11 ][ 167 ],
   alphaCSR[ 11 ][ 168 ],
   alphaCSR[ 11 ][ 169 ],
   alphaCSR[ 11 ][ 170 ],
   alphaCSR[ 11 ][ 171 ],
   alphaCSR[ 11 ][ 172 ],
   alphaCSR[ 11 ][ 173 ],
   alphaCSR[ 11 ][ 174 ],
   alphaCSR[ 11 ][ 175 ],
   alphaCSR[ 11 ][ 176 ],
   alphaCSR[ 11 ][ 177 ],
   alphaCSR[ 11 ][ 178 ],
   alphaCSR[ 11 ][ 179 ],
   alphaCSR[ 11 ][ 180 ],
   alphaCSR[ 11 ][ 181 ],
   alphaCSR[ 11 ][ 182 ],
   alphaCSR[ 11 ][ 183 ],
   alphaCSR[ 11 ][ 184 ],
   alphaCSR[ 11 ][ 185 ],
   alphaCSR[ 11 ][ 186 ],
   alphaCSR[ 11 ][ 187 ],
   alphaCSR[ 11 ][ 188 ],
   alphaCSR[ 11 ][ 189 ],
   alphaCSR[ 11 ][ 190 ],
   alphaCSR[ 11 ][ 191 ],
   alphaCSR[ 11 ][ 192 ],
   alphaCSR[ 11 ][ 193 ],
   alphaCSR[ 11 ][ 194 ],
   alphaCSR[ 11 ][ 195 ],
   alphaCSR[ 11 ][ 196 ],
   alphaCSR[ 11 ][ 197 ],
   alphaCSR[ 11 ][ 198 ],
   alphaCSR[ 11 ][ 199 ],
   alphaCSR[ 11 ][ 200 ],
   alphaCSR[ 11 ][ 201 ],
   alphaCSR[ 11 ][ 202 ],
   alphaCSR[ 11 ][ 203 ],
   alphaCSR[ 11 ][ 204 ],
   alphaCSR[ 11 ][ 205 ],
   alphaCSR[ 11 ][ 206 ],
   alphaCSR[ 11 ][ 207 ],
   alphaCSR[ 11 ][ 208 ],
   alphaCSR[ 11 ][ 209 ],
   alphaCSR[ 11 ][ 210 ],
   alphaCSR[ 11 ][ 211 ],
   alphaCSR[ 11 ][ 212 ],
   alphaCSR[ 11 ][ 213 ],
   alphaCSR[ 11 ][ 214 ],
   alphaCSR[ 11 ][ 215 ],
   alphaCSR[ 11 ][ 216 ],
   alphaCSR[ 11 ][ 217 ],
   alphaCSR[ 11 ][ 218 ],
   alphaCSR[ 11 ][ 219 ],
   alphaCSR[ 11 ][ 220 ],
   alphaCSR[ 11 ][ 221 ],
   alphaCSR[ 11 ][ 222 ],
   alphaCSR[ 11 ][ 223 ],
   alphaCSR[ 11 ][ 224 ],
   alphaCSR[ 11 ][ 225 ],
   alphaCSR[ 11 ][ 226 ],
   alphaCSR[ 11 ][ 227 ],
   alphaCSR[ 11 ][ 228 ],
   alphaCSR[ 11 ][ 229 ],
   alphaCSR[ 11 ][ 230 ],
   alphaCSR[ 11 ][ 231 ],
   alphaCSR[ 11 ][ 232 ],
   alphaCSR[ 11 ][ 233 ],
   alphaCSR[ 11 ][ 234 ],
   alphaCSR[ 11 ][ 235 ],
   alphaCSR[ 11 ][ 236 ],
   alphaCSR[ 11 ][ 237 ],
   alphaCSR[ 11 ][ 238 ],
   alphaCSR[ 11 ][ 239 ],
   alphaCSR[ 11 ][ 240 ],
   alphaCSR[ 11 ][ 241 ],
   alphaCSR[ 11 ][ 242 ],
   alphaCSR[ 11 ][ 243 ],
   alphaCSR[ 11 ][ 244 ],
   alphaCSR[ 11 ][ 245 ],
   alphaCSR[ 11 ][ 246 ],
   alphaCSR[ 11 ][ 247 ],
   alphaCSR[ 11 ][ 248 ],
   alphaCSR[ 11 ][ 249 ],
   alphaCSR[ 11 ][ 250 ],
   alphaCSR[ 11 ][ 251 ],
   alphaCSR[ 11 ][ 252 ],
   alphaCSR[ 11 ][ 253 ],
   alphaCSR[ 11 ][ 254 ],
   alphaCSR[ 11 ][ 255 ],
   alphaCSR[ 11 ][ 256 ],
   alphaCSR[ 11 ][ 257 ],
   alphaCSR[ 11 ][ 258 ],
   alphaCSR[ 11 ][ 259 ],
   alphaCSR[ 11 ][ 260 ],
   alphaCSR[ 11 ][ 261 ],
   alphaCSR[ 11 ][ 262 ],
   alphaCSR[ 11 ][ 263 ],
   alphaCSR[ 11 ][ 264 ],
   alphaCSR[ 11 ][ 265 ],
   alphaCSR[ 11 ][ 266 ],
   alphaCSR[ 11 ][ 267 ],
   alphaCSR[ 11 ][ 268 ],
   alphaCSR[ 11 ][ 269 ],
   alphaCSR[ 11 ][ 270 ],
   alphaCSR[ 11 ][ 271 ],
   alphaCSR[ 11 ][ 272 ],
   alphaCSR[ 11 ][ 273 ],
   alphaCSR[ 11 ][ 274 ],
   alphaCSR[ 11 ][ 275 ],
   alphaCSR[ 11 ][ 276 ],
   alphaCSR[ 11 ][ 277 ],
   alphaCSR[ 11 ][ 278 ],
   alphaCSR[ 11 ][ 279 ],
   alphaCSR[ 11 ][ 280 ],
   alphaCSR[ 11 ][ 281 ],
   alphaCSR[ 11 ][ 282 ],
   alphaCSR[ 11 ][ 283 ],
   alphaCSR[ 11 ][ 284 ],
   alphaCSR[ 11 ][ 285 ],
   alphaCSR[ 11 ][ 286 ],
   alphaCSR[ 11 ][ 287 ],
   alphaCSR[ 11 ][ 288 ],
   alphaCSR[ 11 ][ 289 ],
   alphaCSR[ 11 ][ 290 ],
   alphaCSR[ 11 ][ 291 ],
   alphaCSR[ 11 ][ 292 ],
   alphaCSR[ 11 ][ 293 ],
   alphaCSR[ 11 ][ 294 ],
   alphaCSR[ 11 ][ 295 ],
   alphaCSR[ 11 ][ 296 ],
   alphaCSR[ 11 ][ 297 ],
   alphaCSR[ 11 ][ 298 ],
   alphaCSR[ 11 ][ 299 ],
   alphaCSR[ 11 ][ 300 ],
   alphaCSR[ 11 ][ 301 ],
   alphaCSR[ 11 ][ 302 ],
   alphaCSR[ 11 ][ 303 ],
   alphaCSR[ 11 ][ 304 ],
   alphaCSR[ 11 ][ 305 ],
   alphaCSR[ 11 ][ 306 ],
   alphaCSR[ 11 ][ 307 ],
   alphaCSR[ 11 ][ 308 ],
   alphaCSR[ 11 ][ 309 ],
   alphaCSR[ 11 ][ 310 ],
   alphaCSR[ 11 ][ 311 ],
   alphaCSR[ 11 ][ 312 ],
   alphaCSR[ 11 ][ 313 ],
   alphaCSR[ 11 ][ 314 ],
   alphaCSR[ 11 ][ 315 ],
   alphaCSR[ 11 ][ 316 ],
   alphaCSR[ 11 ][ 317 ],
   alphaCSR[ 11 ][ 318 ],
   alphaCSR[ 11 ][ 319 ],
   alphaCSR[ 11 ][ 320 ],
   alphaCSR[ 11 ][ 321 ],
   alphaCSR[ 11 ][ 322 ],
   alphaCSR[ 11 ][ 323 ],
   alphaCSR[ 11 ][ 324 ],
   alphaCSR[ 11 ][ 325 ],
   alphaCSR[ 11 ][ 326 ],
   alphaCSR[ 11 ][ 327 ],
   alphaCSR[ 11 ][ 328 ],
   alphaCSR[ 11 ][ 329 ],
   alphaCSR[ 11 ][ 330 ],
   alphaCSR[ 11 ][ 331 ],
   alphaCSR[ 11 ][ 332 ],
   alphaCSR[ 11 ][ 333 ],
   alphaCSR[ 11 ][ 334 ],
   alphaCSR[ 11 ][ 335 ],
   alphaCSR[ 11 ][ 336 ],
   alphaCSR[ 11 ][ 337 ],
   alphaCSR[ 11 ][ 338 ],
   alphaCSR[ 11 ][ 339 ],
   alphaCSR[ 11 ][ 340 ],
   alphaCSR[ 11 ][ 341 ],
   alphaCSR[ 11 ][ 342 ],
   alphaCSR[ 11 ][ 343 ],
   alphaCSR[ 11 ][ 344 ],
   alphaCSR[ 11 ][ 345 ],
   alphaCSR[ 11 ][ 346 ],
   alphaCSR[ 11 ][ 347 ],
   alphaCSR[ 11 ][ 348 ],
   alphaCSR[ 11 ][ 349 ],
   alphaCSR[ 11 ][ 350 ],
   alphaCSR[ 11 ][ 351 ],
   alphaCSR[ 11 ][ 352 ],
   alphaCSR[ 11 ][ 353 ],
   alphaCSR[ 11 ][ 354 ],
   alphaCSR[ 11 ][ 355 ],
   alphaCSR[ 11 ][ 356 ],
   alphaCSR[ 11 ][ 357 ],
   alphaCSR[ 11 ][ 358 ],
   alphaCSR[ 11 ][ 359 ],
   alphaCSR[ 11 ][ 360 ],
   alphaCSR[ 11 ][ 361 ],
   alphaCSR[ 11 ][ 362 ],
   alphaCSR[ 11 ][ 363 ],
   alphaCSR[ 11 ][ 364 ],
   alphaCSR[ 11 ][ 365 ],
   alphaCSR[ 11 ][ 366 ],
   alphaCSR[ 11 ][ 367 ],
   alphaCSR[ 11 ][ 368 ],
   alphaCSR[ 11 ][ 369 ],
   alphaCSR[ 11 ][ 370 ],
   alphaCSR[ 11 ][ 371 ],
   alphaCSR[ 11 ][ 372 ],
   alphaCSR[ 11 ][ 373 ],
   alphaCSR[ 11 ][ 374 ],
   alphaCSR[ 11 ][ 375 ],
   alphaCSR[ 11 ][ 376 ],
   alphaCSR[ 11 ][ 377 ],
   alphaCSR[ 11 ][ 378 ],
   alphaCSR[ 11 ][ 379 ],
   alphaCSR[ 11 ][ 380 ],
   alphaCSR[ 11 ][ 381 ],
   alphaCSR[ 11 ][ 382 ],
   alphaCSR[ 11 ][ 383 ],
   alphaCSR[ 12 ][ 0 ],
   alphaCSR[ 12 ][ 1 ],
   alphaCSR[ 12 ][ 2 ],
   alphaCSR[ 12 ][ 3 ],
   alphaCSR[ 12 ][ 4 ],
   alphaCSR[ 12 ][ 5 ],
   alphaCSR[ 12 ][ 6 ],
   alphaCSR[ 12 ][ 7 ],
   alphaCSR[ 12 ][ 8 ],
   alphaCSR[ 12 ][ 9 ],
   alphaCSR[ 12 ][ 10 ],
   alphaCSR[ 12 ][ 11 ],
   alphaCSR[ 12 ][ 12 ],
   alphaCSR[ 12 ][ 13 ],
   alphaCSR[ 12 ][ 14 ],
   alphaCSR[ 12 ][ 15 ],
   alphaCSR[ 12 ][ 16 ],
   alphaCSR[ 12 ][ 17 ],
   alphaCSR[ 12 ][ 18 ],
   alphaCSR[ 12 ][ 19 ],
   alphaCSR[ 12 ][ 20 ],
   alphaCSR[ 12 ][ 21 ],
   alphaCSR[ 12 ][ 22 ],
   alphaCSR[ 12 ][ 23 ],
   alphaCSR[ 12 ][ 24 ],
   alphaCSR[ 12 ][ 25 ],
   alphaCSR[ 12 ][ 26 ],
   alphaCSR[ 12 ][ 27 ],
   alphaCSR[ 12 ][ 28 ],
   alphaCSR[ 12 ][ 29 ],
   alphaCSR[ 12 ][ 30 ],
   alphaCSR[ 12 ][ 31 ],
   alphaCSR[ 12 ][ 32 ],
   alphaCSR[ 12 ][ 33 ],
   alphaCSR[ 12 ][ 34 ],
   alphaCSR[ 12 ][ 35 ],
   alphaCSR[ 12 ][ 36 ],
   alphaCSR[ 12 ][ 37 ],
   alphaCSR[ 12 ][ 38 ],
   alphaCSR[ 12 ][ 39 ],
   alphaCSR[ 12 ][ 40 ],
   alphaCSR[ 12 ][ 41 ],
   alphaCSR[ 12 ][ 42 ],
   alphaCSR[ 12 ][ 43 ],
   alphaCSR[ 12 ][ 44 ],
   alphaCSR[ 12 ][ 45 ],
   alphaCSR[ 12 ][ 46 ],
   alphaCSR[ 12 ][ 47 ],
   alphaCSR[ 12 ][ 48 ],
   alphaCSR[ 12 ][ 49 ],
   alphaCSR[ 12 ][ 50 ],
   alphaCSR[ 12 ][ 51 ],
   alphaCSR[ 12 ][ 52 ],
   alphaCSR[ 12 ][ 53 ],
   alphaCSR[ 12 ][ 54 ],
   alphaCSR[ 12 ][ 55 ],
   alphaCSR[ 12 ][ 56 ],
   alphaCSR[ 12 ][ 57 ],
   alphaCSR[ 12 ][ 58 ],
   alphaCSR[ 12 ][ 59 ],
   alphaCSR[ 12 ][ 60 ],
   alphaCSR[ 12 ][ 61 ],
   alphaCSR[ 12 ][ 62 ],
   alphaCSR[ 12 ][ 63 ],
   alphaCSR[ 12 ][ 64 ],
   alphaCSR[ 12 ][ 65 ],
   alphaCSR[ 12 ][ 66 ],
   alphaCSR[ 12 ][ 67 ],
   alphaCSR[ 12 ][ 68 ],
   alphaCSR[ 12 ][ 69 ],
   alphaCSR[ 12 ][ 70 ],
   alphaCSR[ 12 ][ 71 ],
   alphaCSR[ 12 ][ 72 ],
   alphaCSR[ 12 ][ 73 ],
   alphaCSR[ 12 ][ 74 ],
   alphaCSR[ 12 ][ 75 ],
   alphaCSR[ 12 ][ 76 ],
   alphaCSR[ 12 ][ 77 ],
   alphaCSR[ 12 ][ 78 ],
   alphaCSR[ 12 ][ 79 ],
   alphaCSR[ 12 ][ 80 ],
   alphaCSR[ 12 ][ 81 ],
   alphaCSR[ 12 ][ 82 ],
   alphaCSR[ 12 ][ 83 ],
   alphaCSR[ 12 ][ 84 ],
   alphaCSR[ 12 ][ 85 ],
   alphaCSR[ 12 ][ 86 ],
   alphaCSR[ 12 ][ 87 ],
   alphaCSR[ 12 ][ 88 ],
   alphaCSR[ 12 ][ 89 ],
   alphaCSR[ 12 ][ 90 ],
   alphaCSR[ 12 ][ 91 ],
   alphaCSR[ 12 ][ 92 ],
   alphaCSR[ 12 ][ 93 ],
   alphaCSR[ 12 ][ 94 ],
   alphaCSR[ 12 ][ 95 ],
   alphaCSR[ 12 ][ 96 ],
   alphaCSR[ 12 ][ 97 ],
   alphaCSR[ 12 ][ 98 ],
   alphaCSR[ 12 ][ 99 ],
   alphaCSR[ 12 ][ 100 ],
   alphaCSR[ 12 ][ 101 ],
   alphaCSR[ 12 ][ 102 ],
   alphaCSR[ 12 ][ 103 ],
   alphaCSR[ 12 ][ 104 ],
   alphaCSR[ 12 ][ 105 ],
   alphaCSR[ 12 ][ 106 ],
   alphaCSR[ 12 ][ 107 ],
   alphaCSR[ 12 ][ 108 ],
   alphaCSR[ 12 ][ 109 ],
   alphaCSR[ 12 ][ 110 ],
   alphaCSR[ 12 ][ 111 ],
   alphaCSR[ 12 ][ 112 ],
   alphaCSR[ 12 ][ 113 ],
   alphaCSR[ 12 ][ 114 ],
   alphaCSR[ 12 ][ 115 ],
   alphaCSR[ 12 ][ 116 ],
   alphaCSR[ 12 ][ 117 ],
   alphaCSR[ 12 ][ 118 ],
   alphaCSR[ 12 ][ 119 ],
   alphaCSR[ 12 ][ 120 ],
   alphaCSR[ 12 ][ 121 ],
   alphaCSR[ 12 ][ 122 ],
   alphaCSR[ 12 ][ 123 ],
   alphaCSR[ 12 ][ 124 ],
   alphaCSR[ 12 ][ 125 ],
   alphaCSR[ 12 ][ 126 ],
   alphaCSR[ 12 ][ 127 ],
   alphaCSR[ 12 ][ 128 ],
   alphaCSR[ 12 ][ 129 ],
   alphaCSR[ 12 ][ 130 ],
   alphaCSR[ 12 ][ 131 ],
   alphaCSR[ 12 ][ 132 ],
   alphaCSR[ 12 ][ 133 ],
   alphaCSR[ 12 ][ 134 ],
   alphaCSR[ 12 ][ 135 ],
   alphaCSR[ 12 ][ 136 ],
   alphaCSR[ 12 ][ 137 ],
   alphaCSR[ 12 ][ 138 ],
   alphaCSR[ 12 ][ 139 ],
   alphaCSR[ 12 ][ 140 ],
   alphaCSR[ 12 ][ 141 ],
   alphaCSR[ 12 ][ 142 ],
   alphaCSR[ 12 ][ 143 ],
   alphaCSR[ 12 ][ 144 ],
   alphaCSR[ 12 ][ 145 ],
   alphaCSR[ 12 ][ 146 ],
   alphaCSR[ 12 ][ 147 ],
   alphaCSR[ 12 ][ 148 ],
   alphaCSR[ 12 ][ 149 ],
   alphaCSR[ 12 ][ 150 ],
   alphaCSR[ 12 ][ 151 ],
   alphaCSR[ 12 ][ 152 ],
   alphaCSR[ 12 ][ 153 ],
   alphaCSR[ 12 ][ 154 ],
   alphaCSR[ 12 ][ 155 ],
   alphaCSR[ 12 ][ 156 ],
   alphaCSR[ 12 ][ 157 ],
   alphaCSR[ 12 ][ 158 ],
   alphaCSR[ 12 ][ 159 ],
   alphaCSR[ 12 ][ 160 ],
   alphaCSR[ 12 ][ 161 ],
   alphaCSR[ 12 ][ 162 ],
   alphaCSR[ 12 ][ 163 ],
   alphaCSR[ 12 ][ 164 ],
   alphaCSR[ 12 ][ 165 ],
   alphaCSR[ 12 ][ 166 ],
   alphaCSR[ 12 ][ 167 ],
   alphaCSR[ 12 ][ 168 ],
   alphaCSR[ 12 ][ 169 ],
   alphaCSR[ 12 ][ 170 ],
   alphaCSR[ 12 ][ 171 ],
   alphaCSR[ 12 ][ 172 ],
   alphaCSR[ 12 ][ 173 ],
   alphaCSR[ 12 ][ 174 ],
   alphaCSR[ 12 ][ 175 ],
   alphaCSR[ 12 ][ 176 ],
   alphaCSR[ 12 ][ 177 ],
   alphaCSR[ 12 ][ 178 ],
   alphaCSR[ 12 ][ 179 ],
   alphaCSR[ 12 ][ 180 ],
   alphaCSR[ 12 ][ 181 ],
   alphaCSR[ 12 ][ 182 ],
   alphaCSR[ 12 ][ 183 ],
   alphaCSR[ 12 ][ 184 ],
   alphaCSR[ 12 ][ 185 ],
   alphaCSR[ 12 ][ 186 ],
   alphaCSR[ 12 ][ 187 ],
   alphaCSR[ 12 ][ 188 ],
   alphaCSR[ 12 ][ 189 ],
   alphaCSR[ 12 ][ 190 ],
   alphaCSR[ 12 ][ 191 ],
   alphaCSR[ 12 ][ 192 ],
   alphaCSR[ 12 ][ 193 ],
   alphaCSR[ 12 ][ 194 ],
   alphaCSR[ 12 ][ 195 ],
   alphaCSR[ 12 ][ 196 ],
   alphaCSR[ 12 ][ 197 ],
   alphaCSR[ 12 ][ 198 ],
   alphaCSR[ 12 ][ 199 ],
   alphaCSR[ 12 ][ 200 ],
   alphaCSR[ 12 ][ 201 ],
   alphaCSR[ 12 ][ 202 ],
   alphaCSR[ 12 ][ 203 ],
   alphaCSR[ 12 ][ 204 ],
   alphaCSR[ 12 ][ 205 ],
   alphaCSR[ 12 ][ 206 ],
   alphaCSR[ 12 ][ 207 ],
   alphaCSR[ 12 ][ 208 ],
   alphaCSR[ 12 ][ 209 ],
   alphaCSR[ 12 ][ 210 ],
   alphaCSR[ 12 ][ 211 ],
   alphaCSR[ 12 ][ 212 ],
   alphaCSR[ 12 ][ 213 ],
   alphaCSR[ 12 ][ 214 ],
   alphaCSR[ 12 ][ 215 ],
   alphaCSR[ 12 ][ 216 ],
   alphaCSR[ 12 ][ 217 ],
   alphaCSR[ 12 ][ 218 ],
   alphaCSR[ 12 ][ 219 ],
   alphaCSR[ 12 ][ 220 ],
   alphaCSR[ 12 ][ 221 ],
   alphaCSR[ 12 ][ 222 ],
   alphaCSR[ 12 ][ 223 ],
   alphaCSR[ 12 ][ 224 ],
   alphaCSR[ 12 ][ 225 ],
   alphaCSR[ 12 ][ 226 ],
   alphaCSR[ 12 ][ 227 ],
   alphaCSR[ 12 ][ 228 ],
   alphaCSR[ 12 ][ 229 ],
   alphaCSR[ 12 ][ 230 ],
   alphaCSR[ 12 ][ 231 ],
   alphaCSR[ 12 ][ 232 ],
   alphaCSR[ 12 ][ 233 ],
   alphaCSR[ 12 ][ 234 ],
   alphaCSR[ 12 ][ 235 ],
   alphaCSR[ 12 ][ 236 ],
   alphaCSR[ 12 ][ 237 ],
   alphaCSR[ 12 ][ 238 ],
   alphaCSR[ 12 ][ 239 ],
   alphaCSR[ 12 ][ 240 ],
   alphaCSR[ 12 ][ 241 ],
   alphaCSR[ 12 ][ 242 ],
   alphaCSR[ 12 ][ 243 ],
   alphaCSR[ 12 ][ 244 ],
   alphaCSR[ 12 ][ 245 ],
   alphaCSR[ 12 ][ 246 ],
   alphaCSR[ 12 ][ 247 ],
   alphaCSR[ 12 ][ 248 ],
   alphaCSR[ 12 ][ 249 ],
   alphaCSR[ 12 ][ 250 ],
   alphaCSR[ 12 ][ 251 ],
   alphaCSR[ 12 ][ 252 ],
   alphaCSR[ 12 ][ 253 ],
   alphaCSR[ 12 ][ 254 ],
   alphaCSR[ 12 ][ 255 ],
   alphaCSR[ 12 ][ 256 ],
   alphaCSR[ 12 ][ 257 ],
   alphaCSR[ 12 ][ 258 ],
   alphaCSR[ 12 ][ 259 ],
   alphaCSR[ 12 ][ 260 ],
   alphaCSR[ 12 ][ 261 ],
   alphaCSR[ 12 ][ 262 ],
   alphaCSR[ 12 ][ 263 ],
   alphaCSR[ 12 ][ 264 ],
   alphaCSR[ 12 ][ 265 ],
   alphaCSR[ 12 ][ 266 ],
   alphaCSR[ 12 ][ 267 ],
   alphaCSR[ 12 ][ 268 ],
   alphaCSR[ 12 ][ 269 ],
   alphaCSR[ 12 ][ 270 ],
   alphaCSR[ 12 ][ 271 ],
   alphaCSR[ 12 ][ 272 ],
   alphaCSR[ 12 ][ 273 ],
   alphaCSR[ 12 ][ 274 ],
   alphaCSR[ 12 ][ 275 ],
   alphaCSR[ 12 ][ 276 ],
   alphaCSR[ 12 ][ 277 ],
   alphaCSR[ 12 ][ 278 ],
   alphaCSR[ 12 ][ 279 ],
   alphaCSR[ 12 ][ 280 ],
   alphaCSR[ 12 ][ 281 ],
   alphaCSR[ 12 ][ 282 ],
   alphaCSR[ 12 ][ 283 ],
   alphaCSR[ 12 ][ 284 ],
   alphaCSR[ 12 ][ 285 ],
   alphaCSR[ 12 ][ 286 ],
   alphaCSR[ 12 ][ 287 ],
   alphaCSR[ 12 ][ 288 ],
   alphaCSR[ 12 ][ 289 ],
   alphaCSR[ 12 ][ 290 ],
   alphaCSR[ 12 ][ 291 ],
   alphaCSR[ 12 ][ 292 ],
   alphaCSR[ 12 ][ 293 ],
   alphaCSR[ 12 ][ 294 ],
   alphaCSR[ 12 ][ 295 ],
   alphaCSR[ 12 ][ 296 ],
   alphaCSR[ 12 ][ 297 ],
   alphaCSR[ 12 ][ 298 ],
   alphaCSR[ 12 ][ 299 ],
   alphaCSR[ 12 ][ 300 ],
   alphaCSR[ 12 ][ 301 ],
   alphaCSR[ 12 ][ 302 ],
   alphaCSR[ 12 ][ 303 ],
   alphaCSR[ 12 ][ 304 ],
   alphaCSR[ 12 ][ 305 ],
   alphaCSR[ 12 ][ 306 ],
   alphaCSR[ 12 ][ 307 ],
   alphaCSR[ 12 ][ 308 ],
   alphaCSR[ 12 ][ 309 ],
   alphaCSR[ 12 ][ 310 ],
   alphaCSR[ 12 ][ 311 ],
   alphaCSR[ 12 ][ 312 ],
   alphaCSR[ 12 ][ 313 ],
   alphaCSR[ 12 ][ 314 ],
   alphaCSR[ 12 ][ 315 ],
   alphaCSR[ 12 ][ 316 ],
   alphaCSR[ 12 ][ 317 ],
   alphaCSR[ 12 ][ 318 ],
   alphaCSR[ 12 ][ 319 ],
   alphaCSR[ 12 ][ 320 ],
   alphaCSR[ 12 ][ 321 ],
   alphaCSR[ 12 ][ 322 ],
   alphaCSR[ 12 ][ 323 ],
   alphaCSR[ 12 ][ 324 ],
   alphaCSR[ 12 ][ 325 ],
   alphaCSR[ 12 ][ 326 ],
   alphaCSR[ 12 ][ 327 ],
   alphaCSR[ 12 ][ 328 ],
   alphaCSR[ 12 ][ 329 ],
   alphaCSR[ 12 ][ 330 ],
   alphaCSR[ 12 ][ 331 ],
   alphaCSR[ 12 ][ 332 ],
   alphaCSR[ 12 ][ 333 ],
   alphaCSR[ 12 ][ 334 ],
   alphaCSR[ 12 ][ 335 ],
   alphaCSR[ 12 ][ 336 ],
   alphaCSR[ 12 ][ 337 ],
   alphaCSR[ 12 ][ 338 ],
   alphaCSR[ 12 ][ 339 ],
   alphaCSR[ 12 ][ 340 ],
   alphaCSR[ 12 ][ 341 ],
   alphaCSR[ 12 ][ 342 ],
   alphaCSR[ 12 ][ 343 ],
   alphaCSR[ 12 ][ 344 ],
   alphaCSR[ 12 ][ 345 ],
   alphaCSR[ 12 ][ 346 ],
   alphaCSR[ 12 ][ 347 ],
   alphaCSR[ 12 ][ 348 ],
   alphaCSR[ 12 ][ 349 ],
   alphaCSR[ 12 ][ 350 ],
   alphaCSR[ 12 ][ 351 ],
   alphaCSR[ 12 ][ 352 ],
   alphaCSR[ 12 ][ 353 ],
   alphaCSR[ 12 ][ 354 ],
   alphaCSR[ 12 ][ 355 ],
   alphaCSR[ 12 ][ 356 ],
   alphaCSR[ 12 ][ 357 ],
   alphaCSR[ 12 ][ 358 ],
   alphaCSR[ 12 ][ 359 ],
   alphaCSR[ 12 ][ 360 ],
   alphaCSR[ 12 ][ 361 ],
   alphaCSR[ 12 ][ 362 ],
   alphaCSR[ 12 ][ 363 ],
   alphaCSR[ 12 ][ 364 ],
   alphaCSR[ 12 ][ 365 ],
   alphaCSR[ 12 ][ 366 ],
   alphaCSR[ 12 ][ 367 ],
   alphaCSR[ 12 ][ 368 ],
   alphaCSR[ 12 ][ 369 ],
   alphaCSR[ 12 ][ 370 ],
   alphaCSR[ 12 ][ 371 ],
   alphaCSR[ 12 ][ 372 ],
   alphaCSR[ 12 ][ 373 ],
   alphaCSR[ 12 ][ 374 ],
   alphaCSR[ 12 ][ 375 ],
   alphaCSR[ 12 ][ 376 ],
   alphaCSR[ 12 ][ 377 ],
   alphaCSR[ 12 ][ 378 ],
   alphaCSR[ 12 ][ 379 ],
   alphaCSR[ 12 ][ 380 ],
   alphaCSR[ 12 ][ 381 ],
   alphaCSR[ 12 ][ 382 ],
   alphaCSR[ 12 ][ 383 ],
   alphaCSR[ 13 ][ 0 ],
   alphaCSR[ 13 ][ 1 ],
   alphaCSR[ 13 ][ 2 ],
   alphaCSR[ 13 ][ 3 ],
   alphaCSR[ 13 ][ 4 ],
   alphaCSR[ 13 ][ 5 ],
   alphaCSR[ 13 ][ 6 ],
   alphaCSR[ 13 ][ 7 ],
   alphaCSR[ 13 ][ 8 ],
   alphaCSR[ 13 ][ 9 ],
   alphaCSR[ 13 ][ 10 ],
   alphaCSR[ 13 ][ 11 ],
   alphaCSR[ 13 ][ 12 ],
   alphaCSR[ 13 ][ 13 ],
   alphaCSR[ 13 ][ 14 ],
   alphaCSR[ 13 ][ 15 ],
   alphaCSR[ 13 ][ 16 ],
   alphaCSR[ 13 ][ 17 ],
   alphaCSR[ 13 ][ 18 ],
   alphaCSR[ 13 ][ 19 ],
   alphaCSR[ 13 ][ 20 ],
   alphaCSR[ 13 ][ 21 ],
   alphaCSR[ 13 ][ 22 ],
   alphaCSR[ 13 ][ 23 ],
   alphaCSR[ 13 ][ 24 ],
   alphaCSR[ 13 ][ 25 ],
   alphaCSR[ 13 ][ 26 ],
   alphaCSR[ 13 ][ 27 ],
   alphaCSR[ 13 ][ 28 ],
   alphaCSR[ 13 ][ 29 ],
   alphaCSR[ 13 ][ 30 ],
   alphaCSR[ 13 ][ 31 ],
   alphaCSR[ 13 ][ 32 ],
   alphaCSR[ 13 ][ 33 ],
   alphaCSR[ 13 ][ 34 ],
   alphaCSR[ 13 ][ 35 ],
   alphaCSR[ 13 ][ 36 ],
   alphaCSR[ 13 ][ 37 ],
   alphaCSR[ 13 ][ 38 ],
   alphaCSR[ 13 ][ 39 ],
   alphaCSR[ 13 ][ 40 ],
   alphaCSR[ 13 ][ 41 ],
   alphaCSR[ 13 ][ 42 ],
   alphaCSR[ 13 ][ 43 ],
   alphaCSR[ 13 ][ 44 ],
   alphaCSR[ 13 ][ 45 ],
   alphaCSR[ 13 ][ 46 ],
   alphaCSR[ 13 ][ 47 ],
   alphaCSR[ 13 ][ 48 ],
   alphaCSR[ 13 ][ 49 ],
   alphaCSR[ 13 ][ 50 ],
   alphaCSR[ 13 ][ 51 ],
   alphaCSR[ 13 ][ 52 ],
   alphaCSR[ 13 ][ 53 ],
   alphaCSR[ 13 ][ 54 ],
   alphaCSR[ 13 ][ 55 ],
   alphaCSR[ 13 ][ 56 ],
   alphaCSR[ 13 ][ 57 ],
   alphaCSR[ 13 ][ 58 ],
   alphaCSR[ 13 ][ 59 ],
   alphaCSR[ 13 ][ 60 ],
   alphaCSR[ 13 ][ 61 ],
   alphaCSR[ 13 ][ 62 ],
   alphaCSR[ 13 ][ 63 ],
   alphaCSR[ 13 ][ 64 ],
   alphaCSR[ 13 ][ 65 ],
   alphaCSR[ 13 ][ 66 ],
   alphaCSR[ 13 ][ 67 ],
   alphaCSR[ 13 ][ 68 ],
   alphaCSR[ 13 ][ 69 ],
   alphaCSR[ 13 ][ 70 ],
   alphaCSR[ 13 ][ 71 ],
   alphaCSR[ 13 ][ 72 ],
   alphaCSR[ 13 ][ 73 ],
   alphaCSR[ 13 ][ 74 ],
   alphaCSR[ 13 ][ 75 ],
   alphaCSR[ 13 ][ 76 ],
   alphaCSR[ 13 ][ 77 ],
   alphaCSR[ 13 ][ 78 ],
   alphaCSR[ 13 ][ 79 ],
   alphaCSR[ 13 ][ 80 ],
   alphaCSR[ 13 ][ 81 ],
   alphaCSR[ 13 ][ 82 ],
   alphaCSR[ 13 ][ 83 ],
   alphaCSR[ 13 ][ 84 ],
   alphaCSR[ 13 ][ 85 ],
   alphaCSR[ 13 ][ 86 ],
   alphaCSR[ 13 ][ 87 ],
   alphaCSR[ 13 ][ 88 ],
   alphaCSR[ 13 ][ 89 ],
   alphaCSR[ 13 ][ 90 ],
   alphaCSR[ 13 ][ 91 ],
   alphaCSR[ 13 ][ 92 ],
   alphaCSR[ 13 ][ 93 ],
   alphaCSR[ 13 ][ 94 ],
   alphaCSR[ 13 ][ 95 ],
   alphaCSR[ 13 ][ 96 ],
   alphaCSR[ 13 ][ 97 ],
   alphaCSR[ 13 ][ 98 ],
   alphaCSR[ 13 ][ 99 ],
   alphaCSR[ 13 ][ 100 ],
   alphaCSR[ 13 ][ 101 ],
   alphaCSR[ 13 ][ 102 ],
   alphaCSR[ 13 ][ 103 ],
   alphaCSR[ 13 ][ 104 ],
   alphaCSR[ 13 ][ 105 ],
   alphaCSR[ 13 ][ 106 ],
   alphaCSR[ 13 ][ 107 ],
   alphaCSR[ 13 ][ 108 ],
   alphaCSR[ 13 ][ 109 ],
   alphaCSR[ 13 ][ 110 ],
   alphaCSR[ 13 ][ 111 ],
   alphaCSR[ 13 ][ 112 ],
   alphaCSR[ 13 ][ 113 ],
   alphaCSR[ 13 ][ 114 ],
   alphaCSR[ 13 ][ 115 ],
   alphaCSR[ 13 ][ 116 ],
   alphaCSR[ 13 ][ 117 ],
   alphaCSR[ 13 ][ 118 ],
   alphaCSR[ 13 ][ 119 ],
   alphaCSR[ 13 ][ 120 ],
   alphaCSR[ 13 ][ 121 ],
   alphaCSR[ 13 ][ 122 ],
   alphaCSR[ 13 ][ 123 ],
   alphaCSR[ 13 ][ 124 ],
   alphaCSR[ 13 ][ 125 ],
   alphaCSR[ 13 ][ 126 ],
   alphaCSR[ 13 ][ 127 ],
   alphaCSR[ 13 ][ 128 ],
   alphaCSR[ 13 ][ 129 ],
   alphaCSR[ 13 ][ 130 ],
   alphaCSR[ 13 ][ 131 ],
   alphaCSR[ 13 ][ 132 ],
   alphaCSR[ 13 ][ 133 ],
   alphaCSR[ 13 ][ 134 ],
   alphaCSR[ 13 ][ 135 ],
   alphaCSR[ 13 ][ 136 ],
   alphaCSR[ 13 ][ 137 ],
   alphaCSR[ 13 ][ 138 ],
   alphaCSR[ 13 ][ 139 ],
   alphaCSR[ 13 ][ 140 ],
   alphaCSR[ 13 ][ 141 ],
   alphaCSR[ 13 ][ 142 ],
   alphaCSR[ 13 ][ 143 ],
   alphaCSR[ 13 ][ 144 ],
   alphaCSR[ 13 ][ 145 ],
   alphaCSR[ 13 ][ 146 ],
   alphaCSR[ 13 ][ 147 ],
   alphaCSR[ 13 ][ 148 ],
   alphaCSR[ 13 ][ 149 ],
   alphaCSR[ 13 ][ 150 ],
   alphaCSR[ 13 ][ 151 ],
   alphaCSR[ 13 ][ 152 ],
   alphaCSR[ 13 ][ 153 ],
   alphaCSR[ 13 ][ 154 ],
   alphaCSR[ 13 ][ 155 ],
   alphaCSR[ 13 ][ 156 ],
   alphaCSR[ 13 ][ 157 ],
   alphaCSR[ 13 ][ 158 ],
   alphaCSR[ 13 ][ 159 ],
   alphaCSR[ 13 ][ 160 ],
   alphaCSR[ 13 ][ 161 ],
   alphaCSR[ 13 ][ 162 ],
   alphaCSR[ 13 ][ 163 ],
   alphaCSR[ 13 ][ 164 ],
   alphaCSR[ 13 ][ 165 ],
   alphaCSR[ 13 ][ 166 ],
   alphaCSR[ 13 ][ 167 ],
   alphaCSR[ 13 ][ 168 ],
   alphaCSR[ 13 ][ 169 ],
   alphaCSR[ 13 ][ 170 ],
   alphaCSR[ 13 ][ 171 ],
   alphaCSR[ 13 ][ 172 ],
   alphaCSR[ 13 ][ 173 ],
   alphaCSR[ 13 ][ 174 ],
   alphaCSR[ 13 ][ 175 ],
   alphaCSR[ 13 ][ 176 ],
   alphaCSR[ 13 ][ 177 ],
   alphaCSR[ 13 ][ 178 ],
   alphaCSR[ 13 ][ 179 ],
   alphaCSR[ 13 ][ 180 ],
   alphaCSR[ 13 ][ 181 ],
   alphaCSR[ 13 ][ 182 ],
   alphaCSR[ 13 ][ 183 ],
   alphaCSR[ 13 ][ 184 ],
   alphaCSR[ 13 ][ 185 ],
   alphaCSR[ 13 ][ 186 ],
   alphaCSR[ 13 ][ 187 ],
   alphaCSR[ 13 ][ 188 ],
   alphaCSR[ 13 ][ 189 ],
   alphaCSR[ 13 ][ 190 ],
   alphaCSR[ 13 ][ 191 ],
   alphaCSR[ 13 ][ 192 ],
   alphaCSR[ 13 ][ 193 ],
   alphaCSR[ 13 ][ 194 ],
   alphaCSR[ 13 ][ 195 ],
   alphaCSR[ 13 ][ 196 ],
   alphaCSR[ 13 ][ 197 ],
   alphaCSR[ 13 ][ 198 ],
   alphaCSR[ 13 ][ 199 ],
   alphaCSR[ 13 ][ 200 ],
   alphaCSR[ 13 ][ 201 ],
   alphaCSR[ 13 ][ 202 ],
   alphaCSR[ 13 ][ 203 ],
   alphaCSR[ 13 ][ 204 ],
   alphaCSR[ 13 ][ 205 ],
   alphaCSR[ 13 ][ 206 ],
   alphaCSR[ 13 ][ 207 ],
   alphaCSR[ 13 ][ 208 ],
   alphaCSR[ 13 ][ 209 ],
   alphaCSR[ 13 ][ 210 ],
   alphaCSR[ 13 ][ 211 ],
   alphaCSR[ 13 ][ 212 ],
   alphaCSR[ 13 ][ 213 ],
   alphaCSR[ 13 ][ 214 ],
   alphaCSR[ 13 ][ 215 ],
   alphaCSR[ 13 ][ 216 ],
   alphaCSR[ 13 ][ 217 ],
   alphaCSR[ 13 ][ 218 ],
   alphaCSR[ 13 ][ 219 ],
   alphaCSR[ 13 ][ 220 ],
   alphaCSR[ 13 ][ 221 ],
   alphaCSR[ 13 ][ 222 ],
   alphaCSR[ 13 ][ 223 ],
   alphaCSR[ 13 ][ 224 ],
   alphaCSR[ 13 ][ 225 ],
   alphaCSR[ 13 ][ 226 ],
   alphaCSR[ 13 ][ 227 ],
   alphaCSR[ 13 ][ 228 ],
   alphaCSR[ 13 ][ 229 ],
   alphaCSR[ 13 ][ 230 ],
   alphaCSR[ 13 ][ 231 ],
   alphaCSR[ 13 ][ 232 ],
   alphaCSR[ 13 ][ 233 ],
   alphaCSR[ 13 ][ 234 ],
   alphaCSR[ 13 ][ 235 ],
   alphaCSR[ 13 ][ 236 ],
   alphaCSR[ 13 ][ 237 ],
   alphaCSR[ 13 ][ 238 ],
   alphaCSR[ 13 ][ 239 ],
   alphaCSR[ 13 ][ 240 ],
   alphaCSR[ 13 ][ 241 ],
   alphaCSR[ 13 ][ 242 ],
   alphaCSR[ 13 ][ 243 ],
   alphaCSR[ 13 ][ 244 ],
   alphaCSR[ 13 ][ 245 ],
   alphaCSR[ 13 ][ 246 ],
   alphaCSR[ 13 ][ 247 ],
   alphaCSR[ 13 ][ 248 ],
   alphaCSR[ 13 ][ 249 ],
   alphaCSR[ 13 ][ 250 ],
   alphaCSR[ 13 ][ 251 ],
   alphaCSR[ 13 ][ 252 ],
   alphaCSR[ 13 ][ 253 ],
   alphaCSR[ 13 ][ 254 ],
   alphaCSR[ 13 ][ 255 ],
   alphaCSR[ 13 ][ 256 ],
   alphaCSR[ 13 ][ 257 ],
   alphaCSR[ 13 ][ 258 ],
   alphaCSR[ 13 ][ 259 ],
   alphaCSR[ 13 ][ 260 ],
   alphaCSR[ 13 ][ 261 ],
   alphaCSR[ 13 ][ 262 ],
   alphaCSR[ 13 ][ 263 ],
   alphaCSR[ 13 ][ 264 ],
   alphaCSR[ 13 ][ 265 ],
   alphaCSR[ 13 ][ 266 ],
   alphaCSR[ 13 ][ 267 ],
   alphaCSR[ 13 ][ 268 ],
   alphaCSR[ 13 ][ 269 ],
   alphaCSR[ 13 ][ 270 ],
   alphaCSR[ 13 ][ 271 ],
   alphaCSR[ 13 ][ 272 ],
   alphaCSR[ 13 ][ 273 ],
   alphaCSR[ 13 ][ 274 ],
   alphaCSR[ 13 ][ 275 ],
   alphaCSR[ 13 ][ 276 ],
   alphaCSR[ 13 ][ 277 ],
   alphaCSR[ 13 ][ 278 ],
   alphaCSR[ 13 ][ 279 ],
   alphaCSR[ 13 ][ 280 ],
   alphaCSR[ 13 ][ 281 ],
   alphaCSR[ 13 ][ 282 ],
   alphaCSR[ 13 ][ 283 ],
   alphaCSR[ 13 ][ 284 ],
   alphaCSR[ 13 ][ 285 ],
   alphaCSR[ 13 ][ 286 ],
   alphaCSR[ 13 ][ 287 ],
   alphaCSR[ 13 ][ 288 ],
   alphaCSR[ 13 ][ 289 ],
   alphaCSR[ 13 ][ 290 ],
   alphaCSR[ 13 ][ 291 ],
   alphaCSR[ 13 ][ 292 ],
   alphaCSR[ 13 ][ 293 ],
   alphaCSR[ 13 ][ 294 ],
   alphaCSR[ 13 ][ 295 ],
   alphaCSR[ 13 ][ 296 ],
   alphaCSR[ 13 ][ 297 ],
   alphaCSR[ 13 ][ 298 ],
   alphaCSR[ 13 ][ 299 ],
   alphaCSR[ 13 ][ 300 ],
   alphaCSR[ 13 ][ 301 ],
   alphaCSR[ 13 ][ 302 ],
   alphaCSR[ 13 ][ 303 ],
   alphaCSR[ 13 ][ 304 ],
   alphaCSR[ 13 ][ 305 ],
   alphaCSR[ 13 ][ 306 ],
   alphaCSR[ 13 ][ 307 ],
   alphaCSR[ 13 ][ 308 ],
   alphaCSR[ 13 ][ 309 ],
   alphaCSR[ 13 ][ 310 ],
   alphaCSR[ 13 ][ 311 ],
   alphaCSR[ 13 ][ 312 ],
   alphaCSR[ 13 ][ 313 ],
   alphaCSR[ 13 ][ 314 ],
   alphaCSR[ 13 ][ 315 ],
   alphaCSR[ 13 ][ 316 ],
   alphaCSR[ 13 ][ 317 ],
   alphaCSR[ 13 ][ 318 ],
   alphaCSR[ 13 ][ 319 ],
   alphaCSR[ 13 ][ 320 ],
   alphaCSR[ 13 ][ 321 ],
   alphaCSR[ 13 ][ 322 ],
   alphaCSR[ 13 ][ 323 ],
   alphaCSR[ 13 ][ 324 ],
   alphaCSR[ 13 ][ 325 ],
   alphaCSR[ 13 ][ 326 ],
   alphaCSR[ 13 ][ 327 ],
   alphaCSR[ 13 ][ 328 ],
   alphaCSR[ 13 ][ 329 ],
   alphaCSR[ 13 ][ 330 ],
   alphaCSR[ 13 ][ 331 ],
   alphaCSR[ 13 ][ 332 ],
   alphaCSR[ 13 ][ 333 ],
   alphaCSR[ 13 ][ 334 ],
   alphaCSR[ 13 ][ 335 ],
   alphaCSR[ 13 ][ 336 ],
   alphaCSR[ 13 ][ 337 ],
   alphaCSR[ 13 ][ 338 ],
   alphaCSR[ 13 ][ 339 ],
   alphaCSR[ 13 ][ 340 ],
   alphaCSR[ 13 ][ 341 ],
   alphaCSR[ 13 ][ 342 ],
   alphaCSR[ 13 ][ 343 ],
   alphaCSR[ 13 ][ 344 ],
   alphaCSR[ 13 ][ 345 ],
   alphaCSR[ 13 ][ 346 ],
   alphaCSR[ 13 ][ 347 ],
   alphaCSR[ 13 ][ 348 ],
   alphaCSR[ 13 ][ 349 ],
   alphaCSR[ 13 ][ 350 ],
   alphaCSR[ 13 ][ 351 ],
   alphaCSR[ 13 ][ 352 ],
   alphaCSR[ 13 ][ 353 ],
   alphaCSR[ 13 ][ 354 ],
   alphaCSR[ 13 ][ 355 ],
   alphaCSR[ 13 ][ 356 ],
   alphaCSR[ 13 ][ 357 ],
   alphaCSR[ 13 ][ 358 ],
   alphaCSR[ 13 ][ 359 ],
   alphaCSR[ 13 ][ 360 ],
   alphaCSR[ 13 ][ 361 ],
   alphaCSR[ 13 ][ 362 ],
   alphaCSR[ 13 ][ 363 ],
   alphaCSR[ 13 ][ 364 ],
   alphaCSR[ 13 ][ 365 ],
   alphaCSR[ 13 ][ 366 ],
   alphaCSR[ 13 ][ 367 ],
   alphaCSR[ 13 ][ 368 ],
   alphaCSR[ 13 ][ 369 ],
   alphaCSR[ 13 ][ 370 ],
   alphaCSR[ 13 ][ 371 ],
   alphaCSR[ 13 ][ 372 ],
   alphaCSR[ 13 ][ 373 ],
   alphaCSR[ 13 ][ 374 ],
   alphaCSR[ 13 ][ 375 ],
   alphaCSR[ 13 ][ 376 ],
   alphaCSR[ 13 ][ 377 ],
   alphaCSR[ 13 ][ 378 ],
   alphaCSR[ 13 ][ 379 ],
   alphaCSR[ 13 ][ 380 ],
   alphaCSR[ 13 ][ 381 ],
   alphaCSR[ 13 ][ 382 ],
   alphaCSR[ 13 ][ 383 ],
   alphaCSR[ 14 ][ 0 ],
   alphaCSR[ 14 ][ 1 ],
   alphaCSR[ 14 ][ 2 ],
   alphaCSR[ 14 ][ 3 ],
   alphaCSR[ 14 ][ 4 ],
   alphaCSR[ 14 ][ 5 ],
   alphaCSR[ 14 ][ 6 ],
   alphaCSR[ 14 ][ 7 ],
   alphaCSR[ 14 ][ 8 ],
   alphaCSR[ 14 ][ 9 ],
   alphaCSR[ 14 ][ 10 ],
   alphaCSR[ 14 ][ 11 ],
   alphaCSR[ 14 ][ 12 ],
   alphaCSR[ 14 ][ 13 ],
   alphaCSR[ 14 ][ 14 ],
   alphaCSR[ 14 ][ 15 ],
   alphaCSR[ 14 ][ 16 ],
   alphaCSR[ 14 ][ 17 ],
   alphaCSR[ 14 ][ 18 ],
   alphaCSR[ 14 ][ 19 ],
   alphaCSR[ 14 ][ 20 ],
   alphaCSR[ 14 ][ 21 ],
   alphaCSR[ 14 ][ 22 ],
   alphaCSR[ 14 ][ 23 ],
   alphaCSR[ 14 ][ 24 ],
   alphaCSR[ 14 ][ 25 ],
   alphaCSR[ 14 ][ 26 ],
   alphaCSR[ 14 ][ 27 ],
   alphaCSR[ 14 ][ 28 ],
   alphaCSR[ 14 ][ 29 ],
   alphaCSR[ 14 ][ 30 ],
   alphaCSR[ 14 ][ 31 ],
   alphaCSR[ 14 ][ 32 ],
   alphaCSR[ 14 ][ 33 ],
   alphaCSR[ 14 ][ 34 ],
   alphaCSR[ 14 ][ 35 ],
   alphaCSR[ 14 ][ 36 ],
   alphaCSR[ 14 ][ 37 ],
   alphaCSR[ 14 ][ 38 ],
   alphaCSR[ 14 ][ 39 ],
   alphaCSR[ 14 ][ 40 ],
   alphaCSR[ 14 ][ 41 ],
   alphaCSR[ 14 ][ 42 ],
   alphaCSR[ 14 ][ 43 ],
   alphaCSR[ 14 ][ 44 ],
   alphaCSR[ 14 ][ 45 ],
   alphaCSR[ 14 ][ 46 ],
   alphaCSR[ 14 ][ 47 ],
   alphaCSR[ 14 ][ 48 ],
   alphaCSR[ 14 ][ 49 ],
   alphaCSR[ 14 ][ 50 ],
   alphaCSR[ 14 ][ 51 ],
   alphaCSR[ 14 ][ 52 ],
   alphaCSR[ 14 ][ 53 ],
   alphaCSR[ 14 ][ 54 ],
   alphaCSR[ 14 ][ 55 ],
   alphaCSR[ 14 ][ 56 ],
   alphaCSR[ 14 ][ 57 ],
   alphaCSR[ 14 ][ 58 ],
   alphaCSR[ 14 ][ 59 ],
   alphaCSR[ 14 ][ 60 ],
   alphaCSR[ 14 ][ 61 ],
   alphaCSR[ 14 ][ 62 ],
   alphaCSR[ 14 ][ 63 ],
   alphaCSR[ 14 ][ 64 ],
   alphaCSR[ 14 ][ 65 ],
   alphaCSR[ 14 ][ 66 ],
   alphaCSR[ 14 ][ 67 ],
   alphaCSR[ 14 ][ 68 ],
   alphaCSR[ 14 ][ 69 ],
   alphaCSR[ 14 ][ 70 ],
   alphaCSR[ 14 ][ 71 ],
   alphaCSR[ 14 ][ 72 ],
   alphaCSR[ 14 ][ 73 ],
   alphaCSR[ 14 ][ 74 ],
   alphaCSR[ 14 ][ 75 ],
   alphaCSR[ 14 ][ 76 ],
   alphaCSR[ 14 ][ 77 ],
   alphaCSR[ 14 ][ 78 ],
   alphaCSR[ 14 ][ 79 ],
   alphaCSR[ 14 ][ 80 ],
   alphaCSR[ 14 ][ 81 ],
   alphaCSR[ 14 ][ 82 ],
   alphaCSR[ 14 ][ 83 ],
   alphaCSR[ 14 ][ 84 ],
   alphaCSR[ 14 ][ 85 ],
   alphaCSR[ 14 ][ 86 ],
   alphaCSR[ 14 ][ 87 ],
   alphaCSR[ 14 ][ 88 ],
   alphaCSR[ 14 ][ 89 ],
   alphaCSR[ 14 ][ 90 ],
   alphaCSR[ 14 ][ 91 ],
   alphaCSR[ 14 ][ 92 ],
   alphaCSR[ 14 ][ 93 ],
   alphaCSR[ 14 ][ 94 ],
   alphaCSR[ 14 ][ 95 ],
   alphaCSR[ 14 ][ 96 ],
   alphaCSR[ 14 ][ 97 ],
   alphaCSR[ 14 ][ 98 ],
   alphaCSR[ 14 ][ 99 ],
   alphaCSR[ 14 ][ 100 ],
   alphaCSR[ 14 ][ 101 ],
   alphaCSR[ 14 ][ 102 ],
   alphaCSR[ 14 ][ 103 ],
   alphaCSR[ 14 ][ 104 ],
   alphaCSR[ 14 ][ 105 ],
   alphaCSR[ 14 ][ 106 ],
   alphaCSR[ 14 ][ 107 ],
   alphaCSR[ 14 ][ 108 ],
   alphaCSR[ 14 ][ 109 ],
   alphaCSR[ 14 ][ 110 ],
   alphaCSR[ 14 ][ 111 ],
   alphaCSR[ 14 ][ 112 ],
   alphaCSR[ 14 ][ 113 ],
   alphaCSR[ 14 ][ 114 ],
   alphaCSR[ 14 ][ 115 ],
   alphaCSR[ 14 ][ 116 ],
   alphaCSR[ 14 ][ 117 ],
   alphaCSR[ 14 ][ 118 ],
   alphaCSR[ 14 ][ 119 ],
   alphaCSR[ 14 ][ 120 ],
   alphaCSR[ 14 ][ 121 ],
   alphaCSR[ 14 ][ 122 ],
   alphaCSR[ 14 ][ 123 ],
   alphaCSR[ 14 ][ 124 ],
   alphaCSR[ 14 ][ 125 ],
   alphaCSR[ 14 ][ 126 ],
   alphaCSR[ 14 ][ 127 ],
   alphaCSR[ 14 ][ 128 ],
   alphaCSR[ 14 ][ 129 ],
   alphaCSR[ 14 ][ 130 ],
   alphaCSR[ 14 ][ 131 ],
   alphaCSR[ 14 ][ 132 ],
   alphaCSR[ 14 ][ 133 ],
   alphaCSR[ 14 ][ 134 ],
   alphaCSR[ 14 ][ 135 ],
   alphaCSR[ 14 ][ 136 ],
   alphaCSR[ 14 ][ 137 ],
   alphaCSR[ 14 ][ 138 ],
   alphaCSR[ 14 ][ 139 ],
   alphaCSR[ 14 ][ 140 ],
   alphaCSR[ 14 ][ 141 ],
   alphaCSR[ 14 ][ 142 ],
   alphaCSR[ 14 ][ 143 ],
   alphaCSR[ 14 ][ 144 ],
   alphaCSR[ 14 ][ 145 ],
   alphaCSR[ 14 ][ 146 ],
   alphaCSR[ 14 ][ 147 ],
   alphaCSR[ 14 ][ 148 ],
   alphaCSR[ 14 ][ 149 ],
   alphaCSR[ 14 ][ 150 ],
   alphaCSR[ 14 ][ 151 ],
   alphaCSR[ 14 ][ 152 ],
   alphaCSR[ 14 ][ 153 ],
   alphaCSR[ 14 ][ 154 ],
   alphaCSR[ 14 ][ 155 ],
   alphaCSR[ 14 ][ 156 ],
   alphaCSR[ 14 ][ 157 ],
   alphaCSR[ 14 ][ 158 ],
   alphaCSR[ 14 ][ 159 ],
   alphaCSR[ 14 ][ 160 ],
   alphaCSR[ 14 ][ 161 ],
   alphaCSR[ 14 ][ 162 ],
   alphaCSR[ 14 ][ 163 ],
   alphaCSR[ 14 ][ 164 ],
   alphaCSR[ 14 ][ 165 ],
   alphaCSR[ 14 ][ 166 ],
   alphaCSR[ 14 ][ 167 ],
   alphaCSR[ 14 ][ 168 ],
   alphaCSR[ 14 ][ 169 ],
   alphaCSR[ 14 ][ 170 ],
   alphaCSR[ 14 ][ 171 ],
   alphaCSR[ 14 ][ 172 ],
   alphaCSR[ 14 ][ 173 ],
   alphaCSR[ 14 ][ 174 ],
   alphaCSR[ 14 ][ 175 ],
   alphaCSR[ 14 ][ 176 ],
   alphaCSR[ 14 ][ 177 ],
   alphaCSR[ 14 ][ 178 ],
   alphaCSR[ 14 ][ 179 ],
   alphaCSR[ 14 ][ 180 ],
   alphaCSR[ 14 ][ 181 ],
   alphaCSR[ 14 ][ 182 ],
   alphaCSR[ 14 ][ 183 ],
   alphaCSR[ 14 ][ 184 ],
   alphaCSR[ 14 ][ 185 ],
   alphaCSR[ 14 ][ 186 ],
   alphaCSR[ 14 ][ 187 ],
   alphaCSR[ 14 ][ 188 ],
   alphaCSR[ 14 ][ 189 ],
   alphaCSR[ 14 ][ 190 ],
   alphaCSR[ 14 ][ 191 ],
   alphaCSR[ 14 ][ 192 ],
   alphaCSR[ 14 ][ 193 ],
   alphaCSR[ 14 ][ 194 ],
   alphaCSR[ 14 ][ 195 ],
   alphaCSR[ 14 ][ 196 ],
   alphaCSR[ 14 ][ 197 ],
   alphaCSR[ 14 ][ 198 ],
   alphaCSR[ 14 ][ 199 ],
   alphaCSR[ 14 ][ 200 ],
   alphaCSR[ 14 ][ 201 ],
   alphaCSR[ 14 ][ 202 ],
   alphaCSR[ 14 ][ 203 ],
   alphaCSR[ 14 ][ 204 ],
   alphaCSR[ 14 ][ 205 ],
   alphaCSR[ 14 ][ 206 ],
   alphaCSR[ 14 ][ 207 ],
   alphaCSR[ 14 ][ 208 ],
   alphaCSR[ 14 ][ 209 ],
   alphaCSR[ 14 ][ 210 ],
   alphaCSR[ 14 ][ 211 ],
   alphaCSR[ 14 ][ 212 ],
   alphaCSR[ 14 ][ 213 ],
   alphaCSR[ 14 ][ 214 ],
   alphaCSR[ 14 ][ 215 ],
   alphaCSR[ 14 ][ 216 ],
   alphaCSR[ 14 ][ 217 ],
   alphaCSR[ 14 ][ 218 ],
   alphaCSR[ 14 ][ 219 ],
   alphaCSR[ 14 ][ 220 ],
   alphaCSR[ 14 ][ 221 ],
   alphaCSR[ 14 ][ 222 ],
   alphaCSR[ 14 ][ 223 ],
   alphaCSR[ 14 ][ 224 ],
   alphaCSR[ 14 ][ 225 ],
   alphaCSR[ 14 ][ 226 ],
   alphaCSR[ 14 ][ 227 ],
   alphaCSR[ 14 ][ 228 ],
   alphaCSR[ 14 ][ 229 ],
   alphaCSR[ 14 ][ 230 ],
   alphaCSR[ 14 ][ 231 ],
   alphaCSR[ 14 ][ 232 ],
   alphaCSR[ 14 ][ 233 ],
   alphaCSR[ 14 ][ 234 ],
   alphaCSR[ 14 ][ 235 ],
   alphaCSR[ 14 ][ 236 ],
   alphaCSR[ 14 ][ 237 ],
   alphaCSR[ 14 ][ 238 ],
   alphaCSR[ 14 ][ 239 ],
   alphaCSR[ 14 ][ 240 ],
   alphaCSR[ 14 ][ 241 ],
   alphaCSR[ 14 ][ 242 ],
   alphaCSR[ 14 ][ 243 ],
   alphaCSR[ 14 ][ 244 ],
   alphaCSR[ 14 ][ 245 ],
   alphaCSR[ 14 ][ 246 ],
   alphaCSR[ 14 ][ 247 ],
   alphaCSR[ 14 ][ 248 ],
   alphaCSR[ 14 ][ 249 ],
   alphaCSR[ 14 ][ 250 ],
   alphaCSR[ 14 ][ 251 ],
   alphaCSR[ 14 ][ 252 ],
   alphaCSR[ 14 ][ 253 ],
   alphaCSR[ 14 ][ 254 ],
   alphaCSR[ 14 ][ 255 ],
   alphaCSR[ 14 ][ 256 ],
   alphaCSR[ 14 ][ 257 ],
   alphaCSR[ 14 ][ 258 ],
   alphaCSR[ 14 ][ 259 ],
   alphaCSR[ 14 ][ 260 ],
   alphaCSR[ 14 ][ 261 ],
   alphaCSR[ 14 ][ 262 ],
   alphaCSR[ 14 ][ 263 ],
   alphaCSR[ 14 ][ 264 ],
   alphaCSR[ 14 ][ 265 ],
   alphaCSR[ 14 ][ 266 ],
   alphaCSR[ 14 ][ 267 ],
   alphaCSR[ 14 ][ 268 ],
   alphaCSR[ 14 ][ 269 ],
   alphaCSR[ 14 ][ 270 ],
   alphaCSR[ 14 ][ 271 ],
   alphaCSR[ 14 ][ 272 ],
   alphaCSR[ 14 ][ 273 ],
   alphaCSR[ 14 ][ 274 ],
   alphaCSR[ 14 ][ 275 ],
   alphaCSR[ 14 ][ 276 ],
   alphaCSR[ 14 ][ 277 ],
   alphaCSR[ 14 ][ 278 ],
   alphaCSR[ 14 ][ 279 ],
   alphaCSR[ 14 ][ 280 ],
   alphaCSR[ 14 ][ 281 ],
   alphaCSR[ 14 ][ 282 ],
   alphaCSR[ 14 ][ 283 ],
   alphaCSR[ 14 ][ 284 ],
   alphaCSR[ 14 ][ 285 ],
   alphaCSR[ 14 ][ 286 ],
   alphaCSR[ 14 ][ 287 ],
   alphaCSR[ 14 ][ 288 ],
   alphaCSR[ 14 ][ 289 ],
   alphaCSR[ 14 ][ 290 ],
   alphaCSR[ 14 ][ 291 ],
   alphaCSR[ 14 ][ 292 ],
   alphaCSR[ 14 ][ 293 ],
   alphaCSR[ 14 ][ 294 ],
   alphaCSR[ 14 ][ 295 ],
   alphaCSR[ 14 ][ 296 ],
   alphaCSR[ 14 ][ 297 ],
   alphaCSR[ 14 ][ 298 ],
   alphaCSR[ 14 ][ 299 ],
   alphaCSR[ 14 ][ 300 ],
   alphaCSR[ 14 ][ 301 ],
   alphaCSR[ 14 ][ 302 ],
   alphaCSR[ 14 ][ 303 ],
   alphaCSR[ 14 ][ 304 ],
   alphaCSR[ 14 ][ 305 ],
   alphaCSR[ 14 ][ 306 ],
   alphaCSR[ 14 ][ 307 ],
   alphaCSR[ 14 ][ 308 ],
   alphaCSR[ 14 ][ 309 ],
   alphaCSR[ 14 ][ 310 ],
   alphaCSR[ 14 ][ 311 ],
   alphaCSR[ 14 ][ 312 ],
   alphaCSR[ 14 ][ 313 ],
   alphaCSR[ 14 ][ 314 ],
   alphaCSR[ 14 ][ 315 ],
   alphaCSR[ 14 ][ 316 ],
   alphaCSR[ 14 ][ 317 ],
   alphaCSR[ 14 ][ 318 ],
   alphaCSR[ 14 ][ 319 ],
   alphaCSR[ 14 ][ 320 ],
   alphaCSR[ 14 ][ 321 ],
   alphaCSR[ 14 ][ 322 ],
   alphaCSR[ 14 ][ 323 ],
   alphaCSR[ 14 ][ 324 ],
   alphaCSR[ 14 ][ 325 ],
   alphaCSR[ 14 ][ 326 ],
   alphaCSR[ 14 ][ 327 ],
   alphaCSR[ 14 ][ 328 ],
   alphaCSR[ 14 ][ 329 ],
   alphaCSR[ 14 ][ 330 ],
   alphaCSR[ 14 ][ 331 ],
   alphaCSR[ 14 ][ 332 ],
   alphaCSR[ 14 ][ 333 ],
   alphaCSR[ 14 ][ 334 ],
   alphaCSR[ 14 ][ 335 ],
   alphaCSR[ 14 ][ 336 ],
   alphaCSR[ 14 ][ 337 ],
   alphaCSR[ 14 ][ 338 ],
   alphaCSR[ 14 ][ 339 ],
   alphaCSR[ 14 ][ 340 ],
   alphaCSR[ 14 ][ 341 ],
   alphaCSR[ 14 ][ 342 ],
   alphaCSR[ 14 ][ 343 ],
   alphaCSR[ 14 ][ 344 ],
   alphaCSR[ 14 ][ 345 ],
   alphaCSR[ 14 ][ 346 ],
   alphaCSR[ 14 ][ 347 ],
   alphaCSR[ 14 ][ 348 ],
   alphaCSR[ 14 ][ 349 ],
   alphaCSR[ 14 ][ 350 ],
   alphaCSR[ 14 ][ 351 ],
   alphaCSR[ 14 ][ 352 ],
   alphaCSR[ 14 ][ 353 ],
   alphaCSR[ 14 ][ 354 ],
   alphaCSR[ 14 ][ 355 ],
   alphaCSR[ 14 ][ 356 ],
   alphaCSR[ 14 ][ 357 ],
   alphaCSR[ 14 ][ 358 ],
   alphaCSR[ 14 ][ 359 ],
   alphaCSR[ 14 ][ 360 ],
   alphaCSR[ 14 ][ 361 ],
   alphaCSR[ 14 ][ 362 ],
   alphaCSR[ 14 ][ 363 ],
   alphaCSR[ 14 ][ 364 ],
   alphaCSR[ 14 ][ 365 ],
   alphaCSR[ 14 ][ 366 ],
   alphaCSR[ 14 ][ 367 ],
   alphaCSR[ 14 ][ 368 ],
   alphaCSR[ 14 ][ 369 ],
   alphaCSR[ 14 ][ 370 ],
   alphaCSR[ 14 ][ 371 ],
   alphaCSR[ 14 ][ 372 ],
   alphaCSR[ 14 ][ 373 ],
   alphaCSR[ 14 ][ 374 ],
   alphaCSR[ 14 ][ 375 ],
   alphaCSR[ 14 ][ 376 ],
   alphaCSR[ 14 ][ 377 ],
   alphaCSR[ 14 ][ 378 ],
   alphaCSR[ 14 ][ 379 ],
   alphaCSR[ 14 ][ 380 ],
   alphaCSR[ 14 ][ 381 ],
   alphaCSR[ 14 ][ 382 ],
   alphaCSR[ 14 ][ 383 ],
   alphaCSR[ 15 ][ 0 ],
   alphaCSR[ 15 ][ 1 ],
   alphaCSR[ 15 ][ 2 ],
   alphaCSR[ 15 ][ 3 ],
   alphaCSR[ 15 ][ 4 ],
   alphaCSR[ 15 ][ 5 ],
   alphaCSR[ 15 ][ 6 ],
   alphaCSR[ 15 ][ 7 ],
   alphaCSR[ 15 ][ 8 ],
   alphaCSR[ 15 ][ 9 ],
   alphaCSR[ 15 ][ 10 ],
   alphaCSR[ 15 ][ 11 ],
   alphaCSR[ 15 ][ 12 ],
   alphaCSR[ 15 ][ 13 ],
   alphaCSR[ 15 ][ 14 ],
   alphaCSR[ 15 ][ 15 ],
   alphaCSR[ 15 ][ 16 ],
   alphaCSR[ 15 ][ 17 ],
   alphaCSR[ 15 ][ 18 ],
   alphaCSR[ 15 ][ 19 ],
   alphaCSR[ 15 ][ 20 ],
   alphaCSR[ 15 ][ 21 ],
   alphaCSR[ 15 ][ 22 ],
   alphaCSR[ 15 ][ 23 ],
   alphaCSR[ 15 ][ 24 ],
   alphaCSR[ 15 ][ 25 ],
   alphaCSR[ 15 ][ 26 ],
   alphaCSR[ 15 ][ 27 ],
   alphaCSR[ 15 ][ 28 ],
   alphaCSR[ 15 ][ 29 ],
   alphaCSR[ 15 ][ 30 ],
   alphaCSR[ 15 ][ 31 ],
   alphaCSR[ 15 ][ 32 ],
   alphaCSR[ 15 ][ 33 ],
   alphaCSR[ 15 ][ 34 ],
   alphaCSR[ 15 ][ 35 ],
   alphaCSR[ 15 ][ 36 ],
   alphaCSR[ 15 ][ 37 ],
   alphaCSR[ 15 ][ 38 ],
   alphaCSR[ 15 ][ 39 ],
   alphaCSR[ 15 ][ 40 ],
   alphaCSR[ 15 ][ 41 ],
   alphaCSR[ 15 ][ 42 ],
   alphaCSR[ 15 ][ 43 ],
   alphaCSR[ 15 ][ 44 ],
   alphaCSR[ 15 ][ 45 ],
   alphaCSR[ 15 ][ 46 ],
   alphaCSR[ 15 ][ 47 ],
   alphaCSR[ 15 ][ 48 ],
   alphaCSR[ 15 ][ 49 ],
   alphaCSR[ 15 ][ 50 ],
   alphaCSR[ 15 ][ 51 ],
   alphaCSR[ 15 ][ 52 ],
   alphaCSR[ 15 ][ 53 ],
   alphaCSR[ 15 ][ 54 ],
   alphaCSR[ 15 ][ 55 ],
   alphaCSR[ 15 ][ 56 ],
   alphaCSR[ 15 ][ 57 ],
   alphaCSR[ 15 ][ 58 ],
   alphaCSR[ 15 ][ 59 ],
   alphaCSR[ 15 ][ 60 ],
   alphaCSR[ 15 ][ 61 ],
   alphaCSR[ 15 ][ 62 ],
   alphaCSR[ 15 ][ 63 ],
   alphaCSR[ 15 ][ 64 ],
   alphaCSR[ 15 ][ 65 ],
   alphaCSR[ 15 ][ 66 ],
   alphaCSR[ 15 ][ 67 ],
   alphaCSR[ 15 ][ 68 ],
   alphaCSR[ 15 ][ 69 ],
   alphaCSR[ 15 ][ 70 ],
   alphaCSR[ 15 ][ 71 ],
   alphaCSR[ 15 ][ 72 ],
   alphaCSR[ 15 ][ 73 ],
   alphaCSR[ 15 ][ 74 ],
   alphaCSR[ 15 ][ 75 ],
   alphaCSR[ 15 ][ 76 ],
   alphaCSR[ 15 ][ 77 ],
   alphaCSR[ 15 ][ 78 ],
   alphaCSR[ 15 ][ 79 ],
   alphaCSR[ 15 ][ 80 ],
   alphaCSR[ 15 ][ 81 ],
   alphaCSR[ 15 ][ 82 ],
   alphaCSR[ 15 ][ 83 ],
   alphaCSR[ 15 ][ 84 ],
   alphaCSR[ 15 ][ 85 ],
   alphaCSR[ 15 ][ 86 ],
   alphaCSR[ 15 ][ 87 ],
   alphaCSR[ 15 ][ 88 ],
   alphaCSR[ 15 ][ 89 ],
   alphaCSR[ 15 ][ 90 ],
   alphaCSR[ 15 ][ 91 ],
   alphaCSR[ 15 ][ 92 ],
   alphaCSR[ 15 ][ 93 ],
   alphaCSR[ 15 ][ 94 ],
   alphaCSR[ 15 ][ 95 ],
   alphaCSR[ 15 ][ 96 ],
   alphaCSR[ 15 ][ 97 ],
   alphaCSR[ 15 ][ 98 ],
   alphaCSR[ 15 ][ 99 ],
   alphaCSR[ 15 ][ 100 ],
   alphaCSR[ 15 ][ 101 ],
   alphaCSR[ 15 ][ 102 ],
   alphaCSR[ 15 ][ 103 ],
   alphaCSR[ 15 ][ 104 ],
   alphaCSR[ 15 ][ 105 ],
   alphaCSR[ 15 ][ 106 ],
   alphaCSR[ 15 ][ 107 ],
   alphaCSR[ 15 ][ 108 ],
   alphaCSR[ 15 ][ 109 ],
   alphaCSR[ 15 ][ 110 ],
   alphaCSR[ 15 ][ 111 ],
   alphaCSR[ 15 ][ 112 ],
   alphaCSR[ 15 ][ 113 ],
   alphaCSR[ 15 ][ 114 ],
   alphaCSR[ 15 ][ 115 ],
   alphaCSR[ 15 ][ 116 ],
   alphaCSR[ 15 ][ 117 ],
   alphaCSR[ 15 ][ 118 ],
   alphaCSR[ 15 ][ 119 ],
   alphaCSR[ 15 ][ 120 ],
   alphaCSR[ 15 ][ 121 ],
   alphaCSR[ 15 ][ 122 ],
   alphaCSR[ 15 ][ 123 ],
   alphaCSR[ 15 ][ 124 ],
   alphaCSR[ 15 ][ 125 ],
   alphaCSR[ 15 ][ 126 ],
   alphaCSR[ 15 ][ 127 ],
   alphaCSR[ 15 ][ 128 ],
   alphaCSR[ 15 ][ 129 ],
   alphaCSR[ 15 ][ 130 ],
   alphaCSR[ 15 ][ 131 ],
   alphaCSR[ 15 ][ 132 ],
   alphaCSR[ 15 ][ 133 ],
   alphaCSR[ 15 ][ 134 ],
   alphaCSR[ 15 ][ 135 ],
   alphaCSR[ 15 ][ 136 ],
   alphaCSR[ 15 ][ 137 ],
   alphaCSR[ 15 ][ 138 ],
   alphaCSR[ 15 ][ 139 ],
   alphaCSR[ 15 ][ 140 ],
   alphaCSR[ 15 ][ 141 ],
   alphaCSR[ 15 ][ 142 ],
   alphaCSR[ 15 ][ 143 ],
   alphaCSR[ 15 ][ 144 ],
   alphaCSR[ 15 ][ 145 ],
   alphaCSR[ 15 ][ 146 ],
   alphaCSR[ 15 ][ 147 ],
   alphaCSR[ 15 ][ 148 ],
   alphaCSR[ 15 ][ 149 ],
   alphaCSR[ 15 ][ 150 ],
   alphaCSR[ 15 ][ 151 ],
   alphaCSR[ 15 ][ 152 ],
   alphaCSR[ 15 ][ 153 ],
   alphaCSR[ 15 ][ 154 ],
   alphaCSR[ 15 ][ 155 ],
   alphaCSR[ 15 ][ 156 ],
   alphaCSR[ 15 ][ 157 ],
   alphaCSR[ 15 ][ 158 ],
   alphaCSR[ 15 ][ 159 ],
   alphaCSR[ 15 ][ 160 ],
   alphaCSR[ 15 ][ 161 ],
   alphaCSR[ 15 ][ 162 ],
   alphaCSR[ 15 ][ 163 ],
   alphaCSR[ 15 ][ 164 ],
   alphaCSR[ 15 ][ 165 ],
   alphaCSR[ 15 ][ 166 ],
   alphaCSR[ 15 ][ 167 ],
   alphaCSR[ 15 ][ 168 ],
   alphaCSR[ 15 ][ 169 ],
   alphaCSR[ 15 ][ 170 ],
   alphaCSR[ 15 ][ 171 ],
   alphaCSR[ 15 ][ 172 ],
   alphaCSR[ 15 ][ 173 ],
   alphaCSR[ 15 ][ 174 ],
   alphaCSR[ 15 ][ 175 ],
   alphaCSR[ 15 ][ 176 ],
   alphaCSR[ 15 ][ 177 ],
   alphaCSR[ 15 ][ 178 ],
   alphaCSR[ 15 ][ 179 ],
   alphaCSR[ 15 ][ 180 ],
   alphaCSR[ 15 ][ 181 ],
   alphaCSR[ 15 ][ 182 ],
   alphaCSR[ 15 ][ 183 ],
   alphaCSR[ 15 ][ 184 ],
   alphaCSR[ 15 ][ 185 ],
   alphaCSR[ 15 ][ 186 ],
   alphaCSR[ 15 ][ 187 ],
   alphaCSR[ 15 ][ 188 ],
   alphaCSR[ 15 ][ 189 ],
   alphaCSR[ 15 ][ 190 ],
   alphaCSR[ 15 ][ 191 ],
   alphaCSR[ 15 ][ 192 ],
   alphaCSR[ 15 ][ 193 ],
   alphaCSR[ 15 ][ 194 ],
   alphaCSR[ 15 ][ 195 ],
   alphaCSR[ 15 ][ 196 ],
   alphaCSR[ 15 ][ 197 ],
   alphaCSR[ 15 ][ 198 ],
   alphaCSR[ 15 ][ 199 ],
   alphaCSR[ 15 ][ 200 ],
   alphaCSR[ 15 ][ 201 ],
   alphaCSR[ 15 ][ 202 ],
   alphaCSR[ 15 ][ 203 ],
   alphaCSR[ 15 ][ 204 ],
   alphaCSR[ 15 ][ 205 ],
   alphaCSR[ 15 ][ 206 ],
   alphaCSR[ 15 ][ 207 ],
   alphaCSR[ 15 ][ 208 ],
   alphaCSR[ 15 ][ 209 ],
   alphaCSR[ 15 ][ 210 ],
   alphaCSR[ 15 ][ 211 ],
   alphaCSR[ 15 ][ 212 ],
   alphaCSR[ 15 ][ 213 ],
   alphaCSR[ 15 ][ 214 ],
   alphaCSR[ 15 ][ 215 ],
   alphaCSR[ 15 ][ 216 ],
   alphaCSR[ 15 ][ 217 ],
   alphaCSR[ 15 ][ 218 ],
   alphaCSR[ 15 ][ 219 ],
   alphaCSR[ 15 ][ 220 ],
   alphaCSR[ 15 ][ 221 ],
   alphaCSR[ 15 ][ 222 ],
   alphaCSR[ 15 ][ 223 ],
   alphaCSR[ 15 ][ 224 ],
   alphaCSR[ 15 ][ 225 ],
   alphaCSR[ 15 ][ 226 ],
   alphaCSR[ 15 ][ 227 ],
   alphaCSR[ 15 ][ 228 ],
   alphaCSR[ 15 ][ 229 ],
   alphaCSR[ 15 ][ 230 ],
   alphaCSR[ 15 ][ 231 ],
   alphaCSR[ 15 ][ 232 ],
   alphaCSR[ 15 ][ 233 ],
   alphaCSR[ 15 ][ 234 ],
   alphaCSR[ 15 ][ 235 ],
   alphaCSR[ 15 ][ 236 ],
   alphaCSR[ 15 ][ 237 ],
   alphaCSR[ 15 ][ 238 ],
   alphaCSR[ 15 ][ 239 ],
   alphaCSR[ 15 ][ 240 ],
   alphaCSR[ 15 ][ 241 ],
   alphaCSR[ 15 ][ 242 ],
   alphaCSR[ 15 ][ 243 ],
   alphaCSR[ 15 ][ 244 ],
   alphaCSR[ 15 ][ 245 ],
   alphaCSR[ 15 ][ 246 ],
   alphaCSR[ 15 ][ 247 ],
   alphaCSR[ 15 ][ 248 ],
   alphaCSR[ 15 ][ 249 ],
   alphaCSR[ 15 ][ 250 ],
   alphaCSR[ 15 ][ 251 ],
   alphaCSR[ 15 ][ 252 ],
   alphaCSR[ 15 ][ 253 ],
   alphaCSR[ 15 ][ 254 ],
   alphaCSR[ 15 ][ 255 ],
   alphaCSR[ 15 ][ 256 ],
   alphaCSR[ 15 ][ 257 ],
   alphaCSR[ 15 ][ 258 ],
   alphaCSR[ 15 ][ 259 ],
   alphaCSR[ 15 ][ 260 ],
   alphaCSR[ 15 ][ 261 ],
   alphaCSR[ 15 ][ 262 ],
   alphaCSR[ 15 ][ 263 ],
   alphaCSR[ 15 ][ 264 ],
   alphaCSR[ 15 ][ 265 ],
   alphaCSR[ 15 ][ 266 ],
   alphaCSR[ 15 ][ 267 ],
   alphaCSR[ 15 ][ 268 ],
   alphaCSR[ 15 ][ 269 ],
   alphaCSR[ 15 ][ 270 ],
   alphaCSR[ 15 ][ 271 ],
   alphaCSR[ 15 ][ 272 ],
   alphaCSR[ 15 ][ 273 ],
   alphaCSR[ 15 ][ 274 ],
   alphaCSR[ 15 ][ 275 ],
   alphaCSR[ 15 ][ 276 ],
   alphaCSR[ 15 ][ 277 ],
   alphaCSR[ 15 ][ 278 ],
   alphaCSR[ 15 ][ 279 ],
   alphaCSR[ 15 ][ 280 ],
   alphaCSR[ 15 ][ 281 ],
   alphaCSR[ 15 ][ 282 ],
   alphaCSR[ 15 ][ 283 ],
   alphaCSR[ 15 ][ 284 ],
   alphaCSR[ 15 ][ 285 ],
   alphaCSR[ 15 ][ 286 ],
   alphaCSR[ 15 ][ 287 ],
   alphaCSR[ 15 ][ 288 ],
   alphaCSR[ 15 ][ 289 ],
   alphaCSR[ 15 ][ 290 ],
   alphaCSR[ 15 ][ 291 ],
   alphaCSR[ 15 ][ 292 ],
   alphaCSR[ 15 ][ 293 ],
   alphaCSR[ 15 ][ 294 ],
   alphaCSR[ 15 ][ 295 ],
   alphaCSR[ 15 ][ 296 ],
   alphaCSR[ 15 ][ 297 ],
   alphaCSR[ 15 ][ 298 ],
   alphaCSR[ 15 ][ 299 ],
   alphaCSR[ 15 ][ 300 ],
   alphaCSR[ 15 ][ 301 ],
   alphaCSR[ 15 ][ 302 ],
   alphaCSR[ 15 ][ 303 ],
   alphaCSR[ 15 ][ 304 ],
   alphaCSR[ 15 ][ 305 ],
   alphaCSR[ 15 ][ 306 ],
   alphaCSR[ 15 ][ 307 ],
   alphaCSR[ 15 ][ 308 ],
   alphaCSR[ 15 ][ 309 ],
   alphaCSR[ 15 ][ 310 ],
   alphaCSR[ 15 ][ 311 ],
   alphaCSR[ 15 ][ 312 ],
   alphaCSR[ 15 ][ 313 ],
   alphaCSR[ 15 ][ 314 ],
   alphaCSR[ 15 ][ 315 ],
   alphaCSR[ 15 ][ 316 ],
   alphaCSR[ 15 ][ 317 ],
   alphaCSR[ 15 ][ 318 ],
   alphaCSR[ 15 ][ 319 ],
   alphaCSR[ 15 ][ 320 ],
   alphaCSR[ 15 ][ 321 ],
   alphaCSR[ 15 ][ 322 ],
   alphaCSR[ 15 ][ 323 ],
   alphaCSR[ 15 ][ 324 ],
   alphaCSR[ 15 ][ 325 ],
   alphaCSR[ 15 ][ 326 ],
   alphaCSR[ 15 ][ 327 ],
   alphaCSR[ 15 ][ 328 ],
   alphaCSR[ 15 ][ 329 ],
   alphaCSR[ 15 ][ 330 ],
   alphaCSR[ 15 ][ 331 ],
   alphaCSR[ 15 ][ 332 ],
   alphaCSR[ 15 ][ 333 ],
   alphaCSR[ 15 ][ 334 ],
   alphaCSR[ 15 ][ 335 ],
   alphaCSR[ 15 ][ 336 ],
   alphaCSR[ 15 ][ 337 ],
   alphaCSR[ 15 ][ 338 ],
   alphaCSR[ 15 ][ 339 ],
   alphaCSR[ 15 ][ 340 ],
   alphaCSR[ 15 ][ 341 ],
   alphaCSR[ 15 ][ 342 ],
   alphaCSR[ 15 ][ 343 ],
   alphaCSR[ 15 ][ 344 ],
   alphaCSR[ 15 ][ 345 ],
   alphaCSR[ 15 ][ 346 ],
   alphaCSR[ 15 ][ 347 ],
   alphaCSR[ 15 ][ 348 ],
   alphaCSR[ 15 ][ 349 ],
   alphaCSR[ 15 ][ 350 ],
   alphaCSR[ 15 ][ 351 ],
   alphaCSR[ 15 ][ 352 ],
   alphaCSR[ 15 ][ 353 ],
   alphaCSR[ 15 ][ 354 ],
   alphaCSR[ 15 ][ 355 ],
   alphaCSR[ 15 ][ 356 ],
   alphaCSR[ 15 ][ 357 ],
   alphaCSR[ 15 ][ 358 ],
   alphaCSR[ 15 ][ 359 ],
   alphaCSR[ 15 ][ 360 ],
   alphaCSR[ 15 ][ 361 ],
   alphaCSR[ 15 ][ 362 ],
   alphaCSR[ 15 ][ 363 ],
   alphaCSR[ 15 ][ 364 ],
   alphaCSR[ 15 ][ 365 ],
   alphaCSR[ 15 ][ 366 ],
   alphaCSR[ 15 ][ 367 ],
   alphaCSR[ 15 ][ 368 ],
   alphaCSR[ 15 ][ 369 ],
   alphaCSR[ 15 ][ 370 ],
   alphaCSR[ 15 ][ 371 ],
   alphaCSR[ 15 ][ 372 ],
   alphaCSR[ 15 ][ 373 ],
   alphaCSR[ 15 ][ 374 ],
   alphaCSR[ 15 ][ 375 ],
   alphaCSR[ 15 ][ 376 ],
   alphaCSR[ 15 ][ 377 ],
   alphaCSR[ 15 ][ 378 ],
   alphaCSR[ 15 ][ 379 ],
   alphaCSR[ 15 ][ 380 ],
   alphaCSR[ 15 ][ 381 ],
   alphaCSR[ 15 ][ 382 ],
   alphaCSR[ 15 ][ 383 ],
   alphaCSR[ 16 ][ 0 ],
   alphaCSR[ 16 ][ 1 ],
   alphaCSR[ 16 ][ 2 ],
   alphaCSR[ 16 ][ 3 ],
   alphaCSR[ 16 ][ 4 ],
   alphaCSR[ 16 ][ 5 ],
   alphaCSR[ 16 ][ 6 ],
   alphaCSR[ 16 ][ 7 ],
   alphaCSR[ 16 ][ 8 ],
   alphaCSR[ 16 ][ 9 ],
   alphaCSR[ 16 ][ 10 ],
   alphaCSR[ 16 ][ 11 ],
   alphaCSR[ 16 ][ 12 ],
   alphaCSR[ 16 ][ 13 ],
   alphaCSR[ 16 ][ 14 ],
   alphaCSR[ 16 ][ 15 ],
   alphaCSR[ 16 ][ 16 ],
   alphaCSR[ 16 ][ 17 ],
   alphaCSR[ 16 ][ 18 ],
   alphaCSR[ 16 ][ 19 ],
   alphaCSR[ 16 ][ 20 ],
   alphaCSR[ 16 ][ 21 ],
   alphaCSR[ 16 ][ 22 ],
   alphaCSR[ 16 ][ 23 ],
   alphaCSR[ 16 ][ 24 ],
   alphaCSR[ 16 ][ 25 ],
   alphaCSR[ 16 ][ 26 ],
   alphaCSR[ 16 ][ 27 ],
   alphaCSR[ 16 ][ 28 ],
   alphaCSR[ 16 ][ 29 ],
   alphaCSR[ 16 ][ 30 ],
   alphaCSR[ 16 ][ 31 ],
   alphaCSR[ 16 ][ 32 ],
   alphaCSR[ 16 ][ 33 ],
   alphaCSR[ 16 ][ 34 ],
   alphaCSR[ 16 ][ 35 ],
   alphaCSR[ 16 ][ 36 ],
   alphaCSR[ 16 ][ 37 ],
   alphaCSR[ 16 ][ 38 ],
   alphaCSR[ 16 ][ 39 ],
   alphaCSR[ 16 ][ 40 ],
   alphaCSR[ 16 ][ 41 ],
   alphaCSR[ 16 ][ 42 ],
   alphaCSR[ 16 ][ 43 ],
   alphaCSR[ 16 ][ 44 ],
   alphaCSR[ 16 ][ 45 ],
   alphaCSR[ 16 ][ 46 ],
   alphaCSR[ 16 ][ 47 ],
   alphaCSR[ 16 ][ 48 ],
   alphaCSR[ 16 ][ 49 ],
   alphaCSR[ 16 ][ 50 ],
   alphaCSR[ 16 ][ 51 ],
   alphaCSR[ 16 ][ 52 ],
   alphaCSR[ 16 ][ 53 ],
   alphaCSR[ 16 ][ 54 ],
   alphaCSR[ 16 ][ 55 ],
   alphaCSR[ 16 ][ 56 ],
   alphaCSR[ 16 ][ 57 ],
   alphaCSR[ 16 ][ 58 ],
   alphaCSR[ 16 ][ 59 ],
   alphaCSR[ 16 ][ 60 ],
   alphaCSR[ 16 ][ 61 ],
   alphaCSR[ 16 ][ 62 ],
   alphaCSR[ 16 ][ 63 ],
   alphaCSR[ 16 ][ 64 ],
   alphaCSR[ 16 ][ 65 ],
   alphaCSR[ 16 ][ 66 ],
   alphaCSR[ 16 ][ 67 ],
   alphaCSR[ 16 ][ 68 ],
   alphaCSR[ 16 ][ 69 ],
   alphaCSR[ 16 ][ 70 ],
   alphaCSR[ 16 ][ 71 ],
   alphaCSR[ 16 ][ 72 ],
   alphaCSR[ 16 ][ 73 ],
   alphaCSR[ 16 ][ 74 ],
   alphaCSR[ 16 ][ 75 ],
   alphaCSR[ 16 ][ 76 ],
   alphaCSR[ 16 ][ 77 ],
   alphaCSR[ 16 ][ 78 ],
   alphaCSR[ 16 ][ 79 ],
   alphaCSR[ 16 ][ 80 ],
   alphaCSR[ 16 ][ 81 ],
   alphaCSR[ 16 ][ 82 ],
   alphaCSR[ 16 ][ 83 ],
   alphaCSR[ 16 ][ 84 ],
   alphaCSR[ 16 ][ 85 ],
   alphaCSR[ 16 ][ 86 ],
   alphaCSR[ 16 ][ 87 ],
   alphaCSR[ 16 ][ 88 ],
   alphaCSR[ 16 ][ 89 ],
   alphaCSR[ 16 ][ 90 ],
   alphaCSR[ 16 ][ 91 ],
   alphaCSR[ 16 ][ 92 ],
   alphaCSR[ 16 ][ 93 ],
   alphaCSR[ 16 ][ 94 ],
   alphaCSR[ 16 ][ 95 ],
   alphaCSR[ 16 ][ 96 ],
   alphaCSR[ 16 ][ 97 ],
   alphaCSR[ 16 ][ 98 ],
   alphaCSR[ 16 ][ 99 ],
   alphaCSR[ 16 ][ 100 ],
   alphaCSR[ 16 ][ 101 ],
   alphaCSR[ 16 ][ 102 ],
   alphaCSR[ 16 ][ 103 ],
   alphaCSR[ 16 ][ 104 ],
   alphaCSR[ 16 ][ 105 ],
   alphaCSR[ 16 ][ 106 ],
   alphaCSR[ 16 ][ 107 ],
   alphaCSR[ 16 ][ 108 ],
   alphaCSR[ 16 ][ 109 ],
   alphaCSR[ 16 ][ 110 ],
   alphaCSR[ 16 ][ 111 ],
   alphaCSR[ 16 ][ 112 ],
   alphaCSR[ 16 ][ 113 ],
   alphaCSR[ 16 ][ 114 ],
   alphaCSR[ 16 ][ 115 ],
   alphaCSR[ 16 ][ 116 ],
   alphaCSR[ 16 ][ 117 ],
   alphaCSR[ 16 ][ 118 ],
   alphaCSR[ 16 ][ 119 ],
   alphaCSR[ 16 ][ 120 ],
   alphaCSR[ 16 ][ 121 ],
   alphaCSR[ 16 ][ 122 ],
   alphaCSR[ 16 ][ 123 ],
   alphaCSR[ 16 ][ 124 ],
   alphaCSR[ 16 ][ 125 ],
   alphaCSR[ 16 ][ 126 ],
   alphaCSR[ 16 ][ 127 ],
   alphaCSR[ 16 ][ 128 ],
   alphaCSR[ 16 ][ 129 ],
   alphaCSR[ 16 ][ 130 ],
   alphaCSR[ 16 ][ 131 ],
   alphaCSR[ 16 ][ 132 ],
   alphaCSR[ 16 ][ 133 ],
   alphaCSR[ 16 ][ 134 ],
   alphaCSR[ 16 ][ 135 ],
   alphaCSR[ 16 ][ 136 ],
   alphaCSR[ 16 ][ 137 ],
   alphaCSR[ 16 ][ 138 ],
   alphaCSR[ 16 ][ 139 ],
   alphaCSR[ 16 ][ 140 ],
   alphaCSR[ 16 ][ 141 ],
   alphaCSR[ 16 ][ 142 ],
   alphaCSR[ 16 ][ 143 ],
   alphaCSR[ 16 ][ 144 ],
   alphaCSR[ 16 ][ 145 ],
   alphaCSR[ 16 ][ 146 ],
   alphaCSR[ 16 ][ 147 ],
   alphaCSR[ 16 ][ 148 ],
   alphaCSR[ 16 ][ 149 ],
   alphaCSR[ 16 ][ 150 ],
   alphaCSR[ 16 ][ 151 ],
   alphaCSR[ 16 ][ 152 ],
   alphaCSR[ 16 ][ 153 ],
   alphaCSR[ 16 ][ 154 ],
   alphaCSR[ 16 ][ 155 ],
   alphaCSR[ 16 ][ 156 ],
   alphaCSR[ 16 ][ 157 ],
   alphaCSR[ 16 ][ 158 ],
   alphaCSR[ 16 ][ 159 ],
   alphaCSR[ 16 ][ 160 ],
   alphaCSR[ 16 ][ 161 ],
   alphaCSR[ 16 ][ 162 ],
   alphaCSR[ 16 ][ 163 ],
   alphaCSR[ 16 ][ 164 ],
   alphaCSR[ 16 ][ 165 ],
   alphaCSR[ 16 ][ 166 ],
   alphaCSR[ 16 ][ 167 ],
   alphaCSR[ 16 ][ 168 ],
   alphaCSR[ 16 ][ 169 ],
   alphaCSR[ 16 ][ 170 ],
   alphaCSR[ 16 ][ 171 ],
   alphaCSR[ 16 ][ 172 ],
   alphaCSR[ 16 ][ 173 ],
   alphaCSR[ 16 ][ 174 ],
   alphaCSR[ 16 ][ 175 ],
   alphaCSR[ 16 ][ 176 ],
   alphaCSR[ 16 ][ 177 ],
   alphaCSR[ 16 ][ 178 ],
   alphaCSR[ 16 ][ 179 ],
   alphaCSR[ 16 ][ 180 ],
   alphaCSR[ 16 ][ 181 ],
   alphaCSR[ 16 ][ 182 ],
   alphaCSR[ 16 ][ 183 ],
   alphaCSR[ 16 ][ 184 ],
   alphaCSR[ 16 ][ 185 ],
   alphaCSR[ 16 ][ 186 ],
   alphaCSR[ 16 ][ 187 ],
   alphaCSR[ 16 ][ 188 ],
   alphaCSR[ 16 ][ 189 ],
   alphaCSR[ 16 ][ 190 ],
   alphaCSR[ 16 ][ 191 ],
   alphaCSR[ 16 ][ 192 ],
   alphaCSR[ 16 ][ 193 ],
   alphaCSR[ 16 ][ 194 ],
   alphaCSR[ 16 ][ 195 ],
   alphaCSR[ 16 ][ 196 ],
   alphaCSR[ 16 ][ 197 ],
   alphaCSR[ 16 ][ 198 ],
   alphaCSR[ 16 ][ 199 ],
   alphaCSR[ 16 ][ 200 ],
   alphaCSR[ 16 ][ 201 ],
   alphaCSR[ 16 ][ 202 ],
   alphaCSR[ 16 ][ 203 ],
   alphaCSR[ 16 ][ 204 ],
   alphaCSR[ 16 ][ 205 ],
   alphaCSR[ 16 ][ 206 ],
   alphaCSR[ 16 ][ 207 ],
   alphaCSR[ 16 ][ 208 ],
   alphaCSR[ 16 ][ 209 ],
   alphaCSR[ 16 ][ 210 ],
   alphaCSR[ 16 ][ 211 ],
   alphaCSR[ 16 ][ 212 ],
   alphaCSR[ 16 ][ 213 ],
   alphaCSR[ 16 ][ 214 ],
   alphaCSR[ 16 ][ 215 ],
   alphaCSR[ 16 ][ 216 ],
   alphaCSR[ 16 ][ 217 ],
   alphaCSR[ 16 ][ 218 ],
   alphaCSR[ 16 ][ 219 ],
   alphaCSR[ 16 ][ 220 ],
   alphaCSR[ 16 ][ 221 ],
   alphaCSR[ 16 ][ 222 ],
   alphaCSR[ 16 ][ 223 ],
   alphaCSR[ 16 ][ 224 ],
   alphaCSR[ 16 ][ 225 ],
   alphaCSR[ 16 ][ 226 ],
   alphaCSR[ 16 ][ 227 ],
   alphaCSR[ 16 ][ 228 ],
   alphaCSR[ 16 ][ 229 ],
   alphaCSR[ 16 ][ 230 ],
   alphaCSR[ 16 ][ 231 ],
   alphaCSR[ 16 ][ 232 ],
   alphaCSR[ 16 ][ 233 ],
   alphaCSR[ 16 ][ 234 ],
   alphaCSR[ 16 ][ 235 ],
   alphaCSR[ 16 ][ 236 ],
   alphaCSR[ 16 ][ 237 ],
   alphaCSR[ 16 ][ 238 ],
   alphaCSR[ 16 ][ 239 ],
   alphaCSR[ 16 ][ 240 ],
   alphaCSR[ 16 ][ 241 ],
   alphaCSR[ 16 ][ 242 ],
   alphaCSR[ 16 ][ 243 ],
   alphaCSR[ 16 ][ 244 ],
   alphaCSR[ 16 ][ 245 ],
   alphaCSR[ 16 ][ 246 ],
   alphaCSR[ 16 ][ 247 ],
   alphaCSR[ 16 ][ 248 ],
   alphaCSR[ 16 ][ 249 ],
   alphaCSR[ 16 ][ 250 ],
   alphaCSR[ 16 ][ 251 ],
   alphaCSR[ 16 ][ 252 ],
   alphaCSR[ 16 ][ 253 ],
   alphaCSR[ 16 ][ 254 ],
   alphaCSR[ 16 ][ 255 ],
   alphaCSR[ 16 ][ 256 ],
   alphaCSR[ 16 ][ 257 ],
   alphaCSR[ 16 ][ 258 ],
   alphaCSR[ 16 ][ 259 ],
   alphaCSR[ 16 ][ 260 ],
   alphaCSR[ 16 ][ 261 ],
   alphaCSR[ 16 ][ 262 ],
   alphaCSR[ 16 ][ 263 ],
   alphaCSR[ 16 ][ 264 ],
   alphaCSR[ 16 ][ 265 ],
   alphaCSR[ 16 ][ 266 ],
   alphaCSR[ 16 ][ 267 ],
   alphaCSR[ 16 ][ 268 ],
   alphaCSR[ 16 ][ 269 ],
   alphaCSR[ 16 ][ 270 ],
   alphaCSR[ 16 ][ 271 ],
   alphaCSR[ 16 ][ 272 ],
   alphaCSR[ 16 ][ 273 ],
   alphaCSR[ 16 ][ 274 ],
   alphaCSR[ 16 ][ 275 ],
   alphaCSR[ 16 ][ 276 ],
   alphaCSR[ 16 ][ 277 ],
   alphaCSR[ 16 ][ 278 ],
   alphaCSR[ 16 ][ 279 ],
   alphaCSR[ 16 ][ 280 ],
   alphaCSR[ 16 ][ 281 ],
   alphaCSR[ 16 ][ 282 ],
   alphaCSR[ 16 ][ 283 ],
   alphaCSR[ 16 ][ 284 ],
   alphaCSR[ 16 ][ 285 ],
   alphaCSR[ 16 ][ 286 ],
   alphaCSR[ 16 ][ 287 ],
   alphaCSR[ 16 ][ 288 ],
   alphaCSR[ 16 ][ 289 ],
   alphaCSR[ 16 ][ 290 ],
   alphaCSR[ 16 ][ 291 ],
   alphaCSR[ 16 ][ 292 ],
   alphaCSR[ 16 ][ 293 ],
   alphaCSR[ 16 ][ 294 ],
   alphaCSR[ 16 ][ 295 ],
   alphaCSR[ 16 ][ 296 ],
   alphaCSR[ 16 ][ 297 ],
   alphaCSR[ 16 ][ 298 ],
   alphaCSR[ 16 ][ 299 ],
   alphaCSR[ 16 ][ 300 ],
   alphaCSR[ 16 ][ 301 ],
   alphaCSR[ 16 ][ 302 ],
   alphaCSR[ 16 ][ 303 ],
   alphaCSR[ 16 ][ 304 ],
   alphaCSR[ 16 ][ 305 ],
   alphaCSR[ 16 ][ 306 ],
   alphaCSR[ 16 ][ 307 ],
   alphaCSR[ 16 ][ 308 ],
   alphaCSR[ 16 ][ 309 ],
   alphaCSR[ 16 ][ 310 ],
   alphaCSR[ 16 ][ 311 ],
   alphaCSR[ 16 ][ 312 ],
   alphaCSR[ 16 ][ 313 ],
   alphaCSR[ 16 ][ 314 ],
   alphaCSR[ 16 ][ 315 ],
   alphaCSR[ 16 ][ 316 ],
   alphaCSR[ 16 ][ 317 ],
   alphaCSR[ 16 ][ 318 ],
   alphaCSR[ 16 ][ 319 ],
   alphaCSR[ 16 ][ 320 ],
   alphaCSR[ 16 ][ 321 ],
   alphaCSR[ 16 ][ 322 ],
   alphaCSR[ 16 ][ 323 ],
   alphaCSR[ 16 ][ 324 ],
   alphaCSR[ 16 ][ 325 ],
   alphaCSR[ 16 ][ 326 ],
   alphaCSR[ 16 ][ 327 ],
   alphaCSR[ 16 ][ 328 ],
   alphaCSR[ 16 ][ 329 ],
   alphaCSR[ 16 ][ 330 ],
   alphaCSR[ 16 ][ 331 ],
   alphaCSR[ 16 ][ 332 ],
   alphaCSR[ 16 ][ 333 ],
   alphaCSR[ 16 ][ 334 ],
   alphaCSR[ 16 ][ 335 ],
   alphaCSR[ 16 ][ 336 ],
   alphaCSR[ 16 ][ 337 ],
   alphaCSR[ 16 ][ 338 ],
   alphaCSR[ 16 ][ 339 ],
   alphaCSR[ 16 ][ 340 ],
   alphaCSR[ 16 ][ 341 ],
   alphaCSR[ 16 ][ 342 ],
   alphaCSR[ 16 ][ 343 ],
   alphaCSR[ 16 ][ 344 ],
   alphaCSR[ 16 ][ 345 ],
   alphaCSR[ 16 ][ 346 ],
   alphaCSR[ 16 ][ 347 ],
   alphaCSR[ 16 ][ 348 ],
   alphaCSR[ 16 ][ 349 ],
   alphaCSR[ 16 ][ 350 ],
   alphaCSR[ 16 ][ 351 ],
   alphaCSR[ 16 ][ 352 ],
   alphaCSR[ 16 ][ 353 ],
   alphaCSR[ 16 ][ 354 ],
   alphaCSR[ 16 ][ 355 ],
   alphaCSR[ 16 ][ 356 ],
   alphaCSR[ 16 ][ 357 ],
   alphaCSR[ 16 ][ 358 ],
   alphaCSR[ 16 ][ 359 ],
   alphaCSR[ 16 ][ 360 ],
   alphaCSR[ 16 ][ 361 ],
   alphaCSR[ 16 ][ 362 ],
   alphaCSR[ 16 ][ 363 ],
   alphaCSR[ 16 ][ 364 ],
   alphaCSR[ 16 ][ 365 ],
   alphaCSR[ 16 ][ 366 ],
   alphaCSR[ 16 ][ 367 ],
   alphaCSR[ 16 ][ 368 ],
   alphaCSR[ 16 ][ 369 ],
   alphaCSR[ 16 ][ 370 ],
   alphaCSR[ 16 ][ 371 ],
   alphaCSR[ 16 ][ 372 ],
   alphaCSR[ 16 ][ 373 ],
   alphaCSR[ 16 ][ 374 ],
   alphaCSR[ 16 ][ 375 ],
   alphaCSR[ 16 ][ 376 ],
   alphaCSR[ 16 ][ 377 ],
   alphaCSR[ 16 ][ 378 ],
   alphaCSR[ 16 ][ 379 ],
   alphaCSR[ 16 ][ 380 ],
   alphaCSR[ 16 ][ 381 ],
   alphaCSR[ 16 ][ 382 ],
   alphaCSR[ 16 ][ 383 ],
   alphaCSR[ 17 ][ 0 ],
   alphaCSR[ 17 ][ 1 ],
   alphaCSR[ 17 ][ 2 ],
   alphaCSR[ 17 ][ 3 ],
   alphaCSR[ 17 ][ 4 ],
   alphaCSR[ 17 ][ 5 ],
   alphaCSR[ 17 ][ 6 ],
   alphaCSR[ 17 ][ 7 ],
   alphaCSR[ 17 ][ 8 ],
   alphaCSR[ 17 ][ 9 ],
   alphaCSR[ 17 ][ 10 ],
   alphaCSR[ 17 ][ 11 ],
   alphaCSR[ 17 ][ 12 ],
   alphaCSR[ 17 ][ 13 ],
   alphaCSR[ 17 ][ 14 ],
   alphaCSR[ 17 ][ 15 ],
   alphaCSR[ 17 ][ 16 ],
   alphaCSR[ 17 ][ 17 ],
   alphaCSR[ 17 ][ 18 ],
   alphaCSR[ 17 ][ 19 ],
   alphaCSR[ 17 ][ 20 ],
   alphaCSR[ 17 ][ 21 ],
   alphaCSR[ 17 ][ 22 ],
   alphaCSR[ 17 ][ 23 ],
   alphaCSR[ 17 ][ 24 ],
   alphaCSR[ 17 ][ 25 ],
   alphaCSR[ 17 ][ 26 ],
   alphaCSR[ 17 ][ 27 ],
   alphaCSR[ 17 ][ 28 ],
   alphaCSR[ 17 ][ 29 ],
   alphaCSR[ 17 ][ 30 ],
   alphaCSR[ 17 ][ 31 ],
   alphaCSR[ 17 ][ 32 ],
   alphaCSR[ 17 ][ 33 ],
   alphaCSR[ 17 ][ 34 ],
   alphaCSR[ 17 ][ 35 ],
   alphaCSR[ 17 ][ 36 ],
   alphaCSR[ 17 ][ 37 ],
   alphaCSR[ 17 ][ 38 ],
   alphaCSR[ 17 ][ 39 ],
   alphaCSR[ 17 ][ 40 ],
   alphaCSR[ 17 ][ 41 ],
   alphaCSR[ 17 ][ 42 ],
   alphaCSR[ 17 ][ 43 ],
   alphaCSR[ 17 ][ 44 ],
   alphaCSR[ 17 ][ 45 ],
   alphaCSR[ 17 ][ 46 ],
   alphaCSR[ 17 ][ 47 ],
   alphaCSR[ 17 ][ 48 ],
   alphaCSR[ 17 ][ 49 ],
   alphaCSR[ 17 ][ 50 ],
   alphaCSR[ 17 ][ 51 ],
   alphaCSR[ 17 ][ 52 ],
   alphaCSR[ 17 ][ 53 ],
   alphaCSR[ 17 ][ 54 ],
   alphaCSR[ 17 ][ 55 ],
   alphaCSR[ 17 ][ 56 ],
   alphaCSR[ 17 ][ 57 ],
   alphaCSR[ 17 ][ 58 ],
   alphaCSR[ 17 ][ 59 ],
   alphaCSR[ 17 ][ 60 ],
   alphaCSR[ 17 ][ 61 ],
   alphaCSR[ 17 ][ 62 ],
   alphaCSR[ 17 ][ 63 ],
   alphaCSR[ 17 ][ 64 ],
   alphaCSR[ 17 ][ 65 ],
   alphaCSR[ 17 ][ 66 ],
   alphaCSR[ 17 ][ 67 ],
   alphaCSR[ 17 ][ 68 ],
   alphaCSR[ 17 ][ 69 ],
   alphaCSR[ 17 ][ 70 ],
   alphaCSR[ 17 ][ 71 ],
   alphaCSR[ 17 ][ 72 ],
   alphaCSR[ 17 ][ 73 ],
   alphaCSR[ 17 ][ 74 ],
   alphaCSR[ 17 ][ 75 ],
   alphaCSR[ 17 ][ 76 ],
   alphaCSR[ 17 ][ 77 ],
   alphaCSR[ 17 ][ 78 ],
   alphaCSR[ 17 ][ 79 ],
   alphaCSR[ 17 ][ 80 ],
   alphaCSR[ 17 ][ 81 ],
   alphaCSR[ 17 ][ 82 ],
   alphaCSR[ 17 ][ 83 ],
   alphaCSR[ 17 ][ 84 ],
   alphaCSR[ 17 ][ 85 ],
   alphaCSR[ 17 ][ 86 ],
   alphaCSR[ 17 ][ 87 ],
   alphaCSR[ 17 ][ 88 ],
   alphaCSR[ 17 ][ 89 ],
   alphaCSR[ 17 ][ 90 ],
   alphaCSR[ 17 ][ 91 ],
   alphaCSR[ 17 ][ 92 ],
   alphaCSR[ 17 ][ 93 ],
   alphaCSR[ 17 ][ 94 ],
   alphaCSR[ 17 ][ 95 ],
   alphaCSR[ 17 ][ 96 ],
   alphaCSR[ 17 ][ 97 ],
   alphaCSR[ 17 ][ 98 ],
   alphaCSR[ 17 ][ 99 ],
   alphaCSR[ 17 ][ 100 ],
   alphaCSR[ 17 ][ 101 ],
   alphaCSR[ 17 ][ 102 ],
   alphaCSR[ 17 ][ 103 ],
   alphaCSR[ 17 ][ 104 ],
   alphaCSR[ 17 ][ 105 ],
   alphaCSR[ 17 ][ 106 ],
   alphaCSR[ 17 ][ 107 ],
   alphaCSR[ 17 ][ 108 ],
   alphaCSR[ 17 ][ 109 ],
   alphaCSR[ 17 ][ 110 ],
   alphaCSR[ 17 ][ 111 ],
   alphaCSR[ 17 ][ 112 ],
   alphaCSR[ 17 ][ 113 ],
   alphaCSR[ 17 ][ 114 ],
   alphaCSR[ 17 ][ 115 ],
   alphaCSR[ 17 ][ 116 ],
   alphaCSR[ 17 ][ 117 ],
   alphaCSR[ 17 ][ 118 ],
   alphaCSR[ 17 ][ 119 ],
   alphaCSR[ 17 ][ 120 ],
   alphaCSR[ 17 ][ 121 ],
   alphaCSR[ 17 ][ 122 ],
   alphaCSR[ 17 ][ 123 ],
   alphaCSR[ 17 ][ 124 ],
   alphaCSR[ 17 ][ 125 ],
   alphaCSR[ 17 ][ 126 ],
   alphaCSR[ 17 ][ 127 ],
   alphaCSR[ 17 ][ 128 ],
   alphaCSR[ 17 ][ 129 ],
   alphaCSR[ 17 ][ 130 ],
   alphaCSR[ 17 ][ 131 ],
   alphaCSR[ 17 ][ 132 ],
   alphaCSR[ 17 ][ 133 ],
   alphaCSR[ 17 ][ 134 ],
   alphaCSR[ 17 ][ 135 ],
   alphaCSR[ 17 ][ 136 ],
   alphaCSR[ 17 ][ 137 ],
   alphaCSR[ 17 ][ 138 ],
   alphaCSR[ 17 ][ 139 ],
   alphaCSR[ 17 ][ 140 ],
   alphaCSR[ 17 ][ 141 ],
   alphaCSR[ 17 ][ 142 ],
   alphaCSR[ 17 ][ 143 ],
   alphaCSR[ 17 ][ 144 ],
   alphaCSR[ 17 ][ 145 ],
   alphaCSR[ 17 ][ 146 ],
   alphaCSR[ 17 ][ 147 ],
   alphaCSR[ 17 ][ 148 ],
   alphaCSR[ 17 ][ 149 ],
   alphaCSR[ 17 ][ 150 ],
   alphaCSR[ 17 ][ 151 ],
   alphaCSR[ 17 ][ 152 ],
   alphaCSR[ 17 ][ 153 ],
   alphaCSR[ 17 ][ 154 ],
   alphaCSR[ 17 ][ 155 ],
   alphaCSR[ 17 ][ 156 ],
   alphaCSR[ 17 ][ 157 ],
   alphaCSR[ 17 ][ 158 ],
   alphaCSR[ 17 ][ 159 ],
   alphaCSR[ 17 ][ 160 ],
   alphaCSR[ 17 ][ 161 ],
   alphaCSR[ 17 ][ 162 ],
   alphaCSR[ 17 ][ 163 ],
   alphaCSR[ 17 ][ 164 ],
   alphaCSR[ 17 ][ 165 ],
   alphaCSR[ 17 ][ 166 ],
   alphaCSR[ 17 ][ 167 ],
   alphaCSR[ 17 ][ 168 ],
   alphaCSR[ 17 ][ 169 ],
   alphaCSR[ 17 ][ 170 ],
   alphaCSR[ 17 ][ 171 ],
   alphaCSR[ 17 ][ 172 ],
   alphaCSR[ 17 ][ 173 ],
   alphaCSR[ 17 ][ 174 ],
   alphaCSR[ 17 ][ 175 ],
   alphaCSR[ 17 ][ 176 ],
   alphaCSR[ 17 ][ 177 ],
   alphaCSR[ 17 ][ 178 ],
   alphaCSR[ 17 ][ 179 ],
   alphaCSR[ 17 ][ 180 ],
   alphaCSR[ 17 ][ 181 ],
   alphaCSR[ 17 ][ 182 ],
   alphaCSR[ 17 ][ 183 ],
   alphaCSR[ 17 ][ 184 ],
   alphaCSR[ 17 ][ 185 ],
   alphaCSR[ 17 ][ 186 ],
   alphaCSR[ 17 ][ 187 ],
   alphaCSR[ 17 ][ 188 ],
   alphaCSR[ 17 ][ 189 ],
   alphaCSR[ 17 ][ 190 ],
   alphaCSR[ 17 ][ 191 ],
   alphaCSR[ 17 ][ 192 ],
   alphaCSR[ 17 ][ 193 ],
   alphaCSR[ 17 ][ 194 ],
   alphaCSR[ 17 ][ 195 ],
   alphaCSR[ 17 ][ 196 ],
   alphaCSR[ 17 ][ 197 ],
   alphaCSR[ 17 ][ 198 ],
   alphaCSR[ 17 ][ 199 ],
   alphaCSR[ 17 ][ 200 ],
   alphaCSR[ 17 ][ 201 ],
   alphaCSR[ 17 ][ 202 ],
   alphaCSR[ 17 ][ 203 ],
   alphaCSR[ 17 ][ 204 ],
   alphaCSR[ 17 ][ 205 ],
   alphaCSR[ 17 ][ 206 ],
   alphaCSR[ 17 ][ 207 ],
   alphaCSR[ 17 ][ 208 ],
   alphaCSR[ 17 ][ 209 ],
   alphaCSR[ 17 ][ 210 ],
   alphaCSR[ 17 ][ 211 ],
   alphaCSR[ 17 ][ 212 ],
   alphaCSR[ 17 ][ 213 ],
   alphaCSR[ 17 ][ 214 ],
   alphaCSR[ 17 ][ 215 ],
   alphaCSR[ 17 ][ 216 ],
   alphaCSR[ 17 ][ 217 ],
   alphaCSR[ 17 ][ 218 ],
   alphaCSR[ 17 ][ 219 ],
   alphaCSR[ 17 ][ 220 ],
   alphaCSR[ 17 ][ 221 ],
   alphaCSR[ 17 ][ 222 ],
   alphaCSR[ 17 ][ 223 ],
   alphaCSR[ 17 ][ 224 ],
   alphaCSR[ 17 ][ 225 ],
   alphaCSR[ 17 ][ 226 ],
   alphaCSR[ 17 ][ 227 ],
   alphaCSR[ 17 ][ 228 ],
   alphaCSR[ 17 ][ 229 ],
   alphaCSR[ 17 ][ 230 ],
   alphaCSR[ 17 ][ 231 ],
   alphaCSR[ 17 ][ 232 ],
   alphaCSR[ 17 ][ 233 ],
   alphaCSR[ 17 ][ 234 ],
   alphaCSR[ 17 ][ 235 ],
   alphaCSR[ 17 ][ 236 ],
   alphaCSR[ 17 ][ 237 ],
   alphaCSR[ 17 ][ 238 ],
   alphaCSR[ 17 ][ 239 ],
   alphaCSR[ 17 ][ 240 ],
   alphaCSR[ 17 ][ 241 ],
   alphaCSR[ 17 ][ 242 ],
   alphaCSR[ 17 ][ 243 ],
   alphaCSR[ 17 ][ 244 ],
   alphaCSR[ 17 ][ 245 ],
   alphaCSR[ 17 ][ 246 ],
   alphaCSR[ 17 ][ 247 ],
   alphaCSR[ 17 ][ 248 ],
   alphaCSR[ 17 ][ 249 ],
   alphaCSR[ 17 ][ 250 ],
   alphaCSR[ 17 ][ 251 ],
   alphaCSR[ 17 ][ 252 ],
   alphaCSR[ 17 ][ 253 ],
   alphaCSR[ 17 ][ 254 ],
   alphaCSR[ 17 ][ 255 ],
   alphaCSR[ 17 ][ 256 ],
   alphaCSR[ 17 ][ 257 ],
   alphaCSR[ 17 ][ 258 ],
   alphaCSR[ 17 ][ 259 ],
   alphaCSR[ 17 ][ 260 ],
   alphaCSR[ 17 ][ 261 ],
   alphaCSR[ 17 ][ 262 ],
   alphaCSR[ 17 ][ 263 ],
   alphaCSR[ 17 ][ 264 ],
   alphaCSR[ 17 ][ 265 ],
   alphaCSR[ 17 ][ 266 ],
   alphaCSR[ 17 ][ 267 ],
   alphaCSR[ 17 ][ 268 ],
   alphaCSR[ 17 ][ 269 ],
   alphaCSR[ 17 ][ 270 ],
   alphaCSR[ 17 ][ 271 ],
   alphaCSR[ 17 ][ 272 ],
   alphaCSR[ 17 ][ 273 ],
   alphaCSR[ 17 ][ 274 ],
   alphaCSR[ 17 ][ 275 ],
   alphaCSR[ 17 ][ 276 ],
   alphaCSR[ 17 ][ 277 ],
   alphaCSR[ 17 ][ 278 ],
   alphaCSR[ 17 ][ 279 ],
   alphaCSR[ 17 ][ 280 ],
   alphaCSR[ 17 ][ 281 ],
   alphaCSR[ 17 ][ 282 ],
   alphaCSR[ 17 ][ 283 ],
   alphaCSR[ 17 ][ 284 ],
   alphaCSR[ 17 ][ 285 ],
   alphaCSR[ 17 ][ 286 ],
   alphaCSR[ 17 ][ 287 ],
   alphaCSR[ 17 ][ 288 ],
   alphaCSR[ 17 ][ 289 ],
   alphaCSR[ 17 ][ 290 ],
   alphaCSR[ 17 ][ 291 ],
   alphaCSR[ 17 ][ 292 ],
   alphaCSR[ 17 ][ 293 ],
   alphaCSR[ 17 ][ 294 ],
   alphaCSR[ 17 ][ 295 ],
   alphaCSR[ 17 ][ 296 ],
   alphaCSR[ 17 ][ 297 ],
   alphaCSR[ 17 ][ 298 ],
   alphaCSR[ 17 ][ 299 ],
   alphaCSR[ 17 ][ 300 ],
   alphaCSR[ 17 ][ 301 ],
   alphaCSR[ 17 ][ 302 ],
   alphaCSR[ 17 ][ 303 ],
   alphaCSR[ 17 ][ 304 ],
   alphaCSR[ 17 ][ 305 ],
   alphaCSR[ 17 ][ 306 ],
   alphaCSR[ 17 ][ 307 ],
   alphaCSR[ 17 ][ 308 ],
   alphaCSR[ 17 ][ 309 ],
   alphaCSR[ 17 ][ 310 ],
   alphaCSR[ 17 ][ 311 ],
   alphaCSR[ 17 ][ 312 ],
   alphaCSR[ 17 ][ 313 ],
   alphaCSR[ 17 ][ 314 ],
   alphaCSR[ 17 ][ 315 ],
   alphaCSR[ 17 ][ 316 ],
   alphaCSR[ 17 ][ 317 ],
   alphaCSR[ 17 ][ 318 ],
   alphaCSR[ 17 ][ 319 ],
   alphaCSR[ 17 ][ 320 ],
   alphaCSR[ 17 ][ 321 ],
   alphaCSR[ 17 ][ 322 ],
   alphaCSR[ 17 ][ 323 ],
   alphaCSR[ 17 ][ 324 ],
   alphaCSR[ 17 ][ 325 ],
   alphaCSR[ 17 ][ 326 ],
   alphaCSR[ 17 ][ 327 ],
   alphaCSR[ 17 ][ 328 ],
   alphaCSR[ 17 ][ 329 ],
   alphaCSR[ 17 ][ 330 ],
   alphaCSR[ 17 ][ 331 ],
   alphaCSR[ 17 ][ 332 ],
   alphaCSR[ 17 ][ 333 ],
   alphaCSR[ 17 ][ 334 ],
   alphaCSR[ 17 ][ 335 ],
   alphaCSR[ 17 ][ 336 ],
   alphaCSR[ 17 ][ 337 ],
   alphaCSR[ 17 ][ 338 ],
   alphaCSR[ 17 ][ 339 ],
   alphaCSR[ 17 ][ 340 ],
   alphaCSR[ 17 ][ 341 ],
   alphaCSR[ 17 ][ 342 ],
   alphaCSR[ 17 ][ 343 ],
   alphaCSR[ 17 ][ 344 ],
   alphaCSR[ 17 ][ 345 ],
   alphaCSR[ 17 ][ 346 ],
   alphaCSR[ 17 ][ 347 ],
   alphaCSR[ 17 ][ 348 ],
   alphaCSR[ 17 ][ 349 ],
   alphaCSR[ 17 ][ 350 ],
   alphaCSR[ 17 ][ 351 ],
   alphaCSR[ 17 ][ 352 ],
   alphaCSR[ 17 ][ 353 ],
   alphaCSR[ 17 ][ 354 ],
   alphaCSR[ 17 ][ 355 ],
   alphaCSR[ 17 ][ 356 ],
   alphaCSR[ 17 ][ 357 ],
   alphaCSR[ 17 ][ 358 ],
   alphaCSR[ 17 ][ 359 ],
   alphaCSR[ 17 ][ 360 ],
   alphaCSR[ 17 ][ 361 ],
   alphaCSR[ 17 ][ 362 ],
   alphaCSR[ 17 ][ 363 ],
   alphaCSR[ 17 ][ 364 ],
   alphaCSR[ 17 ][ 365 ],
   alphaCSR[ 17 ][ 366 ],
   alphaCSR[ 17 ][ 367 ],
   alphaCSR[ 17 ][ 368 ],
   alphaCSR[ 17 ][ 369 ],
   alphaCSR[ 17 ][ 370 ],
   alphaCSR[ 17 ][ 371 ],
   alphaCSR[ 17 ][ 372 ],
   alphaCSR[ 17 ][ 373 ],
   alphaCSR[ 17 ][ 374 ],
   alphaCSR[ 17 ][ 375 ],
   alphaCSR[ 17 ][ 376 ],
   alphaCSR[ 17 ][ 377 ],
   alphaCSR[ 17 ][ 378 ],
   alphaCSR[ 17 ][ 379 ],
   alphaCSR[ 17 ][ 380 ],
   alphaCSR[ 17 ][ 381 ],
   alphaCSR[ 17 ][ 382 ],
   alphaCSR[ 17 ][ 383 ],
   alphaCSR[ 18 ][ 0 ],
   alphaCSR[ 18 ][ 1 ],
   alphaCSR[ 18 ][ 2 ],
   alphaCSR[ 18 ][ 3 ],
   alphaCSR[ 18 ][ 4 ],
   alphaCSR[ 18 ][ 5 ],
   alphaCSR[ 18 ][ 6 ],
   alphaCSR[ 18 ][ 7 ],
   alphaCSR[ 18 ][ 8 ],
   alphaCSR[ 18 ][ 9 ],
   alphaCSR[ 18 ][ 10 ],
   alphaCSR[ 18 ][ 11 ],
   alphaCSR[ 18 ][ 12 ],
   alphaCSR[ 18 ][ 13 ],
   alphaCSR[ 18 ][ 14 ],
   alphaCSR[ 18 ][ 15 ],
   alphaCSR[ 18 ][ 16 ],
   alphaCSR[ 18 ][ 17 ],
   alphaCSR[ 18 ][ 18 ],
   alphaCSR[ 18 ][ 19 ],
   alphaCSR[ 18 ][ 20 ],
   alphaCSR[ 18 ][ 21 ],
   alphaCSR[ 18 ][ 22 ],
   alphaCSR[ 18 ][ 23 ],
   alphaCSR[ 18 ][ 24 ],
   alphaCSR[ 18 ][ 25 ],
   alphaCSR[ 18 ][ 26 ],
   alphaCSR[ 18 ][ 27 ],
   alphaCSR[ 18 ][ 28 ],
   alphaCSR[ 18 ][ 29 ],
   alphaCSR[ 18 ][ 30 ],
   alphaCSR[ 18 ][ 31 ],
   alphaCSR[ 18 ][ 32 ],
   alphaCSR[ 18 ][ 33 ],
   alphaCSR[ 18 ][ 34 ],
   alphaCSR[ 18 ][ 35 ],
   alphaCSR[ 18 ][ 36 ],
   alphaCSR[ 18 ][ 37 ],
   alphaCSR[ 18 ][ 38 ],
   alphaCSR[ 18 ][ 39 ],
   alphaCSR[ 18 ][ 40 ],
   alphaCSR[ 18 ][ 41 ],
   alphaCSR[ 18 ][ 42 ],
   alphaCSR[ 18 ][ 43 ],
   alphaCSR[ 18 ][ 44 ],
   alphaCSR[ 18 ][ 45 ],
   alphaCSR[ 18 ][ 46 ],
   alphaCSR[ 18 ][ 47 ],
   alphaCSR[ 18 ][ 48 ],
   alphaCSR[ 18 ][ 49 ],
   alphaCSR[ 18 ][ 50 ],
   alphaCSR[ 18 ][ 51 ],
   alphaCSR[ 18 ][ 52 ],
   alphaCSR[ 18 ][ 53 ],
   alphaCSR[ 18 ][ 54 ],
   alphaCSR[ 18 ][ 55 ],
   alphaCSR[ 18 ][ 56 ],
   alphaCSR[ 18 ][ 57 ],
   alphaCSR[ 18 ][ 58 ],
   alphaCSR[ 18 ][ 59 ],
   alphaCSR[ 18 ][ 60 ],
   alphaCSR[ 18 ][ 61 ],
   alphaCSR[ 18 ][ 62 ],
   alphaCSR[ 18 ][ 63 ],
   alphaCSR[ 18 ][ 64 ],
   alphaCSR[ 18 ][ 65 ],
   alphaCSR[ 18 ][ 66 ],
   alphaCSR[ 18 ][ 67 ],
   alphaCSR[ 18 ][ 68 ],
   alphaCSR[ 18 ][ 69 ],
   alphaCSR[ 18 ][ 70 ],
   alphaCSR[ 18 ][ 71 ],
   alphaCSR[ 18 ][ 72 ],
   alphaCSR[ 18 ][ 73 ],
   alphaCSR[ 18 ][ 74 ],
   alphaCSR[ 18 ][ 75 ],
   alphaCSR[ 18 ][ 76 ],
   alphaCSR[ 18 ][ 77 ],
   alphaCSR[ 18 ][ 78 ],
   alphaCSR[ 18 ][ 79 ],
   alphaCSR[ 18 ][ 80 ],
   alphaCSR[ 18 ][ 81 ],
   alphaCSR[ 18 ][ 82 ],
   alphaCSR[ 18 ][ 83 ],
   alphaCSR[ 18 ][ 84 ],
   alphaCSR[ 18 ][ 85 ],
   alphaCSR[ 18 ][ 86 ],
   alphaCSR[ 18 ][ 87 ],
   alphaCSR[ 18 ][ 88 ],
   alphaCSR[ 18 ][ 89 ],
   alphaCSR[ 18 ][ 90 ],
   alphaCSR[ 18 ][ 91 ],
   alphaCSR[ 18 ][ 92 ],
   alphaCSR[ 18 ][ 93 ],
   alphaCSR[ 18 ][ 94 ],
   alphaCSR[ 18 ][ 95 ],
   alphaCSR[ 18 ][ 96 ],
   alphaCSR[ 18 ][ 97 ],
   alphaCSR[ 18 ][ 98 ],
   alphaCSR[ 18 ][ 99 ],
   alphaCSR[ 18 ][ 100 ],
   alphaCSR[ 18 ][ 101 ],
   alphaCSR[ 18 ][ 102 ],
   alphaCSR[ 18 ][ 103 ],
   alphaCSR[ 18 ][ 104 ],
   alphaCSR[ 18 ][ 105 ],
   alphaCSR[ 18 ][ 106 ],
   alphaCSR[ 18 ][ 107 ],
   alphaCSR[ 18 ][ 108 ],
   alphaCSR[ 18 ][ 109 ],
   alphaCSR[ 18 ][ 110 ],
   alphaCSR[ 18 ][ 111 ],
   alphaCSR[ 18 ][ 112 ],
   alphaCSR[ 18 ][ 113 ],
   alphaCSR[ 18 ][ 114 ],
   alphaCSR[ 18 ][ 115 ],
   alphaCSR[ 18 ][ 116 ],
   alphaCSR[ 18 ][ 117 ],
   alphaCSR[ 18 ][ 118 ],
   alphaCSR[ 18 ][ 119 ],
   alphaCSR[ 18 ][ 120 ],
   alphaCSR[ 18 ][ 121 ],
   alphaCSR[ 18 ][ 122 ],
   alphaCSR[ 18 ][ 123 ],
   alphaCSR[ 18 ][ 124 ],
   alphaCSR[ 18 ][ 125 ],
   alphaCSR[ 18 ][ 126 ],
   alphaCSR[ 18 ][ 127 ],
   alphaCSR[ 18 ][ 128 ],
   alphaCSR[ 18 ][ 129 ],
   alphaCSR[ 18 ][ 130 ],
   alphaCSR[ 18 ][ 131 ],
   alphaCSR[ 18 ][ 132 ],
   alphaCSR[ 18 ][ 133 ],
   alphaCSR[ 18 ][ 134 ],
   alphaCSR[ 18 ][ 135 ],
   alphaCSR[ 18 ][ 136 ],
   alphaCSR[ 18 ][ 137 ],
   alphaCSR[ 18 ][ 138 ],
   alphaCSR[ 18 ][ 139 ],
   alphaCSR[ 18 ][ 140 ],
   alphaCSR[ 18 ][ 141 ],
   alphaCSR[ 18 ][ 142 ],
   alphaCSR[ 18 ][ 143 ],
   alphaCSR[ 18 ][ 144 ],
   alphaCSR[ 18 ][ 145 ],
   alphaCSR[ 18 ][ 146 ],
   alphaCSR[ 18 ][ 147 ],
   alphaCSR[ 18 ][ 148 ],
   alphaCSR[ 18 ][ 149 ],
   alphaCSR[ 18 ][ 150 ],
   alphaCSR[ 18 ][ 151 ],
   alphaCSR[ 18 ][ 152 ],
   alphaCSR[ 18 ][ 153 ],
   alphaCSR[ 18 ][ 154 ],
   alphaCSR[ 18 ][ 155 ],
   alphaCSR[ 18 ][ 156 ],
   alphaCSR[ 18 ][ 157 ],
   alphaCSR[ 18 ][ 158 ],
   alphaCSR[ 18 ][ 159 ],
   alphaCSR[ 18 ][ 160 ],
   alphaCSR[ 18 ][ 161 ],
   alphaCSR[ 18 ][ 162 ],
   alphaCSR[ 18 ][ 163 ],
   alphaCSR[ 18 ][ 164 ],
   alphaCSR[ 18 ][ 165 ],
   alphaCSR[ 18 ][ 166 ],
   alphaCSR[ 18 ][ 167 ],
   alphaCSR[ 18 ][ 168 ],
   alphaCSR[ 18 ][ 169 ],
   alphaCSR[ 18 ][ 170 ],
   alphaCSR[ 18 ][ 171 ],
   alphaCSR[ 18 ][ 172 ],
   alphaCSR[ 18 ][ 173 ],
   alphaCSR[ 18 ][ 174 ],
   alphaCSR[ 18 ][ 175 ],
   alphaCSR[ 18 ][ 176 ],
   alphaCSR[ 18 ][ 177 ],
   alphaCSR[ 18 ][ 178 ],
   alphaCSR[ 18 ][ 179 ],
   alphaCSR[ 18 ][ 180 ],
   alphaCSR[ 18 ][ 181 ],
   alphaCSR[ 18 ][ 182 ],
   alphaCSR[ 18 ][ 183 ],
   alphaCSR[ 18 ][ 184 ],
   alphaCSR[ 18 ][ 185 ],
   alphaCSR[ 18 ][ 186 ],
   alphaCSR[ 18 ][ 187 ],
   alphaCSR[ 18 ][ 188 ],
   alphaCSR[ 18 ][ 189 ],
   alphaCSR[ 18 ][ 190 ],
   alphaCSR[ 18 ][ 191 ],
   alphaCSR[ 18 ][ 192 ],
   alphaCSR[ 18 ][ 193 ],
   alphaCSR[ 18 ][ 194 ],
   alphaCSR[ 18 ][ 195 ],
   alphaCSR[ 18 ][ 196 ],
   alphaCSR[ 18 ][ 197 ],
   alphaCSR[ 18 ][ 198 ],
   alphaCSR[ 18 ][ 199 ],
   alphaCSR[ 18 ][ 200 ],
   alphaCSR[ 18 ][ 201 ],
   alphaCSR[ 18 ][ 202 ],
   alphaCSR[ 18 ][ 203 ],
   alphaCSR[ 18 ][ 204 ],
   alphaCSR[ 18 ][ 205 ],
   alphaCSR[ 18 ][ 206 ],
   alphaCSR[ 18 ][ 207 ],
   alphaCSR[ 18 ][ 208 ],
   alphaCSR[ 18 ][ 209 ],
   alphaCSR[ 18 ][ 210 ],
   alphaCSR[ 18 ][ 211 ],
   alphaCSR[ 18 ][ 212 ],
   alphaCSR[ 18 ][ 213 ],
   alphaCSR[ 18 ][ 214 ],
   alphaCSR[ 18 ][ 215 ],
   alphaCSR[ 18 ][ 216 ],
   alphaCSR[ 18 ][ 217 ],
   alphaCSR[ 18 ][ 218 ],
   alphaCSR[ 18 ][ 219 ],
   alphaCSR[ 18 ][ 220 ],
   alphaCSR[ 18 ][ 221 ],
   alphaCSR[ 18 ][ 222 ],
   alphaCSR[ 18 ][ 223 ],
   alphaCSR[ 18 ][ 224 ],
   alphaCSR[ 18 ][ 225 ],
   alphaCSR[ 18 ][ 226 ],
   alphaCSR[ 18 ][ 227 ],
   alphaCSR[ 18 ][ 228 ],
   alphaCSR[ 18 ][ 229 ],
   alphaCSR[ 18 ][ 230 ],
   alphaCSR[ 18 ][ 231 ],
   alphaCSR[ 18 ][ 232 ],
   alphaCSR[ 18 ][ 233 ],
   alphaCSR[ 18 ][ 234 ],
   alphaCSR[ 18 ][ 235 ],
   alphaCSR[ 18 ][ 236 ],
   alphaCSR[ 18 ][ 237 ],
   alphaCSR[ 18 ][ 238 ],
   alphaCSR[ 18 ][ 239 ],
   alphaCSR[ 18 ][ 240 ],
   alphaCSR[ 18 ][ 241 ],
   alphaCSR[ 18 ][ 242 ],
   alphaCSR[ 18 ][ 243 ],
   alphaCSR[ 18 ][ 244 ],
   alphaCSR[ 18 ][ 245 ],
   alphaCSR[ 18 ][ 246 ],
   alphaCSR[ 18 ][ 247 ],
   alphaCSR[ 18 ][ 248 ],
   alphaCSR[ 18 ][ 249 ],
   alphaCSR[ 18 ][ 250 ],
   alphaCSR[ 18 ][ 251 ],
   alphaCSR[ 18 ][ 252 ],
   alphaCSR[ 18 ][ 253 ],
   alphaCSR[ 18 ][ 254 ],
   alphaCSR[ 18 ][ 255 ],
   alphaCSR[ 18 ][ 256 ],
   alphaCSR[ 18 ][ 257 ],
   alphaCSR[ 18 ][ 258 ],
   alphaCSR[ 18 ][ 259 ],
   alphaCSR[ 18 ][ 260 ],
   alphaCSR[ 18 ][ 261 ],
   alphaCSR[ 18 ][ 262 ],
   alphaCSR[ 18 ][ 263 ],
   alphaCSR[ 18 ][ 264 ],
   alphaCSR[ 18 ][ 265 ],
   alphaCSR[ 18 ][ 266 ],
   alphaCSR[ 18 ][ 267 ],
   alphaCSR[ 18 ][ 268 ],
   alphaCSR[ 18 ][ 269 ],
   alphaCSR[ 18 ][ 270 ],
   alphaCSR[ 18 ][ 271 ],
   alphaCSR[ 18 ][ 272 ],
   alphaCSR[ 18 ][ 273 ],
   alphaCSR[ 18 ][ 274 ],
   alphaCSR[ 18 ][ 275 ],
   alphaCSR[ 18 ][ 276 ],
   alphaCSR[ 18 ][ 277 ],
   alphaCSR[ 18 ][ 278 ],
   alphaCSR[ 18 ][ 279 ],
   alphaCSR[ 18 ][ 280 ],
   alphaCSR[ 18 ][ 281 ],
   alphaCSR[ 18 ][ 282 ],
   alphaCSR[ 18 ][ 283 ],
   alphaCSR[ 18 ][ 284 ],
   alphaCSR[ 18 ][ 285 ],
   alphaCSR[ 18 ][ 286 ],
   alphaCSR[ 18 ][ 287 ],
   alphaCSR[ 18 ][ 288 ],
   alphaCSR[ 18 ][ 289 ],
   alphaCSR[ 18 ][ 290 ],
   alphaCSR[ 18 ][ 291 ],
   alphaCSR[ 18 ][ 292 ],
   alphaCSR[ 18 ][ 293 ],
   alphaCSR[ 18 ][ 294 ],
   alphaCSR[ 18 ][ 295 ],
   alphaCSR[ 18 ][ 296 ],
   alphaCSR[ 18 ][ 297 ],
   alphaCSR[ 18 ][ 298 ],
   alphaCSR[ 18 ][ 299 ],
   alphaCSR[ 18 ][ 300 ],
   alphaCSR[ 18 ][ 301 ],
   alphaCSR[ 18 ][ 302 ],
   alphaCSR[ 18 ][ 303 ],
   alphaCSR[ 18 ][ 304 ],
   alphaCSR[ 18 ][ 305 ],
   alphaCSR[ 18 ][ 306 ],
   alphaCSR[ 18 ][ 307 ],
   alphaCSR[ 18 ][ 308 ],
   alphaCSR[ 18 ][ 309 ],
   alphaCSR[ 18 ][ 310 ],
   alphaCSR[ 18 ][ 311 ],
   alphaCSR[ 18 ][ 312 ],
   alphaCSR[ 18 ][ 313 ],
   alphaCSR[ 18 ][ 314 ],
   alphaCSR[ 18 ][ 315 ],
   alphaCSR[ 18 ][ 316 ],
   alphaCSR[ 18 ][ 317 ],
   alphaCSR[ 18 ][ 318 ],
   alphaCSR[ 18 ][ 319 ],
   alphaCSR[ 18 ][ 320 ],
   alphaCSR[ 18 ][ 321 ],
   alphaCSR[ 18 ][ 322 ],
   alphaCSR[ 18 ][ 323 ],
   alphaCSR[ 18 ][ 324 ],
   alphaCSR[ 18 ][ 325 ],
   alphaCSR[ 18 ][ 326 ],
   alphaCSR[ 18 ][ 327 ],
   alphaCSR[ 18 ][ 328 ],
   alphaCSR[ 18 ][ 329 ],
   alphaCSR[ 18 ][ 330 ],
   alphaCSR[ 18 ][ 331 ],
   alphaCSR[ 18 ][ 332 ],
   alphaCSR[ 18 ][ 333 ],
   alphaCSR[ 18 ][ 334 ],
   alphaCSR[ 18 ][ 335 ],
   alphaCSR[ 18 ][ 336 ],
   alphaCSR[ 18 ][ 337 ],
   alphaCSR[ 18 ][ 338 ],
   alphaCSR[ 18 ][ 339 ],
   alphaCSR[ 18 ][ 340 ],
   alphaCSR[ 18 ][ 341 ],
   alphaCSR[ 18 ][ 342 ],
   alphaCSR[ 18 ][ 343 ],
   alphaCSR[ 18 ][ 344 ],
   alphaCSR[ 18 ][ 345 ],
   alphaCSR[ 18 ][ 346 ],
   alphaCSR[ 18 ][ 347 ],
   alphaCSR[ 18 ][ 348 ],
   alphaCSR[ 18 ][ 349 ],
   alphaCSR[ 18 ][ 350 ],
   alphaCSR[ 18 ][ 351 ],
   alphaCSR[ 18 ][ 352 ],
   alphaCSR[ 18 ][ 353 ],
   alphaCSR[ 18 ][ 354 ],
   alphaCSR[ 18 ][ 355 ],
   alphaCSR[ 18 ][ 356 ],
   alphaCSR[ 18 ][ 357 ],
   alphaCSR[ 18 ][ 358 ],
   alphaCSR[ 18 ][ 359 ],
   alphaCSR[ 18 ][ 360 ],
   alphaCSR[ 18 ][ 361 ],
   alphaCSR[ 18 ][ 362 ],
   alphaCSR[ 18 ][ 363 ],
   alphaCSR[ 18 ][ 364 ],
   alphaCSR[ 18 ][ 365 ],
   alphaCSR[ 18 ][ 366 ],
   alphaCSR[ 18 ][ 367 ],
   alphaCSR[ 18 ][ 368 ],
   alphaCSR[ 18 ][ 369 ],
   alphaCSR[ 18 ][ 370 ],
   alphaCSR[ 18 ][ 371 ],
   alphaCSR[ 18 ][ 372 ],
   alphaCSR[ 18 ][ 373 ],
   alphaCSR[ 18 ][ 374 ],
   alphaCSR[ 18 ][ 375 ],
   alphaCSR[ 18 ][ 376 ],
   alphaCSR[ 18 ][ 377 ],
   alphaCSR[ 18 ][ 378 ],
   alphaCSR[ 18 ][ 379 ],
   alphaCSR[ 18 ][ 380 ],
   alphaCSR[ 18 ][ 381 ],
   alphaCSR[ 18 ][ 382 ],
   alphaCSR[ 18 ][ 383 ],
   alphaCSR[ 19 ][ 0 ],
   alphaCSR[ 19 ][ 1 ],
   alphaCSR[ 19 ][ 2 ],
   alphaCSR[ 19 ][ 3 ],
   alphaCSR[ 19 ][ 4 ],
   alphaCSR[ 19 ][ 5 ],
   alphaCSR[ 19 ][ 6 ],
   alphaCSR[ 19 ][ 7 ],
   alphaCSR[ 19 ][ 8 ],
   alphaCSR[ 19 ][ 9 ],
   alphaCSR[ 19 ][ 10 ],
   alphaCSR[ 19 ][ 11 ],
   alphaCSR[ 19 ][ 12 ],
   alphaCSR[ 19 ][ 13 ],
   alphaCSR[ 19 ][ 14 ],
   alphaCSR[ 19 ][ 15 ],
   alphaCSR[ 19 ][ 16 ],
   alphaCSR[ 19 ][ 17 ],
   alphaCSR[ 19 ][ 18 ],
   alphaCSR[ 19 ][ 19 ],
   alphaCSR[ 19 ][ 20 ],
   alphaCSR[ 19 ][ 21 ],
   alphaCSR[ 19 ][ 22 ],
   alphaCSR[ 19 ][ 23 ],
   alphaCSR[ 19 ][ 24 ],
   alphaCSR[ 19 ][ 25 ],
   alphaCSR[ 19 ][ 26 ],
   alphaCSR[ 19 ][ 27 ],
   alphaCSR[ 19 ][ 28 ],
   alphaCSR[ 19 ][ 29 ],
   alphaCSR[ 19 ][ 30 ],
   alphaCSR[ 19 ][ 31 ],
   alphaCSR[ 19 ][ 32 ],
   alphaCSR[ 19 ][ 33 ],
   alphaCSR[ 19 ][ 34 ],
   alphaCSR[ 19 ][ 35 ],
   alphaCSR[ 19 ][ 36 ],
   alphaCSR[ 19 ][ 37 ],
   alphaCSR[ 19 ][ 38 ],
   alphaCSR[ 19 ][ 39 ],
   alphaCSR[ 19 ][ 40 ],
   alphaCSR[ 19 ][ 41 ],
   alphaCSR[ 19 ][ 42 ],
   alphaCSR[ 19 ][ 43 ],
   alphaCSR[ 19 ][ 44 ],
   alphaCSR[ 19 ][ 45 ],
   alphaCSR[ 19 ][ 46 ],
   alphaCSR[ 19 ][ 47 ],
   alphaCSR[ 19 ][ 48 ],
   alphaCSR[ 19 ][ 49 ],
   alphaCSR[ 19 ][ 50 ],
   alphaCSR[ 19 ][ 51 ],
   alphaCSR[ 19 ][ 52 ],
   alphaCSR[ 19 ][ 53 ],
   alphaCSR[ 19 ][ 54 ],
   alphaCSR[ 19 ][ 55 ],
   alphaCSR[ 19 ][ 56 ],
   alphaCSR[ 19 ][ 57 ],
   alphaCSR[ 19 ][ 58 ],
   alphaCSR[ 19 ][ 59 ],
   alphaCSR[ 19 ][ 60 ],
   alphaCSR[ 19 ][ 61 ],
   alphaCSR[ 19 ][ 62 ],
   alphaCSR[ 19 ][ 63 ],
   alphaCSR[ 19 ][ 64 ],
   alphaCSR[ 19 ][ 65 ],
   alphaCSR[ 19 ][ 66 ],
   alphaCSR[ 19 ][ 67 ],
   alphaCSR[ 19 ][ 68 ],
   alphaCSR[ 19 ][ 69 ],
   alphaCSR[ 19 ][ 70 ],
   alphaCSR[ 19 ][ 71 ],
   alphaCSR[ 19 ][ 72 ],
   alphaCSR[ 19 ][ 73 ],
   alphaCSR[ 19 ][ 74 ],
   alphaCSR[ 19 ][ 75 ],
   alphaCSR[ 19 ][ 76 ],
   alphaCSR[ 19 ][ 77 ],
   alphaCSR[ 19 ][ 78 ],
   alphaCSR[ 19 ][ 79 ],
   alphaCSR[ 19 ][ 80 ],
   alphaCSR[ 19 ][ 81 ],
   alphaCSR[ 19 ][ 82 ],
   alphaCSR[ 19 ][ 83 ],
   alphaCSR[ 19 ][ 84 ],
   alphaCSR[ 19 ][ 85 ],
   alphaCSR[ 19 ][ 86 ],
   alphaCSR[ 19 ][ 87 ],
   alphaCSR[ 19 ][ 88 ],
   alphaCSR[ 19 ][ 89 ],
   alphaCSR[ 19 ][ 90 ],
   alphaCSR[ 19 ][ 91 ],
   alphaCSR[ 19 ][ 92 ],
   alphaCSR[ 19 ][ 93 ],
   alphaCSR[ 19 ][ 94 ],
   alphaCSR[ 19 ][ 95 ],
   alphaCSR[ 19 ][ 96 ],
   alphaCSR[ 19 ][ 97 ],
   alphaCSR[ 19 ][ 98 ],
   alphaCSR[ 19 ][ 99 ],
   alphaCSR[ 19 ][ 100 ],
   alphaCSR[ 19 ][ 101 ],
   alphaCSR[ 19 ][ 102 ],
   alphaCSR[ 19 ][ 103 ],
   alphaCSR[ 19 ][ 104 ],
   alphaCSR[ 19 ][ 105 ],
   alphaCSR[ 19 ][ 106 ],
   alphaCSR[ 19 ][ 107 ],
   alphaCSR[ 19 ][ 108 ],
   alphaCSR[ 19 ][ 109 ],
   alphaCSR[ 19 ][ 110 ],
   alphaCSR[ 19 ][ 111 ],
   alphaCSR[ 19 ][ 112 ],
   alphaCSR[ 19 ][ 113 ],
   alphaCSR[ 19 ][ 114 ],
   alphaCSR[ 19 ][ 115 ],
   alphaCSR[ 19 ][ 116 ],
   alphaCSR[ 19 ][ 117 ],
   alphaCSR[ 19 ][ 118 ],
   alphaCSR[ 19 ][ 119 ],
   alphaCSR[ 19 ][ 120 ],
   alphaCSR[ 19 ][ 121 ],
   alphaCSR[ 19 ][ 122 ],
   alphaCSR[ 19 ][ 123 ],
   alphaCSR[ 19 ][ 124 ],
   alphaCSR[ 19 ][ 125 ],
   alphaCSR[ 19 ][ 126 ],
   alphaCSR[ 19 ][ 127 ],
   alphaCSR[ 19 ][ 128 ],
   alphaCSR[ 19 ][ 129 ],
   alphaCSR[ 19 ][ 130 ],
   alphaCSR[ 19 ][ 131 ],
   alphaCSR[ 19 ][ 132 ],
   alphaCSR[ 19 ][ 133 ],
   alphaCSR[ 19 ][ 134 ],
   alphaCSR[ 19 ][ 135 ],
   alphaCSR[ 19 ][ 136 ],
   alphaCSR[ 19 ][ 137 ],
   alphaCSR[ 19 ][ 138 ],
   alphaCSR[ 19 ][ 139 ],
   alphaCSR[ 19 ][ 140 ],
   alphaCSR[ 19 ][ 141 ],
   alphaCSR[ 19 ][ 142 ],
   alphaCSR[ 19 ][ 143 ],
   alphaCSR[ 19 ][ 144 ],
   alphaCSR[ 19 ][ 145 ],
   alphaCSR[ 19 ][ 146 ],
   alphaCSR[ 19 ][ 147 ],
   alphaCSR[ 19 ][ 148 ],
   alphaCSR[ 19 ][ 149 ],
   alphaCSR[ 19 ][ 150 ],
   alphaCSR[ 19 ][ 151 ],
   alphaCSR[ 19 ][ 152 ],
   alphaCSR[ 19 ][ 153 ],
   alphaCSR[ 19 ][ 154 ],
   alphaCSR[ 19 ][ 155 ],
   alphaCSR[ 19 ][ 156 ],
   alphaCSR[ 19 ][ 157 ],
   alphaCSR[ 19 ][ 158 ],
   alphaCSR[ 19 ][ 159 ],
   alphaCSR[ 19 ][ 160 ],
   alphaCSR[ 19 ][ 161 ],
   alphaCSR[ 19 ][ 162 ],
   alphaCSR[ 19 ][ 163 ],
   alphaCSR[ 19 ][ 164 ],
   alphaCSR[ 19 ][ 165 ],
   alphaCSR[ 19 ][ 166 ],
   alphaCSR[ 19 ][ 167 ],
   alphaCSR[ 19 ][ 168 ],
   alphaCSR[ 19 ][ 169 ],
   alphaCSR[ 19 ][ 170 ],
   alphaCSR[ 19 ][ 171 ],
   alphaCSR[ 19 ][ 172 ],
   alphaCSR[ 19 ][ 173 ],
   alphaCSR[ 19 ][ 174 ],
   alphaCSR[ 19 ][ 175 ],
   alphaCSR[ 19 ][ 176 ],
   alphaCSR[ 19 ][ 177 ],
   alphaCSR[ 19 ][ 178 ],
   alphaCSR[ 19 ][ 179 ],
   alphaCSR[ 19 ][ 180 ],
   alphaCSR[ 19 ][ 181 ],
   alphaCSR[ 19 ][ 182 ],
   alphaCSR[ 19 ][ 183 ],
   alphaCSR[ 19 ][ 184 ],
   alphaCSR[ 19 ][ 185 ],
   alphaCSR[ 19 ][ 186 ],
   alphaCSR[ 19 ][ 187 ],
   alphaCSR[ 19 ][ 188 ],
   alphaCSR[ 19 ][ 189 ],
   alphaCSR[ 19 ][ 190 ],
   alphaCSR[ 19 ][ 191 ],
   alphaCSR[ 19 ][ 192 ],
   alphaCSR[ 19 ][ 193 ],
   alphaCSR[ 19 ][ 194 ],
   alphaCSR[ 19 ][ 195 ],
   alphaCSR[ 19 ][ 196 ],
   alphaCSR[ 19 ][ 197 ],
   alphaCSR[ 19 ][ 198 ],
   alphaCSR[ 19 ][ 199 ],
   alphaCSR[ 19 ][ 200 ],
   alphaCSR[ 19 ][ 201 ],
   alphaCSR[ 19 ][ 202 ],
   alphaCSR[ 19 ][ 203 ],
   alphaCSR[ 19 ][ 204 ],
   alphaCSR[ 19 ][ 205 ],
   alphaCSR[ 19 ][ 206 ],
   alphaCSR[ 19 ][ 207 ],
   alphaCSR[ 19 ][ 208 ],
   alphaCSR[ 19 ][ 209 ],
   alphaCSR[ 19 ][ 210 ],
   alphaCSR[ 19 ][ 211 ],
   alphaCSR[ 19 ][ 212 ],
   alphaCSR[ 19 ][ 213 ],
   alphaCSR[ 19 ][ 214 ],
   alphaCSR[ 19 ][ 215 ],
   alphaCSR[ 19 ][ 216 ],
   alphaCSR[ 19 ][ 217 ],
   alphaCSR[ 19 ][ 218 ],
   alphaCSR[ 19 ][ 219 ],
   alphaCSR[ 19 ][ 220 ],
   alphaCSR[ 19 ][ 221 ],
   alphaCSR[ 19 ][ 222 ],
   alphaCSR[ 19 ][ 223 ],
   alphaCSR[ 19 ][ 224 ],
   alphaCSR[ 19 ][ 225 ],
   alphaCSR[ 19 ][ 226 ],
   alphaCSR[ 19 ][ 227 ],
   alphaCSR[ 19 ][ 228 ],
   alphaCSR[ 19 ][ 229 ],
   alphaCSR[ 19 ][ 230 ],
   alphaCSR[ 19 ][ 231 ],
   alphaCSR[ 19 ][ 232 ],
   alphaCSR[ 19 ][ 233 ],
   alphaCSR[ 19 ][ 234 ],
   alphaCSR[ 19 ][ 235 ],
   alphaCSR[ 19 ][ 236 ],
   alphaCSR[ 19 ][ 237 ],
   alphaCSR[ 19 ][ 238 ],
   alphaCSR[ 19 ][ 239 ],
   alphaCSR[ 19 ][ 240 ],
   alphaCSR[ 19 ][ 241 ],
   alphaCSR[ 19 ][ 242 ],
   alphaCSR[ 19 ][ 243 ],
   alphaCSR[ 19 ][ 244 ],
   alphaCSR[ 19 ][ 245 ],
   alphaCSR[ 19 ][ 246 ],
   alphaCSR[ 19 ][ 247 ],
   alphaCSR[ 19 ][ 248 ],
   alphaCSR[ 19 ][ 249 ],
   alphaCSR[ 19 ][ 250 ],
   alphaCSR[ 19 ][ 251 ],
   alphaCSR[ 19 ][ 252 ],
   alphaCSR[ 19 ][ 253 ],
   alphaCSR[ 19 ][ 254 ],
   alphaCSR[ 19 ][ 255 ],
   alphaCSR[ 19 ][ 256 ],
   alphaCSR[ 19 ][ 257 ],
   alphaCSR[ 19 ][ 258 ],
   alphaCSR[ 19 ][ 259 ],
   alphaCSR[ 19 ][ 260 ],
   alphaCSR[ 19 ][ 261 ],
   alphaCSR[ 19 ][ 262 ],
   alphaCSR[ 19 ][ 263 ],
   alphaCSR[ 19 ][ 264 ],
   alphaCSR[ 19 ][ 265 ],
   alphaCSR[ 19 ][ 266 ],
   alphaCSR[ 19 ][ 267 ],
   alphaCSR[ 19 ][ 268 ],
   alphaCSR[ 19 ][ 269 ],
   alphaCSR[ 19 ][ 270 ],
   alphaCSR[ 19 ][ 271 ],
   alphaCSR[ 19 ][ 272 ],
   alphaCSR[ 19 ][ 273 ],
   alphaCSR[ 19 ][ 274 ],
   alphaCSR[ 19 ][ 275 ],
   alphaCSR[ 19 ][ 276 ],
   alphaCSR[ 19 ][ 277 ],
   alphaCSR[ 19 ][ 278 ],
   alphaCSR[ 19 ][ 279 ],
   alphaCSR[ 19 ][ 280 ],
   alphaCSR[ 19 ][ 281 ],
   alphaCSR[ 19 ][ 282 ],
   alphaCSR[ 19 ][ 283 ],
   alphaCSR[ 19 ][ 284 ],
   alphaCSR[ 19 ][ 285 ],
   alphaCSR[ 19 ][ 286 ],
   alphaCSR[ 19 ][ 287 ],
   alphaCSR[ 19 ][ 288 ],
   alphaCSR[ 19 ][ 289 ],
   alphaCSR[ 19 ][ 290 ],
   alphaCSR[ 19 ][ 291 ],
   alphaCSR[ 19 ][ 292 ],
   alphaCSR[ 19 ][ 293 ],
   alphaCSR[ 19 ][ 294 ],
   alphaCSR[ 19 ][ 295 ],
   alphaCSR[ 19 ][ 296 ],
   alphaCSR[ 19 ][ 297 ],
   alphaCSR[ 19 ][ 298 ],
   alphaCSR[ 19 ][ 299 ],
   alphaCSR[ 19 ][ 300 ],
   alphaCSR[ 19 ][ 301 ],
   alphaCSR[ 19 ][ 302 ],
   alphaCSR[ 19 ][ 303 ],
   alphaCSR[ 19 ][ 304 ],
   alphaCSR[ 19 ][ 305 ],
   alphaCSR[ 19 ][ 306 ],
   alphaCSR[ 19 ][ 307 ],
   alphaCSR[ 19 ][ 308 ],
   alphaCSR[ 19 ][ 309 ],
   alphaCSR[ 19 ][ 310 ],
   alphaCSR[ 19 ][ 311 ],
   alphaCSR[ 19 ][ 312 ],
   alphaCSR[ 19 ][ 313 ],
   alphaCSR[ 19 ][ 314 ],
   alphaCSR[ 19 ][ 315 ],
   alphaCSR[ 19 ][ 316 ],
   alphaCSR[ 19 ][ 317 ],
   alphaCSR[ 19 ][ 318 ],
   alphaCSR[ 19 ][ 319 ],
   alphaCSR[ 19 ][ 320 ],
   alphaCSR[ 19 ][ 321 ],
   alphaCSR[ 19 ][ 322 ],
   alphaCSR[ 19 ][ 323 ],
   alphaCSR[ 19 ][ 324 ],
   alphaCSR[ 19 ][ 325 ],
   alphaCSR[ 19 ][ 326 ],
   alphaCSR[ 19 ][ 327 ],
   alphaCSR[ 19 ][ 328 ],
   alphaCSR[ 19 ][ 329 ],
   alphaCSR[ 19 ][ 330 ],
   alphaCSR[ 19 ][ 331 ],
   alphaCSR[ 19 ][ 332 ],
   alphaCSR[ 19 ][ 333 ],
   alphaCSR[ 19 ][ 334 ],
   alphaCSR[ 19 ][ 335 ],
   alphaCSR[ 19 ][ 336 ],
   alphaCSR[ 19 ][ 337 ],
   alphaCSR[ 19 ][ 338 ],
   alphaCSR[ 19 ][ 339 ],
   alphaCSR[ 19 ][ 340 ],
   alphaCSR[ 19 ][ 341 ],
   alphaCSR[ 19 ][ 342 ],
   alphaCSR[ 19 ][ 343 ],
   alphaCSR[ 19 ][ 344 ],
   alphaCSR[ 19 ][ 345 ],
   alphaCSR[ 19 ][ 346 ],
   alphaCSR[ 19 ][ 347 ],
   alphaCSR[ 19 ][ 348 ],
   alphaCSR[ 19 ][ 349 ],
   alphaCSR[ 19 ][ 350 ],
   alphaCSR[ 19 ][ 351 ],
   alphaCSR[ 19 ][ 352 ],
   alphaCSR[ 19 ][ 353 ],
   alphaCSR[ 19 ][ 354 ],
   alphaCSR[ 19 ][ 355 ],
   alphaCSR[ 19 ][ 356 ],
   alphaCSR[ 19 ][ 357 ],
   alphaCSR[ 19 ][ 358 ],
   alphaCSR[ 19 ][ 359 ],
   alphaCSR[ 19 ][ 360 ],
   alphaCSR[ 19 ][ 361 ],
   alphaCSR[ 19 ][ 362 ],
   alphaCSR[ 19 ][ 363 ],
   alphaCSR[ 19 ][ 364 ],
   alphaCSR[ 19 ][ 365 ],
   alphaCSR[ 19 ][ 366 ],
   alphaCSR[ 19 ][ 367 ],
   alphaCSR[ 19 ][ 368 ],
   alphaCSR[ 19 ][ 369 ],
   alphaCSR[ 19 ][ 370 ],
   alphaCSR[ 19 ][ 371 ],
   alphaCSR[ 19 ][ 372 ],
   alphaCSR[ 19 ][ 373 ],
   alphaCSR[ 19 ][ 374 ],
   alphaCSR[ 19 ][ 375 ],
   alphaCSR[ 19 ][ 376 ],
   alphaCSR[ 19 ][ 377 ],
   alphaCSR[ 19 ][ 378 ],
   alphaCSR[ 19 ][ 379 ],
   alphaCSR[ 19 ][ 380 ],
   alphaCSR[ 19 ][ 381 ],
   alphaCSR[ 19 ][ 382 ],
   alphaCSR[ 19 ][ 383 ],
   alphaCSR[ 20 ][ 0 ],
   alphaCSR[ 20 ][ 1 ],
   alphaCSR[ 20 ][ 2 ],
   alphaCSR[ 20 ][ 3 ],
   alphaCSR[ 20 ][ 4 ],
   alphaCSR[ 20 ][ 5 ],
   alphaCSR[ 20 ][ 6 ],
   alphaCSR[ 20 ][ 7 ],
   alphaCSR[ 20 ][ 8 ],
   alphaCSR[ 20 ][ 9 ],
   alphaCSR[ 20 ][ 10 ],
   alphaCSR[ 20 ][ 11 ],
   alphaCSR[ 20 ][ 12 ],
   alphaCSR[ 20 ][ 13 ],
   alphaCSR[ 20 ][ 14 ],
   alphaCSR[ 20 ][ 15 ],
   alphaCSR[ 20 ][ 16 ],
   alphaCSR[ 20 ][ 17 ],
   alphaCSR[ 20 ][ 18 ],
   alphaCSR[ 20 ][ 19 ],
   alphaCSR[ 20 ][ 20 ],
   alphaCSR[ 20 ][ 21 ],
   alphaCSR[ 20 ][ 22 ],
   alphaCSR[ 20 ][ 23 ],
   alphaCSR[ 20 ][ 24 ],
   alphaCSR[ 20 ][ 25 ],
   alphaCSR[ 20 ][ 26 ],
   alphaCSR[ 20 ][ 27 ],
   alphaCSR[ 20 ][ 28 ],
   alphaCSR[ 20 ][ 29 ],
   alphaCSR[ 20 ][ 30 ],
   alphaCSR[ 20 ][ 31 ],
   alphaCSR[ 20 ][ 32 ],
   alphaCSR[ 20 ][ 33 ],
   alphaCSR[ 20 ][ 34 ],
   alphaCSR[ 20 ][ 35 ],
   alphaCSR[ 20 ][ 36 ],
   alphaCSR[ 20 ][ 37 ],
   alphaCSR[ 20 ][ 38 ],
   alphaCSR[ 20 ][ 39 ],
   alphaCSR[ 20 ][ 40 ],
   alphaCSR[ 20 ][ 41 ],
   alphaCSR[ 20 ][ 42 ],
   alphaCSR[ 20 ][ 43 ],
   alphaCSR[ 20 ][ 44 ],
   alphaCSR[ 20 ][ 45 ],
   alphaCSR[ 20 ][ 46 ],
   alphaCSR[ 20 ][ 47 ],
   alphaCSR[ 20 ][ 48 ],
   alphaCSR[ 20 ][ 49 ],
   alphaCSR[ 20 ][ 50 ],
   alphaCSR[ 20 ][ 51 ],
   alphaCSR[ 20 ][ 52 ],
   alphaCSR[ 20 ][ 53 ],
   alphaCSR[ 20 ][ 54 ],
   alphaCSR[ 20 ][ 55 ],
   alphaCSR[ 20 ][ 56 ],
   alphaCSR[ 20 ][ 57 ],
   alphaCSR[ 20 ][ 58 ],
   alphaCSR[ 20 ][ 59 ],
   alphaCSR[ 20 ][ 60 ],
   alphaCSR[ 20 ][ 61 ],
   alphaCSR[ 20 ][ 62 ],
   alphaCSR[ 20 ][ 63 ],
   alphaCSR[ 20 ][ 64 ],
   alphaCSR[ 20 ][ 65 ],
   alphaCSR[ 20 ][ 66 ],
   alphaCSR[ 20 ][ 67 ],
   alphaCSR[ 20 ][ 68 ],
   alphaCSR[ 20 ][ 69 ],
   alphaCSR[ 20 ][ 70 ],
   alphaCSR[ 20 ][ 71 ],
   alphaCSR[ 20 ][ 72 ],
   alphaCSR[ 20 ][ 73 ],
   alphaCSR[ 20 ][ 74 ],
   alphaCSR[ 20 ][ 75 ],
   alphaCSR[ 20 ][ 76 ],
   alphaCSR[ 20 ][ 77 ],
   alphaCSR[ 20 ][ 78 ],
   alphaCSR[ 20 ][ 79 ],
   alphaCSR[ 20 ][ 80 ],
   alphaCSR[ 20 ][ 81 ],
   alphaCSR[ 20 ][ 82 ],
   alphaCSR[ 20 ][ 83 ],
   alphaCSR[ 20 ][ 84 ],
   alphaCSR[ 20 ][ 85 ],
   alphaCSR[ 20 ][ 86 ],
   alphaCSR[ 20 ][ 87 ],
   alphaCSR[ 20 ][ 88 ],
   alphaCSR[ 20 ][ 89 ],
   alphaCSR[ 20 ][ 90 ],
   alphaCSR[ 20 ][ 91 ],
   alphaCSR[ 20 ][ 92 ],
   alphaCSR[ 20 ][ 93 ],
   alphaCSR[ 20 ][ 94 ],
   alphaCSR[ 20 ][ 95 ],
   alphaCSR[ 20 ][ 96 ],
   alphaCSR[ 20 ][ 97 ],
   alphaCSR[ 20 ][ 98 ],
   alphaCSR[ 20 ][ 99 ],
   alphaCSR[ 20 ][ 100 ],
   alphaCSR[ 20 ][ 101 ],
   alphaCSR[ 20 ][ 102 ],
   alphaCSR[ 20 ][ 103 ],
   alphaCSR[ 20 ][ 104 ],
   alphaCSR[ 20 ][ 105 ],
   alphaCSR[ 20 ][ 106 ],
   alphaCSR[ 20 ][ 107 ],
   alphaCSR[ 20 ][ 108 ],
   alphaCSR[ 20 ][ 109 ],
   alphaCSR[ 20 ][ 110 ],
   alphaCSR[ 20 ][ 111 ],
   alphaCSR[ 20 ][ 112 ],
   alphaCSR[ 20 ][ 113 ],
   alphaCSR[ 20 ][ 114 ],
   alphaCSR[ 20 ][ 115 ],
   alphaCSR[ 20 ][ 116 ],
   alphaCSR[ 20 ][ 117 ],
   alphaCSR[ 20 ][ 118 ],
   alphaCSR[ 20 ][ 119 ],
   alphaCSR[ 20 ][ 120 ],
   alphaCSR[ 20 ][ 121 ],
   alphaCSR[ 20 ][ 122 ],
   alphaCSR[ 20 ][ 123 ],
   alphaCSR[ 20 ][ 124 ],
   alphaCSR[ 20 ][ 125 ],
   alphaCSR[ 20 ][ 126 ],
   alphaCSR[ 20 ][ 127 ],
   alphaCSR[ 20 ][ 128 ],
   alphaCSR[ 20 ][ 129 ],
   alphaCSR[ 20 ][ 130 ],
   alphaCSR[ 20 ][ 131 ],
   alphaCSR[ 20 ][ 132 ],
   alphaCSR[ 20 ][ 133 ],
   alphaCSR[ 20 ][ 134 ],
   alphaCSR[ 20 ][ 135 ],
   alphaCSR[ 20 ][ 136 ],
   alphaCSR[ 20 ][ 137 ],
   alphaCSR[ 20 ][ 138 ],
   alphaCSR[ 20 ][ 139 ],
   alphaCSR[ 20 ][ 140 ],
   alphaCSR[ 20 ][ 141 ],
   alphaCSR[ 20 ][ 142 ],
   alphaCSR[ 20 ][ 143 ],
   alphaCSR[ 20 ][ 144 ],
   alphaCSR[ 20 ][ 145 ],
   alphaCSR[ 20 ][ 146 ],
   alphaCSR[ 20 ][ 147 ],
   alphaCSR[ 20 ][ 148 ],
   alphaCSR[ 20 ][ 149 ],
   alphaCSR[ 20 ][ 150 ],
   alphaCSR[ 20 ][ 151 ],
   alphaCSR[ 20 ][ 152 ],
   alphaCSR[ 20 ][ 153 ],
   alphaCSR[ 20 ][ 154 ],
   alphaCSR[ 20 ][ 155 ],
   alphaCSR[ 20 ][ 156 ],
   alphaCSR[ 20 ][ 157 ],
   alphaCSR[ 20 ][ 158 ],
   alphaCSR[ 20 ][ 159 ],
   alphaCSR[ 20 ][ 160 ],
   alphaCSR[ 20 ][ 161 ],
   alphaCSR[ 20 ][ 162 ],
   alphaCSR[ 20 ][ 163 ],
   alphaCSR[ 20 ][ 164 ],
   alphaCSR[ 20 ][ 165 ],
   alphaCSR[ 20 ][ 166 ],
   alphaCSR[ 20 ][ 167 ],
   alphaCSR[ 20 ][ 168 ],
   alphaCSR[ 20 ][ 169 ],
   alphaCSR[ 20 ][ 170 ],
   alphaCSR[ 20 ][ 171 ],
   alphaCSR[ 20 ][ 172 ],
   alphaCSR[ 20 ][ 173 ],
   alphaCSR[ 20 ][ 174 ],
   alphaCSR[ 20 ][ 175 ],
   alphaCSR[ 20 ][ 176 ],
   alphaCSR[ 20 ][ 177 ],
   alphaCSR[ 20 ][ 178 ],
   alphaCSR[ 20 ][ 179 ],
   alphaCSR[ 20 ][ 180 ],
   alphaCSR[ 20 ][ 181 ],
   alphaCSR[ 20 ][ 182 ],
   alphaCSR[ 20 ][ 183 ],
   alphaCSR[ 20 ][ 184 ],
   alphaCSR[ 20 ][ 185 ],
   alphaCSR[ 20 ][ 186 ],
   alphaCSR[ 20 ][ 187 ],
   alphaCSR[ 20 ][ 188 ],
   alphaCSR[ 20 ][ 189 ],
   alphaCSR[ 20 ][ 190 ],
   alphaCSR[ 20 ][ 191 ],
   alphaCSR[ 20 ][ 192 ],
   alphaCSR[ 20 ][ 193 ],
   alphaCSR[ 20 ][ 194 ],
   alphaCSR[ 20 ][ 195 ],
   alphaCSR[ 20 ][ 196 ],
   alphaCSR[ 20 ][ 197 ],
   alphaCSR[ 20 ][ 198 ],
   alphaCSR[ 20 ][ 199 ],
   alphaCSR[ 20 ][ 200 ],
   alphaCSR[ 20 ][ 201 ],
   alphaCSR[ 20 ][ 202 ],
   alphaCSR[ 20 ][ 203 ],
   alphaCSR[ 20 ][ 204 ],
   alphaCSR[ 20 ][ 205 ],
   alphaCSR[ 20 ][ 206 ],
   alphaCSR[ 20 ][ 207 ],
   alphaCSR[ 20 ][ 208 ],
   alphaCSR[ 20 ][ 209 ],
   alphaCSR[ 20 ][ 210 ],
   alphaCSR[ 20 ][ 211 ],
   alphaCSR[ 20 ][ 212 ],
   alphaCSR[ 20 ][ 213 ],
   alphaCSR[ 20 ][ 214 ],
   alphaCSR[ 20 ][ 215 ],
   alphaCSR[ 20 ][ 216 ],
   alphaCSR[ 20 ][ 217 ],
   alphaCSR[ 20 ][ 218 ],
   alphaCSR[ 20 ][ 219 ],
   alphaCSR[ 20 ][ 220 ],
   alphaCSR[ 20 ][ 221 ],
   alphaCSR[ 20 ][ 222 ],
   alphaCSR[ 20 ][ 223 ],
   alphaCSR[ 20 ][ 224 ],
   alphaCSR[ 20 ][ 225 ],
   alphaCSR[ 20 ][ 226 ],
   alphaCSR[ 20 ][ 227 ],
   alphaCSR[ 20 ][ 228 ],
   alphaCSR[ 20 ][ 229 ],
   alphaCSR[ 20 ][ 230 ],
   alphaCSR[ 20 ][ 231 ],
   alphaCSR[ 20 ][ 232 ],
   alphaCSR[ 20 ][ 233 ],
   alphaCSR[ 20 ][ 234 ],
   alphaCSR[ 20 ][ 235 ],
   alphaCSR[ 20 ][ 236 ],
   alphaCSR[ 20 ][ 237 ],
   alphaCSR[ 20 ][ 238 ],
   alphaCSR[ 20 ][ 239 ],
   alphaCSR[ 20 ][ 240 ],
   alphaCSR[ 20 ][ 241 ],
   alphaCSR[ 20 ][ 242 ],
   alphaCSR[ 20 ][ 243 ],
   alphaCSR[ 20 ][ 244 ],
   alphaCSR[ 20 ][ 245 ],
   alphaCSR[ 20 ][ 246 ],
   alphaCSR[ 20 ][ 247 ],
   alphaCSR[ 20 ][ 248 ],
   alphaCSR[ 20 ][ 249 ],
   alphaCSR[ 20 ][ 250 ],
   alphaCSR[ 20 ][ 251 ],
   alphaCSR[ 20 ][ 252 ],
   alphaCSR[ 20 ][ 253 ],
   alphaCSR[ 20 ][ 254 ],
   alphaCSR[ 20 ][ 255 ],
   alphaCSR[ 20 ][ 256 ],
   alphaCSR[ 20 ][ 257 ],
   alphaCSR[ 20 ][ 258 ],
   alphaCSR[ 20 ][ 259 ],
   alphaCSR[ 20 ][ 260 ],
   alphaCSR[ 20 ][ 261 ],
   alphaCSR[ 20 ][ 262 ],
   alphaCSR[ 20 ][ 263 ],
   alphaCSR[ 20 ][ 264 ],
   alphaCSR[ 20 ][ 265 ],
   alphaCSR[ 20 ][ 266 ],
   alphaCSR[ 20 ][ 267 ],
   alphaCSR[ 20 ][ 268 ],
   alphaCSR[ 20 ][ 269 ],
   alphaCSR[ 20 ][ 270 ],
   alphaCSR[ 20 ][ 271 ],
   alphaCSR[ 20 ][ 272 ],
   alphaCSR[ 20 ][ 273 ],
   alphaCSR[ 20 ][ 274 ],
   alphaCSR[ 20 ][ 275 ],
   alphaCSR[ 20 ][ 276 ],
   alphaCSR[ 20 ][ 277 ],
   alphaCSR[ 20 ][ 278 ],
   alphaCSR[ 20 ][ 279 ],
   alphaCSR[ 20 ][ 280 ],
   alphaCSR[ 20 ][ 281 ],
   alphaCSR[ 20 ][ 282 ],
   alphaCSR[ 20 ][ 283 ],
   alphaCSR[ 20 ][ 284 ],
   alphaCSR[ 20 ][ 285 ],
   alphaCSR[ 20 ][ 286 ],
   alphaCSR[ 20 ][ 287 ],
   alphaCSR[ 20 ][ 288 ],
   alphaCSR[ 20 ][ 289 ],
   alphaCSR[ 20 ][ 290 ],
   alphaCSR[ 20 ][ 291 ],
   alphaCSR[ 20 ][ 292 ],
   alphaCSR[ 20 ][ 293 ],
   alphaCSR[ 20 ][ 294 ],
   alphaCSR[ 20 ][ 295 ],
   alphaCSR[ 20 ][ 296 ],
   alphaCSR[ 20 ][ 297 ],
   alphaCSR[ 20 ][ 298 ],
   alphaCSR[ 20 ][ 299 ],
   alphaCSR[ 20 ][ 300 ],
   alphaCSR[ 20 ][ 301 ],
   alphaCSR[ 20 ][ 302 ],
   alphaCSR[ 20 ][ 303 ],
   alphaCSR[ 20 ][ 304 ],
   alphaCSR[ 20 ][ 305 ],
   alphaCSR[ 20 ][ 306 ],
   alphaCSR[ 20 ][ 307 ],
   alphaCSR[ 20 ][ 308 ],
   alphaCSR[ 20 ][ 309 ],
   alphaCSR[ 20 ][ 310 ],
   alphaCSR[ 20 ][ 311 ],
   alphaCSR[ 20 ][ 312 ],
   alphaCSR[ 20 ][ 313 ],
   alphaCSR[ 20 ][ 314 ],
   alphaCSR[ 20 ][ 315 ],
   alphaCSR[ 20 ][ 316 ],
   alphaCSR[ 20 ][ 317 ],
   alphaCSR[ 20 ][ 318 ],
   alphaCSR[ 20 ][ 319 ],
   alphaCSR[ 20 ][ 320 ],
   alphaCSR[ 20 ][ 321 ],
   alphaCSR[ 20 ][ 322 ],
   alphaCSR[ 20 ][ 323 ],
   alphaCSR[ 20 ][ 324 ],
   alphaCSR[ 20 ][ 325 ],
   alphaCSR[ 20 ][ 326 ],
   alphaCSR[ 20 ][ 327 ],
   alphaCSR[ 20 ][ 328 ],
   alphaCSR[ 20 ][ 329 ],
   alphaCSR[ 20 ][ 330 ],
   alphaCSR[ 20 ][ 331 ],
   alphaCSR[ 20 ][ 332 ],
   alphaCSR[ 20 ][ 333 ],
   alphaCSR[ 20 ][ 334 ],
   alphaCSR[ 20 ][ 335 ],
   alphaCSR[ 20 ][ 336 ],
   alphaCSR[ 20 ][ 337 ],
   alphaCSR[ 20 ][ 338 ],
   alphaCSR[ 20 ][ 339 ],
   alphaCSR[ 20 ][ 340 ],
   alphaCSR[ 20 ][ 341 ],
   alphaCSR[ 20 ][ 342 ],
   alphaCSR[ 20 ][ 343 ],
   alphaCSR[ 20 ][ 344 ],
   alphaCSR[ 20 ][ 345 ],
   alphaCSR[ 20 ][ 346 ],
   alphaCSR[ 20 ][ 347 ],
   alphaCSR[ 20 ][ 348 ],
   alphaCSR[ 20 ][ 349 ],
   alphaCSR[ 20 ][ 350 ],
   alphaCSR[ 20 ][ 351 ],
   alphaCSR[ 20 ][ 352 ],
   alphaCSR[ 20 ][ 353 ],
   alphaCSR[ 20 ][ 354 ],
   alphaCSR[ 20 ][ 355 ],
   alphaCSR[ 20 ][ 356 ],
   alphaCSR[ 20 ][ 357 ],
   alphaCSR[ 20 ][ 358 ],
   alphaCSR[ 20 ][ 359 ],
   alphaCSR[ 20 ][ 360 ],
   alphaCSR[ 20 ][ 361 ],
   alphaCSR[ 20 ][ 362 ],
   alphaCSR[ 20 ][ 363 ],
   alphaCSR[ 20 ][ 364 ],
   alphaCSR[ 20 ][ 365 ],
   alphaCSR[ 20 ][ 366 ],
   alphaCSR[ 20 ][ 367 ],
   alphaCSR[ 20 ][ 368 ],
   alphaCSR[ 20 ][ 369 ],
   alphaCSR[ 20 ][ 370 ],
   alphaCSR[ 20 ][ 371 ],
   alphaCSR[ 20 ][ 372 ],
   alphaCSR[ 20 ][ 373 ],
   alphaCSR[ 20 ][ 374 ],
   alphaCSR[ 20 ][ 375 ],
   alphaCSR[ 20 ][ 376 ],
   alphaCSR[ 20 ][ 377 ],
   alphaCSR[ 20 ][ 378 ],
   alphaCSR[ 20 ][ 379 ],
   alphaCSR[ 20 ][ 380 ],
   alphaCSR[ 20 ][ 381 ],
   alphaCSR[ 20 ][ 382 ],
   alphaCSR[ 20 ][ 383 ],
   alphaCSR[ 21 ][ 0 ],
   alphaCSR[ 21 ][ 1 ],
   alphaCSR[ 21 ][ 2 ],
   alphaCSR[ 21 ][ 3 ],
   alphaCSR[ 21 ][ 4 ],
   alphaCSR[ 21 ][ 5 ],
   alphaCSR[ 21 ][ 6 ],
   alphaCSR[ 21 ][ 7 ],
   alphaCSR[ 21 ][ 8 ],
   alphaCSR[ 21 ][ 9 ],
   alphaCSR[ 21 ][ 10 ],
   alphaCSR[ 21 ][ 11 ],
   alphaCSR[ 21 ][ 12 ],
   alphaCSR[ 21 ][ 13 ],
   alphaCSR[ 21 ][ 14 ],
   alphaCSR[ 21 ][ 15 ],
   alphaCSR[ 21 ][ 16 ],
   alphaCSR[ 21 ][ 17 ],
   alphaCSR[ 21 ][ 18 ],
   alphaCSR[ 21 ][ 19 ],
   alphaCSR[ 21 ][ 20 ],
   alphaCSR[ 21 ][ 21 ],
   alphaCSR[ 21 ][ 22 ],
   alphaCSR[ 21 ][ 23 ],
   alphaCSR[ 21 ][ 24 ],
   alphaCSR[ 21 ][ 25 ],
   alphaCSR[ 21 ][ 26 ],
   alphaCSR[ 21 ][ 27 ],
   alphaCSR[ 21 ][ 28 ],
   alphaCSR[ 21 ][ 29 ],
   alphaCSR[ 21 ][ 30 ],
   alphaCSR[ 21 ][ 31 ],
   alphaCSR[ 21 ][ 32 ],
   alphaCSR[ 21 ][ 33 ],
   alphaCSR[ 21 ][ 34 ],
   alphaCSR[ 21 ][ 35 ],
   alphaCSR[ 21 ][ 36 ],
   alphaCSR[ 21 ][ 37 ],
   alphaCSR[ 21 ][ 38 ],
   alphaCSR[ 21 ][ 39 ],
   alphaCSR[ 21 ][ 40 ],
   alphaCSR[ 21 ][ 41 ],
   alphaCSR[ 21 ][ 42 ],
   alphaCSR[ 21 ][ 43 ],
   alphaCSR[ 21 ][ 44 ],
   alphaCSR[ 21 ][ 45 ],
   alphaCSR[ 21 ][ 46 ],
   alphaCSR[ 21 ][ 47 ],
   alphaCSR[ 21 ][ 48 ],
   alphaCSR[ 21 ][ 49 ],
   alphaCSR[ 21 ][ 50 ],
   alphaCSR[ 21 ][ 51 ],
   alphaCSR[ 21 ][ 52 ],
   alphaCSR[ 21 ][ 53 ],
   alphaCSR[ 21 ][ 54 ],
   alphaCSR[ 21 ][ 55 ],
   alphaCSR[ 21 ][ 56 ],
   alphaCSR[ 21 ][ 57 ],
   alphaCSR[ 21 ][ 58 ],
   alphaCSR[ 21 ][ 59 ],
   alphaCSR[ 21 ][ 60 ],
   alphaCSR[ 21 ][ 61 ],
   alphaCSR[ 21 ][ 62 ],
   alphaCSR[ 21 ][ 63 ],
   alphaCSR[ 21 ][ 64 ],
   alphaCSR[ 21 ][ 65 ],
   alphaCSR[ 21 ][ 66 ],
   alphaCSR[ 21 ][ 67 ],
   alphaCSR[ 21 ][ 68 ],
   alphaCSR[ 21 ][ 69 ],
   alphaCSR[ 21 ][ 70 ],
   alphaCSR[ 21 ][ 71 ],
   alphaCSR[ 21 ][ 72 ],
   alphaCSR[ 21 ][ 73 ],
   alphaCSR[ 21 ][ 74 ],
   alphaCSR[ 21 ][ 75 ],
   alphaCSR[ 21 ][ 76 ],
   alphaCSR[ 21 ][ 77 ],
   alphaCSR[ 21 ][ 78 ],
   alphaCSR[ 21 ][ 79 ],
   alphaCSR[ 21 ][ 80 ],
   alphaCSR[ 21 ][ 81 ],
   alphaCSR[ 21 ][ 82 ],
   alphaCSR[ 21 ][ 83 ],
   alphaCSR[ 21 ][ 84 ],
   alphaCSR[ 21 ][ 85 ],
   alphaCSR[ 21 ][ 86 ],
   alphaCSR[ 21 ][ 87 ],
   alphaCSR[ 21 ][ 88 ],
   alphaCSR[ 21 ][ 89 ],
   alphaCSR[ 21 ][ 90 ],
   alphaCSR[ 21 ][ 91 ],
   alphaCSR[ 21 ][ 92 ],
   alphaCSR[ 21 ][ 93 ],
   alphaCSR[ 21 ][ 94 ],
   alphaCSR[ 21 ][ 95 ],
   alphaCSR[ 21 ][ 96 ],
   alphaCSR[ 21 ][ 97 ],
   alphaCSR[ 21 ][ 98 ],
   alphaCSR[ 21 ][ 99 ],
   alphaCSR[ 21 ][ 100 ],
   alphaCSR[ 21 ][ 101 ],
   alphaCSR[ 21 ][ 102 ],
   alphaCSR[ 21 ][ 103 ],
   alphaCSR[ 21 ][ 104 ],
   alphaCSR[ 21 ][ 105 ],
   alphaCSR[ 21 ][ 106 ],
   alphaCSR[ 21 ][ 107 ],
   alphaCSR[ 21 ][ 108 ],
   alphaCSR[ 21 ][ 109 ],
   alphaCSR[ 21 ][ 110 ],
   alphaCSR[ 21 ][ 111 ],
   alphaCSR[ 21 ][ 112 ],
   alphaCSR[ 21 ][ 113 ],
   alphaCSR[ 21 ][ 114 ],
   alphaCSR[ 21 ][ 115 ],
   alphaCSR[ 21 ][ 116 ],
   alphaCSR[ 21 ][ 117 ],
   alphaCSR[ 21 ][ 118 ],
   alphaCSR[ 21 ][ 119 ],
   alphaCSR[ 21 ][ 120 ],
   alphaCSR[ 21 ][ 121 ],
   alphaCSR[ 21 ][ 122 ],
   alphaCSR[ 21 ][ 123 ],
   alphaCSR[ 21 ][ 124 ],
   alphaCSR[ 21 ][ 125 ],
   alphaCSR[ 21 ][ 126 ],
   alphaCSR[ 21 ][ 127 ],
   alphaCSR[ 21 ][ 128 ],
   alphaCSR[ 21 ][ 129 ],
   alphaCSR[ 21 ][ 130 ],
   alphaCSR[ 21 ][ 131 ],
   alphaCSR[ 21 ][ 132 ],
   alphaCSR[ 21 ][ 133 ],
   alphaCSR[ 21 ][ 134 ],
   alphaCSR[ 21 ][ 135 ],
   alphaCSR[ 21 ][ 136 ],
   alphaCSR[ 21 ][ 137 ],
   alphaCSR[ 21 ][ 138 ],
   alphaCSR[ 21 ][ 139 ],
   alphaCSR[ 21 ][ 140 ],
   alphaCSR[ 21 ][ 141 ],
   alphaCSR[ 21 ][ 142 ],
   alphaCSR[ 21 ][ 143 ],
   alphaCSR[ 21 ][ 144 ],
   alphaCSR[ 21 ][ 145 ],
   alphaCSR[ 21 ][ 146 ],
   alphaCSR[ 21 ][ 147 ],
   alphaCSR[ 21 ][ 148 ],
   alphaCSR[ 21 ][ 149 ],
   alphaCSR[ 21 ][ 150 ],
   alphaCSR[ 21 ][ 151 ],
   alphaCSR[ 21 ][ 152 ],
   alphaCSR[ 21 ][ 153 ],
   alphaCSR[ 21 ][ 154 ],
   alphaCSR[ 21 ][ 155 ],
   alphaCSR[ 21 ][ 156 ],
   alphaCSR[ 21 ][ 157 ],
   alphaCSR[ 21 ][ 158 ],
   alphaCSR[ 21 ][ 159 ],
   alphaCSR[ 21 ][ 160 ],
   alphaCSR[ 21 ][ 161 ],
   alphaCSR[ 21 ][ 162 ],
   alphaCSR[ 21 ][ 163 ],
   alphaCSR[ 21 ][ 164 ],
   alphaCSR[ 21 ][ 165 ],
   alphaCSR[ 21 ][ 166 ],
   alphaCSR[ 21 ][ 167 ],
   alphaCSR[ 21 ][ 168 ],
   alphaCSR[ 21 ][ 169 ],
   alphaCSR[ 21 ][ 170 ],
   alphaCSR[ 21 ][ 171 ],
   alphaCSR[ 21 ][ 172 ],
   alphaCSR[ 21 ][ 173 ],
   alphaCSR[ 21 ][ 174 ],
   alphaCSR[ 21 ][ 175 ],
   alphaCSR[ 21 ][ 176 ],
   alphaCSR[ 21 ][ 177 ],
   alphaCSR[ 21 ][ 178 ],
   alphaCSR[ 21 ][ 179 ],
   alphaCSR[ 21 ][ 180 ],
   alphaCSR[ 21 ][ 181 ],
   alphaCSR[ 21 ][ 182 ],
   alphaCSR[ 21 ][ 183 ],
   alphaCSR[ 21 ][ 184 ],
   alphaCSR[ 21 ][ 185 ],
   alphaCSR[ 21 ][ 186 ],
   alphaCSR[ 21 ][ 187 ],
   alphaCSR[ 21 ][ 188 ],
   alphaCSR[ 21 ][ 189 ],
   alphaCSR[ 21 ][ 190 ],
   alphaCSR[ 21 ][ 191 ],
   alphaCSR[ 21 ][ 192 ],
   alphaCSR[ 21 ][ 193 ],
   alphaCSR[ 21 ][ 194 ],
   alphaCSR[ 21 ][ 195 ],
   alphaCSR[ 21 ][ 196 ],
   alphaCSR[ 21 ][ 197 ],
   alphaCSR[ 21 ][ 198 ],
   alphaCSR[ 21 ][ 199 ],
   alphaCSR[ 21 ][ 200 ],
   alphaCSR[ 21 ][ 201 ],
   alphaCSR[ 21 ][ 202 ],
   alphaCSR[ 21 ][ 203 ],
   alphaCSR[ 21 ][ 204 ],
   alphaCSR[ 21 ][ 205 ],
   alphaCSR[ 21 ][ 206 ],
   alphaCSR[ 21 ][ 207 ],
   alphaCSR[ 21 ][ 208 ],
   alphaCSR[ 21 ][ 209 ],
   alphaCSR[ 21 ][ 210 ],
   alphaCSR[ 21 ][ 211 ],
   alphaCSR[ 21 ][ 212 ],
   alphaCSR[ 21 ][ 213 ],
   alphaCSR[ 21 ][ 214 ],
   alphaCSR[ 21 ][ 215 ],
   alphaCSR[ 21 ][ 216 ],
   alphaCSR[ 21 ][ 217 ],
   alphaCSR[ 21 ][ 218 ],
   alphaCSR[ 21 ][ 219 ],
   alphaCSR[ 21 ][ 220 ],
   alphaCSR[ 21 ][ 221 ],
   alphaCSR[ 21 ][ 222 ],
   alphaCSR[ 21 ][ 223 ],
   alphaCSR[ 21 ][ 224 ],
   alphaCSR[ 21 ][ 225 ],
   alphaCSR[ 21 ][ 226 ],
   alphaCSR[ 21 ][ 227 ],
   alphaCSR[ 21 ][ 228 ],
   alphaCSR[ 21 ][ 229 ],
   alphaCSR[ 21 ][ 230 ],
   alphaCSR[ 21 ][ 231 ],
   alphaCSR[ 21 ][ 232 ],
   alphaCSR[ 21 ][ 233 ],
   alphaCSR[ 21 ][ 234 ],
   alphaCSR[ 21 ][ 235 ],
   alphaCSR[ 21 ][ 236 ],
   alphaCSR[ 21 ][ 237 ],
   alphaCSR[ 21 ][ 238 ],
   alphaCSR[ 21 ][ 239 ],
   alphaCSR[ 21 ][ 240 ],
   alphaCSR[ 21 ][ 241 ],
   alphaCSR[ 21 ][ 242 ],
   alphaCSR[ 21 ][ 243 ],
   alphaCSR[ 21 ][ 244 ],
   alphaCSR[ 21 ][ 245 ],
   alphaCSR[ 21 ][ 246 ],
   alphaCSR[ 21 ][ 247 ],
   alphaCSR[ 21 ][ 248 ],
   alphaCSR[ 21 ][ 249 ],
   alphaCSR[ 21 ][ 250 ],
   alphaCSR[ 21 ][ 251 ],
   alphaCSR[ 21 ][ 252 ],
   alphaCSR[ 21 ][ 253 ],
   alphaCSR[ 21 ][ 254 ],
   alphaCSR[ 21 ][ 255 ],
   alphaCSR[ 21 ][ 256 ],
   alphaCSR[ 21 ][ 257 ],
   alphaCSR[ 21 ][ 258 ],
   alphaCSR[ 21 ][ 259 ],
   alphaCSR[ 21 ][ 260 ],
   alphaCSR[ 21 ][ 261 ],
   alphaCSR[ 21 ][ 262 ],
   alphaCSR[ 21 ][ 263 ],
   alphaCSR[ 21 ][ 264 ],
   alphaCSR[ 21 ][ 265 ],
   alphaCSR[ 21 ][ 266 ],
   alphaCSR[ 21 ][ 267 ],
   alphaCSR[ 21 ][ 268 ],
   alphaCSR[ 21 ][ 269 ],
   alphaCSR[ 21 ][ 270 ],
   alphaCSR[ 21 ][ 271 ],
   alphaCSR[ 21 ][ 272 ],
   alphaCSR[ 21 ][ 273 ],
   alphaCSR[ 21 ][ 274 ],
   alphaCSR[ 21 ][ 275 ],
   alphaCSR[ 21 ][ 276 ],
   alphaCSR[ 21 ][ 277 ],
   alphaCSR[ 21 ][ 278 ],
   alphaCSR[ 21 ][ 279 ],
   alphaCSR[ 21 ][ 280 ],
   alphaCSR[ 21 ][ 281 ],
   alphaCSR[ 21 ][ 282 ],
   alphaCSR[ 21 ][ 283 ],
   alphaCSR[ 21 ][ 284 ],
   alphaCSR[ 21 ][ 285 ],
   alphaCSR[ 21 ][ 286 ],
   alphaCSR[ 21 ][ 287 ],
   alphaCSR[ 21 ][ 288 ],
   alphaCSR[ 21 ][ 289 ],
   alphaCSR[ 21 ][ 290 ],
   alphaCSR[ 21 ][ 291 ],
   alphaCSR[ 21 ][ 292 ],
   alphaCSR[ 21 ][ 293 ],
   alphaCSR[ 21 ][ 294 ],
   alphaCSR[ 21 ][ 295 ],
   alphaCSR[ 21 ][ 296 ],
   alphaCSR[ 21 ][ 297 ],
   alphaCSR[ 21 ][ 298 ],
   alphaCSR[ 21 ][ 299 ],
   alphaCSR[ 21 ][ 300 ],
   alphaCSR[ 21 ][ 301 ],
   alphaCSR[ 21 ][ 302 ],
   alphaCSR[ 21 ][ 303 ],
   alphaCSR[ 21 ][ 304 ],
   alphaCSR[ 21 ][ 305 ],
   alphaCSR[ 21 ][ 306 ],
   alphaCSR[ 21 ][ 307 ],
   alphaCSR[ 21 ][ 308 ],
   alphaCSR[ 21 ][ 309 ],
   alphaCSR[ 21 ][ 310 ],
   alphaCSR[ 21 ][ 311 ],
   alphaCSR[ 21 ][ 312 ],
   alphaCSR[ 21 ][ 313 ],
   alphaCSR[ 21 ][ 314 ],
   alphaCSR[ 21 ][ 315 ],
   alphaCSR[ 21 ][ 316 ],
   alphaCSR[ 21 ][ 317 ],
   alphaCSR[ 21 ][ 318 ],
   alphaCSR[ 21 ][ 319 ],
   alphaCSR[ 21 ][ 320 ],
   alphaCSR[ 21 ][ 321 ],
   alphaCSR[ 21 ][ 322 ],
   alphaCSR[ 21 ][ 323 ],
   alphaCSR[ 21 ][ 324 ],
   alphaCSR[ 21 ][ 325 ],
   alphaCSR[ 21 ][ 326 ],
   alphaCSR[ 21 ][ 327 ],
   alphaCSR[ 21 ][ 328 ],
   alphaCSR[ 21 ][ 329 ],
   alphaCSR[ 21 ][ 330 ],
   alphaCSR[ 21 ][ 331 ],
   alphaCSR[ 21 ][ 332 ],
   alphaCSR[ 21 ][ 333 ],
   alphaCSR[ 21 ][ 334 ],
   alphaCSR[ 21 ][ 335 ],
   alphaCSR[ 21 ][ 336 ],
   alphaCSR[ 21 ][ 337 ],
   alphaCSR[ 21 ][ 338 ],
   alphaCSR[ 21 ][ 339 ],
   alphaCSR[ 21 ][ 340 ],
   alphaCSR[ 21 ][ 341 ],
   alphaCSR[ 21 ][ 342 ],
   alphaCSR[ 21 ][ 343 ],
   alphaCSR[ 21 ][ 344 ],
   alphaCSR[ 21 ][ 345 ],
   alphaCSR[ 21 ][ 346 ],
   alphaCSR[ 21 ][ 347 ],
   alphaCSR[ 21 ][ 348 ],
   alphaCSR[ 21 ][ 349 ],
   alphaCSR[ 21 ][ 350 ],
   alphaCSR[ 21 ][ 351 ],
   alphaCSR[ 21 ][ 352 ],
   alphaCSR[ 21 ][ 353 ],
   alphaCSR[ 21 ][ 354 ],
   alphaCSR[ 21 ][ 355 ],
   alphaCSR[ 21 ][ 356 ],
   alphaCSR[ 21 ][ 357 ],
   alphaCSR[ 21 ][ 358 ],
   alphaCSR[ 21 ][ 359 ],
   alphaCSR[ 21 ][ 360 ],
   alphaCSR[ 21 ][ 361 ],
   alphaCSR[ 21 ][ 362 ],
   alphaCSR[ 21 ][ 363 ],
   alphaCSR[ 21 ][ 364 ],
   alphaCSR[ 21 ][ 365 ],
   alphaCSR[ 21 ][ 366 ],
   alphaCSR[ 21 ][ 367 ],
   alphaCSR[ 21 ][ 368 ],
   alphaCSR[ 21 ][ 369 ],
   alphaCSR[ 21 ][ 370 ],
   alphaCSR[ 21 ][ 371 ],
   alphaCSR[ 21 ][ 372 ],
   alphaCSR[ 21 ][ 373 ],
   alphaCSR[ 21 ][ 374 ],
   alphaCSR[ 21 ][ 375 ],
   alphaCSR[ 21 ][ 376 ],
   alphaCSR[ 21 ][ 377 ],
   alphaCSR[ 21 ][ 378 ],
   alphaCSR[ 21 ][ 379 ],
   alphaCSR[ 21 ][ 380 ],
   alphaCSR[ 21 ][ 381 ],
   alphaCSR[ 21 ][ 382 ],
   alphaCSR[ 21 ][ 383 ],
   alphaCSR[ 22 ][ 0 ],
   alphaCSR[ 22 ][ 1 ],
   alphaCSR[ 22 ][ 2 ],
   alphaCSR[ 22 ][ 3 ],
   alphaCSR[ 22 ][ 4 ],
   alphaCSR[ 22 ][ 5 ],
   alphaCSR[ 22 ][ 6 ],
   alphaCSR[ 22 ][ 7 ],
   alphaCSR[ 22 ][ 8 ],
   alphaCSR[ 22 ][ 9 ],
   alphaCSR[ 22 ][ 10 ],
   alphaCSR[ 22 ][ 11 ],
   alphaCSR[ 22 ][ 12 ],
   alphaCSR[ 22 ][ 13 ],
   alphaCSR[ 22 ][ 14 ],
   alphaCSR[ 22 ][ 15 ],
   alphaCSR[ 22 ][ 16 ],
   alphaCSR[ 22 ][ 17 ],
   alphaCSR[ 22 ][ 18 ],
   alphaCSR[ 22 ][ 19 ],
   alphaCSR[ 22 ][ 20 ],
   alphaCSR[ 22 ][ 21 ],
   alphaCSR[ 22 ][ 22 ],
   alphaCSR[ 22 ][ 23 ],
   alphaCSR[ 22 ][ 24 ],
   alphaCSR[ 22 ][ 25 ],
   alphaCSR[ 22 ][ 26 ],
   alphaCSR[ 22 ][ 27 ],
   alphaCSR[ 22 ][ 28 ],
   alphaCSR[ 22 ][ 29 ],
   alphaCSR[ 22 ][ 30 ],
   alphaCSR[ 22 ][ 31 ],
   alphaCSR[ 22 ][ 32 ],
   alphaCSR[ 22 ][ 33 ],
   alphaCSR[ 22 ][ 34 ],
   alphaCSR[ 22 ][ 35 ],
   alphaCSR[ 22 ][ 36 ],
   alphaCSR[ 22 ][ 37 ],
   alphaCSR[ 22 ][ 38 ],
   alphaCSR[ 22 ][ 39 ],
   alphaCSR[ 22 ][ 40 ],
   alphaCSR[ 22 ][ 41 ],
   alphaCSR[ 22 ][ 42 ],
   alphaCSR[ 22 ][ 43 ],
   alphaCSR[ 22 ][ 44 ],
   alphaCSR[ 22 ][ 45 ],
   alphaCSR[ 22 ][ 46 ],
   alphaCSR[ 22 ][ 47 ],
   alphaCSR[ 22 ][ 48 ],
   alphaCSR[ 22 ][ 49 ],
   alphaCSR[ 22 ][ 50 ],
   alphaCSR[ 22 ][ 51 ],
   alphaCSR[ 22 ][ 52 ],
   alphaCSR[ 22 ][ 53 ],
   alphaCSR[ 22 ][ 54 ],
   alphaCSR[ 22 ][ 55 ],
   alphaCSR[ 22 ][ 56 ],
   alphaCSR[ 22 ][ 57 ],
   alphaCSR[ 22 ][ 58 ],
   alphaCSR[ 22 ][ 59 ],
   alphaCSR[ 22 ][ 60 ],
   alphaCSR[ 22 ][ 61 ],
   alphaCSR[ 22 ][ 62 ],
   alphaCSR[ 22 ][ 63 ],
   alphaCSR[ 22 ][ 64 ],
   alphaCSR[ 22 ][ 65 ],
   alphaCSR[ 22 ][ 66 ],
   alphaCSR[ 22 ][ 67 ],
   alphaCSR[ 22 ][ 68 ],
   alphaCSR[ 22 ][ 69 ],
   alphaCSR[ 22 ][ 70 ],
   alphaCSR[ 22 ][ 71 ],
   alphaCSR[ 22 ][ 72 ],
   alphaCSR[ 22 ][ 73 ],
   alphaCSR[ 22 ][ 74 ],
   alphaCSR[ 22 ][ 75 ],
   alphaCSR[ 22 ][ 76 ],
   alphaCSR[ 22 ][ 77 ],
   alphaCSR[ 22 ][ 78 ],
   alphaCSR[ 22 ][ 79 ],
   alphaCSR[ 22 ][ 80 ],
   alphaCSR[ 22 ][ 81 ],
   alphaCSR[ 22 ][ 82 ],
   alphaCSR[ 22 ][ 83 ],
   alphaCSR[ 22 ][ 84 ],
   alphaCSR[ 22 ][ 85 ],
   alphaCSR[ 22 ][ 86 ],
   alphaCSR[ 22 ][ 87 ],
   alphaCSR[ 22 ][ 88 ],
   alphaCSR[ 22 ][ 89 ],
   alphaCSR[ 22 ][ 90 ],
   alphaCSR[ 22 ][ 91 ],
   alphaCSR[ 22 ][ 92 ],
   alphaCSR[ 22 ][ 93 ],
   alphaCSR[ 22 ][ 94 ],
   alphaCSR[ 22 ][ 95 ],
   alphaCSR[ 22 ][ 96 ],
   alphaCSR[ 22 ][ 97 ],
   alphaCSR[ 22 ][ 98 ],
   alphaCSR[ 22 ][ 99 ],
   alphaCSR[ 22 ][ 100 ],
   alphaCSR[ 22 ][ 101 ],
   alphaCSR[ 22 ][ 102 ],
   alphaCSR[ 22 ][ 103 ],
   alphaCSR[ 22 ][ 104 ],
   alphaCSR[ 22 ][ 105 ],
   alphaCSR[ 22 ][ 106 ],
   alphaCSR[ 22 ][ 107 ],
   alphaCSR[ 22 ][ 108 ],
   alphaCSR[ 22 ][ 109 ],
   alphaCSR[ 22 ][ 110 ],
   alphaCSR[ 22 ][ 111 ],
   alphaCSR[ 22 ][ 112 ],
   alphaCSR[ 22 ][ 113 ],
   alphaCSR[ 22 ][ 114 ],
   alphaCSR[ 22 ][ 115 ],
   alphaCSR[ 22 ][ 116 ],
   alphaCSR[ 22 ][ 117 ],
   alphaCSR[ 22 ][ 118 ],
   alphaCSR[ 22 ][ 119 ],
   alphaCSR[ 22 ][ 120 ],
   alphaCSR[ 22 ][ 121 ],
   alphaCSR[ 22 ][ 122 ],
   alphaCSR[ 22 ][ 123 ],
   alphaCSR[ 22 ][ 124 ],
   alphaCSR[ 22 ][ 125 ],
   alphaCSR[ 22 ][ 126 ],
   alphaCSR[ 22 ][ 127 ],
   alphaCSR[ 22 ][ 128 ],
   alphaCSR[ 22 ][ 129 ],
   alphaCSR[ 22 ][ 130 ],
   alphaCSR[ 22 ][ 131 ],
   alphaCSR[ 22 ][ 132 ],
   alphaCSR[ 22 ][ 133 ],
   alphaCSR[ 22 ][ 134 ],
   alphaCSR[ 22 ][ 135 ],
   alphaCSR[ 22 ][ 136 ],
   alphaCSR[ 22 ][ 137 ],
   alphaCSR[ 22 ][ 138 ],
   alphaCSR[ 22 ][ 139 ],
   alphaCSR[ 22 ][ 140 ],
   alphaCSR[ 22 ][ 141 ],
   alphaCSR[ 22 ][ 142 ],
   alphaCSR[ 22 ][ 143 ],
   alphaCSR[ 22 ][ 144 ],
   alphaCSR[ 22 ][ 145 ],
   alphaCSR[ 22 ][ 146 ],
   alphaCSR[ 22 ][ 147 ],
   alphaCSR[ 22 ][ 148 ],
   alphaCSR[ 22 ][ 149 ],
   alphaCSR[ 22 ][ 150 ],
   alphaCSR[ 22 ][ 151 ],
   alphaCSR[ 22 ][ 152 ],
   alphaCSR[ 22 ][ 153 ],
   alphaCSR[ 22 ][ 154 ],
   alphaCSR[ 22 ][ 155 ],
   alphaCSR[ 22 ][ 156 ],
   alphaCSR[ 22 ][ 157 ],
   alphaCSR[ 22 ][ 158 ],
   alphaCSR[ 22 ][ 159 ],
   alphaCSR[ 22 ][ 160 ],
   alphaCSR[ 22 ][ 161 ],
   alphaCSR[ 22 ][ 162 ],
   alphaCSR[ 22 ][ 163 ],
   alphaCSR[ 22 ][ 164 ],
   alphaCSR[ 22 ][ 165 ],
   alphaCSR[ 22 ][ 166 ],
   alphaCSR[ 22 ][ 167 ],
   alphaCSR[ 22 ][ 168 ],
   alphaCSR[ 22 ][ 169 ],
   alphaCSR[ 22 ][ 170 ],
   alphaCSR[ 22 ][ 171 ],
   alphaCSR[ 22 ][ 172 ],
   alphaCSR[ 22 ][ 173 ],
   alphaCSR[ 22 ][ 174 ],
   alphaCSR[ 22 ][ 175 ],
   alphaCSR[ 22 ][ 176 ],
   alphaCSR[ 22 ][ 177 ],
   alphaCSR[ 22 ][ 178 ],
   alphaCSR[ 22 ][ 179 ],
   alphaCSR[ 22 ][ 180 ],
   alphaCSR[ 22 ][ 181 ],
   alphaCSR[ 22 ][ 182 ],
   alphaCSR[ 22 ][ 183 ],
   alphaCSR[ 22 ][ 184 ],
   alphaCSR[ 22 ][ 185 ],
   alphaCSR[ 22 ][ 186 ],
   alphaCSR[ 22 ][ 187 ],
   alphaCSR[ 22 ][ 188 ],
   alphaCSR[ 22 ][ 189 ],
   alphaCSR[ 22 ][ 190 ],
   alphaCSR[ 22 ][ 191 ],
   alphaCSR[ 22 ][ 192 ],
   alphaCSR[ 22 ][ 193 ],
   alphaCSR[ 22 ][ 194 ],
   alphaCSR[ 22 ][ 195 ],
   alphaCSR[ 22 ][ 196 ],
   alphaCSR[ 22 ][ 197 ],
   alphaCSR[ 22 ][ 198 ],
   alphaCSR[ 22 ][ 199 ],
   alphaCSR[ 22 ][ 200 ],
   alphaCSR[ 22 ][ 201 ],
   alphaCSR[ 22 ][ 202 ],
   alphaCSR[ 22 ][ 203 ],
   alphaCSR[ 22 ][ 204 ],
   alphaCSR[ 22 ][ 205 ],
   alphaCSR[ 22 ][ 206 ],
   alphaCSR[ 22 ][ 207 ],
   alphaCSR[ 22 ][ 208 ],
   alphaCSR[ 22 ][ 209 ],
   alphaCSR[ 22 ][ 210 ],
   alphaCSR[ 22 ][ 211 ],
   alphaCSR[ 22 ][ 212 ],
   alphaCSR[ 22 ][ 213 ],
   alphaCSR[ 22 ][ 214 ],
   alphaCSR[ 22 ][ 215 ],
   alphaCSR[ 22 ][ 216 ],
   alphaCSR[ 22 ][ 217 ],
   alphaCSR[ 22 ][ 218 ],
   alphaCSR[ 22 ][ 219 ],
   alphaCSR[ 22 ][ 220 ],
   alphaCSR[ 22 ][ 221 ],
   alphaCSR[ 22 ][ 222 ],
   alphaCSR[ 22 ][ 223 ],
   alphaCSR[ 22 ][ 224 ],
   alphaCSR[ 22 ][ 225 ],
   alphaCSR[ 22 ][ 226 ],
   alphaCSR[ 22 ][ 227 ],
   alphaCSR[ 22 ][ 228 ],
   alphaCSR[ 22 ][ 229 ],
   alphaCSR[ 22 ][ 230 ],
   alphaCSR[ 22 ][ 231 ],
   alphaCSR[ 22 ][ 232 ],
   alphaCSR[ 22 ][ 233 ],
   alphaCSR[ 22 ][ 234 ],
   alphaCSR[ 22 ][ 235 ],
   alphaCSR[ 22 ][ 236 ],
   alphaCSR[ 22 ][ 237 ],
   alphaCSR[ 22 ][ 238 ],
   alphaCSR[ 22 ][ 239 ],
   alphaCSR[ 22 ][ 240 ],
   alphaCSR[ 22 ][ 241 ],
   alphaCSR[ 22 ][ 242 ],
   alphaCSR[ 22 ][ 243 ],
   alphaCSR[ 22 ][ 244 ],
   alphaCSR[ 22 ][ 245 ],
   alphaCSR[ 22 ][ 246 ],
   alphaCSR[ 22 ][ 247 ],
   alphaCSR[ 22 ][ 248 ],
   alphaCSR[ 22 ][ 249 ],
   alphaCSR[ 22 ][ 250 ],
   alphaCSR[ 22 ][ 251 ],
   alphaCSR[ 22 ][ 252 ],
   alphaCSR[ 22 ][ 253 ],
   alphaCSR[ 22 ][ 254 ],
   alphaCSR[ 22 ][ 255 ],
   alphaCSR[ 22 ][ 256 ],
   alphaCSR[ 22 ][ 257 ],
   alphaCSR[ 22 ][ 258 ],
   alphaCSR[ 22 ][ 259 ],
   alphaCSR[ 22 ][ 260 ],
   alphaCSR[ 22 ][ 261 ],
   alphaCSR[ 22 ][ 262 ],
   alphaCSR[ 22 ][ 263 ],
   alphaCSR[ 22 ][ 264 ],
   alphaCSR[ 22 ][ 265 ],
   alphaCSR[ 22 ][ 266 ],
   alphaCSR[ 22 ][ 267 ],
   alphaCSR[ 22 ][ 268 ],
   alphaCSR[ 22 ][ 269 ],
   alphaCSR[ 22 ][ 270 ],
   alphaCSR[ 22 ][ 271 ],
   alphaCSR[ 22 ][ 272 ],
   alphaCSR[ 22 ][ 273 ],
   alphaCSR[ 22 ][ 274 ],
   alphaCSR[ 22 ][ 275 ],
   alphaCSR[ 22 ][ 276 ],
   alphaCSR[ 22 ][ 277 ],
   alphaCSR[ 22 ][ 278 ],
   alphaCSR[ 22 ][ 279 ],
   alphaCSR[ 22 ][ 280 ],
   alphaCSR[ 22 ][ 281 ],
   alphaCSR[ 22 ][ 282 ],
   alphaCSR[ 22 ][ 283 ],
   alphaCSR[ 22 ][ 284 ],
   alphaCSR[ 22 ][ 285 ],
   alphaCSR[ 22 ][ 286 ],
   alphaCSR[ 22 ][ 287 ],
   alphaCSR[ 22 ][ 288 ],
   alphaCSR[ 22 ][ 289 ],
   alphaCSR[ 22 ][ 290 ],
   alphaCSR[ 22 ][ 291 ],
   alphaCSR[ 22 ][ 292 ],
   alphaCSR[ 22 ][ 293 ],
   alphaCSR[ 22 ][ 294 ],
   alphaCSR[ 22 ][ 295 ],
   alphaCSR[ 22 ][ 296 ],
   alphaCSR[ 22 ][ 297 ],
   alphaCSR[ 22 ][ 298 ],
   alphaCSR[ 22 ][ 299 ],
   alphaCSR[ 22 ][ 300 ],
   alphaCSR[ 22 ][ 301 ],
   alphaCSR[ 22 ][ 302 ],
   alphaCSR[ 22 ][ 303 ],
   alphaCSR[ 22 ][ 304 ],
   alphaCSR[ 22 ][ 305 ],
   alphaCSR[ 22 ][ 306 ],
   alphaCSR[ 22 ][ 307 ],
   alphaCSR[ 22 ][ 308 ],
   alphaCSR[ 22 ][ 309 ],
   alphaCSR[ 22 ][ 310 ],
   alphaCSR[ 22 ][ 311 ],
   alphaCSR[ 22 ][ 312 ],
   alphaCSR[ 22 ][ 313 ],
   alphaCSR[ 22 ][ 314 ],
   alphaCSR[ 22 ][ 315 ],
   alphaCSR[ 22 ][ 316 ],
   alphaCSR[ 22 ][ 317 ],
   alphaCSR[ 22 ][ 318 ],
   alphaCSR[ 22 ][ 319 ],
   alphaCSR[ 22 ][ 320 ],
   alphaCSR[ 22 ][ 321 ],
   alphaCSR[ 22 ][ 322 ],
   alphaCSR[ 22 ][ 323 ],
   alphaCSR[ 22 ][ 324 ],
   alphaCSR[ 22 ][ 325 ],
   alphaCSR[ 22 ][ 326 ],
   alphaCSR[ 22 ][ 327 ],
   alphaCSR[ 22 ][ 328 ],
   alphaCSR[ 22 ][ 329 ],
   alphaCSR[ 22 ][ 330 ],
   alphaCSR[ 22 ][ 331 ],
   alphaCSR[ 22 ][ 332 ],
   alphaCSR[ 22 ][ 333 ],
   alphaCSR[ 22 ][ 334 ],
   alphaCSR[ 22 ][ 335 ],
   alphaCSR[ 22 ][ 336 ],
   alphaCSR[ 22 ][ 337 ],
   alphaCSR[ 22 ][ 338 ],
   alphaCSR[ 22 ][ 339 ],
   alphaCSR[ 22 ][ 340 ],
   alphaCSR[ 22 ][ 341 ],
   alphaCSR[ 22 ][ 342 ],
   alphaCSR[ 22 ][ 343 ],
   alphaCSR[ 22 ][ 344 ],
   alphaCSR[ 22 ][ 345 ],
   alphaCSR[ 22 ][ 346 ],
   alphaCSR[ 22 ][ 347 ],
   alphaCSR[ 22 ][ 348 ],
   alphaCSR[ 22 ][ 349 ],
   alphaCSR[ 22 ][ 350 ],
   alphaCSR[ 22 ][ 351 ],
   alphaCSR[ 22 ][ 352 ],
   alphaCSR[ 22 ][ 353 ],
   alphaCSR[ 22 ][ 354 ],
   alphaCSR[ 22 ][ 355 ],
   alphaCSR[ 22 ][ 356 ],
   alphaCSR[ 22 ][ 357 ],
   alphaCSR[ 22 ][ 358 ],
   alphaCSR[ 22 ][ 359 ],
   alphaCSR[ 22 ][ 360 ],
   alphaCSR[ 22 ][ 361 ],
   alphaCSR[ 22 ][ 362 ],
   alphaCSR[ 22 ][ 363 ],
   alphaCSR[ 22 ][ 364 ],
   alphaCSR[ 22 ][ 365 ],
   alphaCSR[ 22 ][ 366 ],
   alphaCSR[ 22 ][ 367 ],
   alphaCSR[ 22 ][ 368 ],
   alphaCSR[ 22 ][ 369 ],
   alphaCSR[ 22 ][ 370 ],
   alphaCSR[ 22 ][ 371 ],
   alphaCSR[ 22 ][ 372 ],
   alphaCSR[ 22 ][ 373 ],
   alphaCSR[ 22 ][ 374 ],
   alphaCSR[ 22 ][ 375 ],
   alphaCSR[ 22 ][ 376 ],
   alphaCSR[ 22 ][ 377 ],
   alphaCSR[ 22 ][ 378 ],
   alphaCSR[ 22 ][ 379 ],
   alphaCSR[ 22 ][ 380 ],
   alphaCSR[ 22 ][ 381 ],
   alphaCSR[ 22 ][ 382 ],
   alphaCSR[ 22 ][ 383 ],
   alphaCSR[ 23 ][ 0 ],
   alphaCSR[ 23 ][ 1 ],
   alphaCSR[ 23 ][ 2 ],
   alphaCSR[ 23 ][ 3 ],
   alphaCSR[ 23 ][ 4 ],
   alphaCSR[ 23 ][ 5 ],
   alphaCSR[ 23 ][ 6 ],
   alphaCSR[ 23 ][ 7 ],
   alphaCSR[ 23 ][ 8 ],
   alphaCSR[ 23 ][ 9 ],
   alphaCSR[ 23 ][ 10 ],
   alphaCSR[ 23 ][ 11 ],
   alphaCSR[ 23 ][ 12 ],
   alphaCSR[ 23 ][ 13 ],
   alphaCSR[ 23 ][ 14 ],
   alphaCSR[ 23 ][ 15 ],
   alphaCSR[ 23 ][ 16 ],
   alphaCSR[ 23 ][ 17 ],
   alphaCSR[ 23 ][ 18 ],
   alphaCSR[ 23 ][ 19 ],
   alphaCSR[ 23 ][ 20 ],
   alphaCSR[ 23 ][ 21 ],
   alphaCSR[ 23 ][ 22 ],
   alphaCSR[ 23 ][ 23 ],
   alphaCSR[ 23 ][ 24 ],
   alphaCSR[ 23 ][ 25 ],
   alphaCSR[ 23 ][ 26 ],
   alphaCSR[ 23 ][ 27 ],
   alphaCSR[ 23 ][ 28 ],
   alphaCSR[ 23 ][ 29 ],
   alphaCSR[ 23 ][ 30 ],
   alphaCSR[ 23 ][ 31 ],
   alphaCSR[ 23 ][ 32 ],
   alphaCSR[ 23 ][ 33 ],
   alphaCSR[ 23 ][ 34 ],
   alphaCSR[ 23 ][ 35 ],
   alphaCSR[ 23 ][ 36 ],
   alphaCSR[ 23 ][ 37 ],
   alphaCSR[ 23 ][ 38 ],
   alphaCSR[ 23 ][ 39 ],
   alphaCSR[ 23 ][ 40 ],
   alphaCSR[ 23 ][ 41 ],
   alphaCSR[ 23 ][ 42 ],
   alphaCSR[ 23 ][ 43 ],
   alphaCSR[ 23 ][ 44 ],
   alphaCSR[ 23 ][ 45 ],
   alphaCSR[ 23 ][ 46 ],
   alphaCSR[ 23 ][ 47 ],
   alphaCSR[ 23 ][ 48 ],
   alphaCSR[ 23 ][ 49 ],
   alphaCSR[ 23 ][ 50 ],
   alphaCSR[ 23 ][ 51 ],
   alphaCSR[ 23 ][ 52 ],
   alphaCSR[ 23 ][ 53 ],
   alphaCSR[ 23 ][ 54 ],
   alphaCSR[ 23 ][ 55 ],
   alphaCSR[ 23 ][ 56 ],
   alphaCSR[ 23 ][ 57 ],
   alphaCSR[ 23 ][ 58 ],
   alphaCSR[ 23 ][ 59 ],
   alphaCSR[ 23 ][ 60 ],
   alphaCSR[ 23 ][ 61 ],
   alphaCSR[ 23 ][ 62 ],
   alphaCSR[ 23 ][ 63 ],
   alphaCSR[ 23 ][ 64 ],
   alphaCSR[ 23 ][ 65 ],
   alphaCSR[ 23 ][ 66 ],
   alphaCSR[ 23 ][ 67 ],
   alphaCSR[ 23 ][ 68 ],
   alphaCSR[ 23 ][ 69 ],
   alphaCSR[ 23 ][ 70 ],
   alphaCSR[ 23 ][ 71 ],
   alphaCSR[ 23 ][ 72 ],
   alphaCSR[ 23 ][ 73 ],
   alphaCSR[ 23 ][ 74 ],
   alphaCSR[ 23 ][ 75 ],
   alphaCSR[ 23 ][ 76 ],
   alphaCSR[ 23 ][ 77 ],
   alphaCSR[ 23 ][ 78 ],
   alphaCSR[ 23 ][ 79 ],
   alphaCSR[ 23 ][ 80 ],
   alphaCSR[ 23 ][ 81 ],
   alphaCSR[ 23 ][ 82 ],
   alphaCSR[ 23 ][ 83 ],
   alphaCSR[ 23 ][ 84 ],
   alphaCSR[ 23 ][ 85 ],
   alphaCSR[ 23 ][ 86 ],
   alphaCSR[ 23 ][ 87 ],
   alphaCSR[ 23 ][ 88 ],
   alphaCSR[ 23 ][ 89 ],
   alphaCSR[ 23 ][ 90 ],
   alphaCSR[ 23 ][ 91 ],
   alphaCSR[ 23 ][ 92 ],
   alphaCSR[ 23 ][ 93 ],
   alphaCSR[ 23 ][ 94 ],
   alphaCSR[ 23 ][ 95 ],
   alphaCSR[ 23 ][ 96 ],
   alphaCSR[ 23 ][ 97 ],
   alphaCSR[ 23 ][ 98 ],
   alphaCSR[ 23 ][ 99 ],
   alphaCSR[ 23 ][ 100 ],
   alphaCSR[ 23 ][ 101 ],
   alphaCSR[ 23 ][ 102 ],
   alphaCSR[ 23 ][ 103 ],
   alphaCSR[ 23 ][ 104 ],
   alphaCSR[ 23 ][ 105 ],
   alphaCSR[ 23 ][ 106 ],
   alphaCSR[ 23 ][ 107 ],
   alphaCSR[ 23 ][ 108 ],
   alphaCSR[ 23 ][ 109 ],
   alphaCSR[ 23 ][ 110 ],
   alphaCSR[ 23 ][ 111 ],
   alphaCSR[ 23 ][ 112 ],
   alphaCSR[ 23 ][ 113 ],
   alphaCSR[ 23 ][ 114 ],
   alphaCSR[ 23 ][ 115 ],
   alphaCSR[ 23 ][ 116 ],
   alphaCSR[ 23 ][ 117 ],
   alphaCSR[ 23 ][ 118 ],
   alphaCSR[ 23 ][ 119 ],
   alphaCSR[ 23 ][ 120 ],
   alphaCSR[ 23 ][ 121 ],
   alphaCSR[ 23 ][ 122 ],
   alphaCSR[ 23 ][ 123 ],
   alphaCSR[ 23 ][ 124 ],
   alphaCSR[ 23 ][ 125 ],
   alphaCSR[ 23 ][ 126 ],
   alphaCSR[ 23 ][ 127 ],
   alphaCSR[ 23 ][ 128 ],
   alphaCSR[ 23 ][ 129 ],
   alphaCSR[ 23 ][ 130 ],
   alphaCSR[ 23 ][ 131 ],
   alphaCSR[ 23 ][ 132 ],
   alphaCSR[ 23 ][ 133 ],
   alphaCSR[ 23 ][ 134 ],
   alphaCSR[ 23 ][ 135 ],
   alphaCSR[ 23 ][ 136 ],
   alphaCSR[ 23 ][ 137 ],
   alphaCSR[ 23 ][ 138 ],
   alphaCSR[ 23 ][ 139 ],
   alphaCSR[ 23 ][ 140 ],
   alphaCSR[ 23 ][ 141 ],
   alphaCSR[ 23 ][ 142 ],
   alphaCSR[ 23 ][ 143 ],
   alphaCSR[ 23 ][ 144 ],
   alphaCSR[ 23 ][ 145 ],
   alphaCSR[ 23 ][ 146 ],
   alphaCSR[ 23 ][ 147 ],
   alphaCSR[ 23 ][ 148 ],
   alphaCSR[ 23 ][ 149 ],
   alphaCSR[ 23 ][ 150 ],
   alphaCSR[ 23 ][ 151 ],
   alphaCSR[ 23 ][ 152 ],
   alphaCSR[ 23 ][ 153 ],
   alphaCSR[ 23 ][ 154 ],
   alphaCSR[ 23 ][ 155 ],
   alphaCSR[ 23 ][ 156 ],
   alphaCSR[ 23 ][ 157 ],
   alphaCSR[ 23 ][ 158 ],
   alphaCSR[ 23 ][ 159 ],
   alphaCSR[ 23 ][ 160 ],
   alphaCSR[ 23 ][ 161 ],
   alphaCSR[ 23 ][ 162 ],
   alphaCSR[ 23 ][ 163 ],
   alphaCSR[ 23 ][ 164 ],
   alphaCSR[ 23 ][ 165 ],
   alphaCSR[ 23 ][ 166 ],
   alphaCSR[ 23 ][ 167 ],
   alphaCSR[ 23 ][ 168 ],
   alphaCSR[ 23 ][ 169 ],
   alphaCSR[ 23 ][ 170 ],
   alphaCSR[ 23 ][ 171 ],
   alphaCSR[ 23 ][ 172 ],
   alphaCSR[ 23 ][ 173 ],
   alphaCSR[ 23 ][ 174 ],
   alphaCSR[ 23 ][ 175 ],
   alphaCSR[ 23 ][ 176 ],
   alphaCSR[ 23 ][ 177 ],
   alphaCSR[ 23 ][ 178 ],
   alphaCSR[ 23 ][ 179 ],
   alphaCSR[ 23 ][ 180 ],
   alphaCSR[ 23 ][ 181 ],
   alphaCSR[ 23 ][ 182 ],
   alphaCSR[ 23 ][ 183 ],
   alphaCSR[ 23 ][ 184 ],
   alphaCSR[ 23 ][ 185 ],
   alphaCSR[ 23 ][ 186 ],
   alphaCSR[ 23 ][ 187 ],
   alphaCSR[ 23 ][ 188 ],
   alphaCSR[ 23 ][ 189 ],
   alphaCSR[ 23 ][ 190 ],
   alphaCSR[ 23 ][ 191 ],
   alphaCSR[ 23 ][ 192 ],
   alphaCSR[ 23 ][ 193 ],
   alphaCSR[ 23 ][ 194 ],
   alphaCSR[ 23 ][ 195 ],
   alphaCSR[ 23 ][ 196 ],
   alphaCSR[ 23 ][ 197 ],
   alphaCSR[ 23 ][ 198 ],
   alphaCSR[ 23 ][ 199 ],
   alphaCSR[ 23 ][ 200 ],
   alphaCSR[ 23 ][ 201 ],
   alphaCSR[ 23 ][ 202 ],
   alphaCSR[ 23 ][ 203 ],
   alphaCSR[ 23 ][ 204 ],
   alphaCSR[ 23 ][ 205 ],
   alphaCSR[ 23 ][ 206 ],
   alphaCSR[ 23 ][ 207 ],
   alphaCSR[ 23 ][ 208 ],
   alphaCSR[ 23 ][ 209 ],
   alphaCSR[ 23 ][ 210 ],
   alphaCSR[ 23 ][ 211 ],
   alphaCSR[ 23 ][ 212 ],
   alphaCSR[ 23 ][ 213 ],
   alphaCSR[ 23 ][ 214 ],
   alphaCSR[ 23 ][ 215 ],
   alphaCSR[ 23 ][ 216 ],
   alphaCSR[ 23 ][ 217 ],
   alphaCSR[ 23 ][ 218 ],
   alphaCSR[ 23 ][ 219 ],
   alphaCSR[ 23 ][ 220 ],
   alphaCSR[ 23 ][ 221 ],
   alphaCSR[ 23 ][ 222 ],
   alphaCSR[ 23 ][ 223 ],
   alphaCSR[ 23 ][ 224 ],
   alphaCSR[ 23 ][ 225 ],
   alphaCSR[ 23 ][ 226 ],
   alphaCSR[ 23 ][ 227 ],
   alphaCSR[ 23 ][ 228 ],
   alphaCSR[ 23 ][ 229 ],
   alphaCSR[ 23 ][ 230 ],
   alphaCSR[ 23 ][ 231 ],
   alphaCSR[ 23 ][ 232 ],
   alphaCSR[ 23 ][ 233 ],
   alphaCSR[ 23 ][ 234 ],
   alphaCSR[ 23 ][ 235 ],
   alphaCSR[ 23 ][ 236 ],
   alphaCSR[ 23 ][ 237 ],
   alphaCSR[ 23 ][ 238 ],
   alphaCSR[ 23 ][ 239 ],
   alphaCSR[ 23 ][ 240 ],
   alphaCSR[ 23 ][ 241 ],
   alphaCSR[ 23 ][ 242 ],
   alphaCSR[ 23 ][ 243 ],
   alphaCSR[ 23 ][ 244 ],
   alphaCSR[ 23 ][ 245 ],
   alphaCSR[ 23 ][ 246 ],
   alphaCSR[ 23 ][ 247 ],
   alphaCSR[ 23 ][ 248 ],
   alphaCSR[ 23 ][ 249 ],
   alphaCSR[ 23 ][ 250 ],
   alphaCSR[ 23 ][ 251 ],
   alphaCSR[ 23 ][ 252 ],
   alphaCSR[ 23 ][ 253 ],
   alphaCSR[ 23 ][ 254 ],
   alphaCSR[ 23 ][ 255 ],
   alphaCSR[ 23 ][ 256 ],
   alphaCSR[ 23 ][ 257 ],
   alphaCSR[ 23 ][ 258 ],
   alphaCSR[ 23 ][ 259 ],
   alphaCSR[ 23 ][ 260 ],
   alphaCSR[ 23 ][ 261 ],
   alphaCSR[ 23 ][ 262 ],
   alphaCSR[ 23 ][ 263 ],
   alphaCSR[ 23 ][ 264 ],
   alphaCSR[ 23 ][ 265 ],
   alphaCSR[ 23 ][ 266 ],
   alphaCSR[ 23 ][ 267 ],
   alphaCSR[ 23 ][ 268 ],
   alphaCSR[ 23 ][ 269 ],
   alphaCSR[ 23 ][ 270 ],
   alphaCSR[ 23 ][ 271 ],
   alphaCSR[ 23 ][ 272 ],
   alphaCSR[ 23 ][ 273 ],
   alphaCSR[ 23 ][ 274 ],
   alphaCSR[ 23 ][ 275 ],
   alphaCSR[ 23 ][ 276 ],
   alphaCSR[ 23 ][ 277 ],
   alphaCSR[ 23 ][ 278 ],
   alphaCSR[ 23 ][ 279 ],
   alphaCSR[ 23 ][ 280 ],
   alphaCSR[ 23 ][ 281 ],
   alphaCSR[ 23 ][ 282 ],
   alphaCSR[ 23 ][ 283 ],
   alphaCSR[ 23 ][ 284 ],
   alphaCSR[ 23 ][ 285 ],
   alphaCSR[ 23 ][ 286 ],
   alphaCSR[ 23 ][ 287 ],
   alphaCSR[ 23 ][ 288 ],
   alphaCSR[ 23 ][ 289 ],
   alphaCSR[ 23 ][ 290 ],
   alphaCSR[ 23 ][ 291 ],
   alphaCSR[ 23 ][ 292 ],
   alphaCSR[ 23 ][ 293 ],
   alphaCSR[ 23 ][ 294 ],
   alphaCSR[ 23 ][ 295 ],
   alphaCSR[ 23 ][ 296 ],
   alphaCSR[ 23 ][ 297 ],
   alphaCSR[ 23 ][ 298 ],
   alphaCSR[ 23 ][ 299 ],
   alphaCSR[ 23 ][ 300 ],
   alphaCSR[ 23 ][ 301 ],
   alphaCSR[ 23 ][ 302 ],
   alphaCSR[ 23 ][ 303 ],
   alphaCSR[ 23 ][ 304 ],
   alphaCSR[ 23 ][ 305 ],
   alphaCSR[ 23 ][ 306 ],
   alphaCSR[ 23 ][ 307 ],
   alphaCSR[ 23 ][ 308 ],
   alphaCSR[ 23 ][ 309 ],
   alphaCSR[ 23 ][ 310 ],
   alphaCSR[ 23 ][ 311 ],
   alphaCSR[ 23 ][ 312 ],
   alphaCSR[ 23 ][ 313 ],
   alphaCSR[ 23 ][ 314 ],
   alphaCSR[ 23 ][ 315 ],
   alphaCSR[ 23 ][ 316 ],
   alphaCSR[ 23 ][ 317 ],
   alphaCSR[ 23 ][ 318 ],
   alphaCSR[ 23 ][ 319 ],
   alphaCSR[ 23 ][ 320 ],
   alphaCSR[ 23 ][ 321 ],
   alphaCSR[ 23 ][ 322 ],
   alphaCSR[ 23 ][ 323 ],
   alphaCSR[ 23 ][ 324 ],
   alphaCSR[ 23 ][ 325 ],
   alphaCSR[ 23 ][ 326 ],
   alphaCSR[ 23 ][ 327 ],
   alphaCSR[ 23 ][ 328 ],
   alphaCSR[ 23 ][ 329 ],
   alphaCSR[ 23 ][ 330 ],
   alphaCSR[ 23 ][ 331 ],
   alphaCSR[ 23 ][ 332 ],
   alphaCSR[ 23 ][ 333 ],
   alphaCSR[ 23 ][ 334 ],
   alphaCSR[ 23 ][ 335 ],
   alphaCSR[ 23 ][ 336 ],
   alphaCSR[ 23 ][ 337 ],
   alphaCSR[ 23 ][ 338 ],
   alphaCSR[ 23 ][ 339 ],
   alphaCSR[ 23 ][ 340 ],
   alphaCSR[ 23 ][ 341 ],
   alphaCSR[ 23 ][ 342 ],
   alphaCSR[ 23 ][ 343 ],
   alphaCSR[ 23 ][ 344 ],
   alphaCSR[ 23 ][ 345 ],
   alphaCSR[ 23 ][ 346 ],
   alphaCSR[ 23 ][ 347 ],
   alphaCSR[ 23 ][ 348 ],
   alphaCSR[ 23 ][ 349 ],
   alphaCSR[ 23 ][ 350 ],
   alphaCSR[ 23 ][ 351 ],
   alphaCSR[ 23 ][ 352 ],
   alphaCSR[ 23 ][ 353 ],
   alphaCSR[ 23 ][ 354 ],
   alphaCSR[ 23 ][ 355 ],
   alphaCSR[ 23 ][ 356 ],
   alphaCSR[ 23 ][ 357 ],
   alphaCSR[ 23 ][ 358 ],
   alphaCSR[ 23 ][ 359 ],
   alphaCSR[ 23 ][ 360 ],
   alphaCSR[ 23 ][ 361 ],
   alphaCSR[ 23 ][ 362 ],
   alphaCSR[ 23 ][ 363 ],
   alphaCSR[ 23 ][ 364 ],
   alphaCSR[ 23 ][ 365 ],
   alphaCSR[ 23 ][ 366 ],
   alphaCSR[ 23 ][ 367 ],
   alphaCSR[ 23 ][ 368 ],
   alphaCSR[ 23 ][ 369 ],
   alphaCSR[ 23 ][ 370 ],
   alphaCSR[ 23 ][ 371 ],
   alphaCSR[ 23 ][ 372 ],
   alphaCSR[ 23 ][ 373 ],
   alphaCSR[ 23 ][ 374 ],
   alphaCSR[ 23 ][ 375 ],
   alphaCSR[ 23 ][ 376 ],
   alphaCSR[ 23 ][ 377 ],
   alphaCSR[ 23 ][ 378 ],
   alphaCSR[ 23 ][ 379 ],
   alphaCSR[ 23 ][ 380 ],
   alphaCSR[ 23 ][ 381 ],
   alphaCSR[ 23 ][ 382 ],
   alphaCSR[ 23 ][ 383 ],
   alphaCSR[ 24 ][ 0 ],
   alphaCSR[ 24 ][ 1 ],
   alphaCSR[ 24 ][ 2 ],
   alphaCSR[ 24 ][ 3 ],
   alphaCSR[ 24 ][ 4 ],
   alphaCSR[ 24 ][ 5 ],
   alphaCSR[ 24 ][ 6 ],
   alphaCSR[ 24 ][ 7 ],
   alphaCSR[ 24 ][ 8 ],
   alphaCSR[ 24 ][ 9 ],
   alphaCSR[ 24 ][ 10 ],
   alphaCSR[ 24 ][ 11 ],
   alphaCSR[ 24 ][ 12 ],
   alphaCSR[ 24 ][ 13 ],
   alphaCSR[ 24 ][ 14 ],
   alphaCSR[ 24 ][ 15 ],
   alphaCSR[ 24 ][ 16 ],
   alphaCSR[ 24 ][ 17 ],
   alphaCSR[ 24 ][ 18 ],
   alphaCSR[ 24 ][ 19 ],
   alphaCSR[ 24 ][ 20 ],
   alphaCSR[ 24 ][ 21 ],
   alphaCSR[ 24 ][ 22 ],
   alphaCSR[ 24 ][ 23 ],
   alphaCSR[ 24 ][ 24 ],
   alphaCSR[ 24 ][ 25 ],
   alphaCSR[ 24 ][ 26 ],
   alphaCSR[ 24 ][ 27 ],
   alphaCSR[ 24 ][ 28 ],
   alphaCSR[ 24 ][ 29 ],
   alphaCSR[ 24 ][ 30 ],
   alphaCSR[ 24 ][ 31 ],
   alphaCSR[ 24 ][ 32 ],
   alphaCSR[ 24 ][ 33 ],
   alphaCSR[ 24 ][ 34 ],
   alphaCSR[ 24 ][ 35 ],
   alphaCSR[ 24 ][ 36 ],
   alphaCSR[ 24 ][ 37 ],
   alphaCSR[ 24 ][ 38 ],
   alphaCSR[ 24 ][ 39 ],
   alphaCSR[ 24 ][ 40 ],
   alphaCSR[ 24 ][ 41 ],
   alphaCSR[ 24 ][ 42 ],
   alphaCSR[ 24 ][ 43 ],
   alphaCSR[ 24 ][ 44 ],
   alphaCSR[ 24 ][ 45 ],
   alphaCSR[ 24 ][ 46 ],
   alphaCSR[ 24 ][ 47 ],
   alphaCSR[ 24 ][ 48 ],
   alphaCSR[ 24 ][ 49 ],
   alphaCSR[ 24 ][ 50 ],
   alphaCSR[ 24 ][ 51 ],
   alphaCSR[ 24 ][ 52 ],
   alphaCSR[ 24 ][ 53 ],
   alphaCSR[ 24 ][ 54 ],
   alphaCSR[ 24 ][ 55 ],
   alphaCSR[ 24 ][ 56 ],
   alphaCSR[ 24 ][ 57 ],
   alphaCSR[ 24 ][ 58 ],
   alphaCSR[ 24 ][ 59 ],
   alphaCSR[ 24 ][ 60 ],
   alphaCSR[ 24 ][ 61 ],
   alphaCSR[ 24 ][ 62 ],
   alphaCSR[ 24 ][ 63 ],
   alphaCSR[ 24 ][ 64 ],
   alphaCSR[ 24 ][ 65 ],
   alphaCSR[ 24 ][ 66 ],
   alphaCSR[ 24 ][ 67 ],
   alphaCSR[ 24 ][ 68 ],
   alphaCSR[ 24 ][ 69 ],
   alphaCSR[ 24 ][ 70 ],
   alphaCSR[ 24 ][ 71 ],
   alphaCSR[ 24 ][ 72 ],
   alphaCSR[ 24 ][ 73 ],
   alphaCSR[ 24 ][ 74 ],
   alphaCSR[ 24 ][ 75 ],
   alphaCSR[ 24 ][ 76 ],
   alphaCSR[ 24 ][ 77 ],
   alphaCSR[ 24 ][ 78 ],
   alphaCSR[ 24 ][ 79 ],
   alphaCSR[ 24 ][ 80 ],
   alphaCSR[ 24 ][ 81 ],
   alphaCSR[ 24 ][ 82 ],
   alphaCSR[ 24 ][ 83 ],
   alphaCSR[ 24 ][ 84 ],
   alphaCSR[ 24 ][ 85 ],
   alphaCSR[ 24 ][ 86 ],
   alphaCSR[ 24 ][ 87 ],
   alphaCSR[ 24 ][ 88 ],
   alphaCSR[ 24 ][ 89 ],
   alphaCSR[ 24 ][ 90 ],
   alphaCSR[ 24 ][ 91 ],
   alphaCSR[ 24 ][ 92 ],
   alphaCSR[ 24 ][ 93 ],
   alphaCSR[ 24 ][ 94 ],
   alphaCSR[ 24 ][ 95 ],
   alphaCSR[ 24 ][ 96 ],
   alphaCSR[ 24 ][ 97 ],
   alphaCSR[ 24 ][ 98 ],
   alphaCSR[ 24 ][ 99 ],
   alphaCSR[ 24 ][ 100 ],
   alphaCSR[ 24 ][ 101 ],
   alphaCSR[ 24 ][ 102 ],
   alphaCSR[ 24 ][ 103 ],
   alphaCSR[ 24 ][ 104 ],
   alphaCSR[ 24 ][ 105 ],
   alphaCSR[ 24 ][ 106 ],
   alphaCSR[ 24 ][ 107 ],
   alphaCSR[ 24 ][ 108 ],
   alphaCSR[ 24 ][ 109 ],
   alphaCSR[ 24 ][ 110 ],
   alphaCSR[ 24 ][ 111 ],
   alphaCSR[ 24 ][ 112 ],
   alphaCSR[ 24 ][ 113 ],
   alphaCSR[ 24 ][ 114 ],
   alphaCSR[ 24 ][ 115 ],
   alphaCSR[ 24 ][ 116 ],
   alphaCSR[ 24 ][ 117 ],
   alphaCSR[ 24 ][ 118 ],
   alphaCSR[ 24 ][ 119 ],
   alphaCSR[ 24 ][ 120 ],
   alphaCSR[ 24 ][ 121 ],
   alphaCSR[ 24 ][ 122 ],
   alphaCSR[ 24 ][ 123 ],
   alphaCSR[ 24 ][ 124 ],
   alphaCSR[ 24 ][ 125 ],
   alphaCSR[ 24 ][ 126 ],
   alphaCSR[ 24 ][ 127 ],
   alphaCSR[ 24 ][ 128 ],
   alphaCSR[ 24 ][ 129 ],
   alphaCSR[ 24 ][ 130 ],
   alphaCSR[ 24 ][ 131 ],
   alphaCSR[ 24 ][ 132 ],
   alphaCSR[ 24 ][ 133 ],
   alphaCSR[ 24 ][ 134 ],
   alphaCSR[ 24 ][ 135 ],
   alphaCSR[ 24 ][ 136 ],
   alphaCSR[ 24 ][ 137 ],
   alphaCSR[ 24 ][ 138 ],
   alphaCSR[ 24 ][ 139 ],
   alphaCSR[ 24 ][ 140 ],
   alphaCSR[ 24 ][ 141 ],
   alphaCSR[ 24 ][ 142 ],
   alphaCSR[ 24 ][ 143 ],
   alphaCSR[ 24 ][ 144 ],
   alphaCSR[ 24 ][ 145 ],
   alphaCSR[ 24 ][ 146 ],
   alphaCSR[ 24 ][ 147 ],
   alphaCSR[ 24 ][ 148 ],
   alphaCSR[ 24 ][ 149 ],
   alphaCSR[ 24 ][ 150 ],
   alphaCSR[ 24 ][ 151 ],
   alphaCSR[ 24 ][ 152 ],
   alphaCSR[ 24 ][ 153 ],
   alphaCSR[ 24 ][ 154 ],
   alphaCSR[ 24 ][ 155 ],
   alphaCSR[ 24 ][ 156 ],
   alphaCSR[ 24 ][ 157 ],
   alphaCSR[ 24 ][ 158 ],
   alphaCSR[ 24 ][ 159 ],
   alphaCSR[ 24 ][ 160 ],
   alphaCSR[ 24 ][ 161 ],
   alphaCSR[ 24 ][ 162 ],
   alphaCSR[ 24 ][ 163 ],
   alphaCSR[ 24 ][ 164 ],
   alphaCSR[ 24 ][ 165 ],
   alphaCSR[ 24 ][ 166 ],
   alphaCSR[ 24 ][ 167 ],
   alphaCSR[ 24 ][ 168 ],
   alphaCSR[ 24 ][ 169 ],
   alphaCSR[ 24 ][ 170 ],
   alphaCSR[ 24 ][ 171 ],
   alphaCSR[ 24 ][ 172 ],
   alphaCSR[ 24 ][ 173 ],
   alphaCSR[ 24 ][ 174 ],
   alphaCSR[ 24 ][ 175 ],
   alphaCSR[ 24 ][ 176 ],
   alphaCSR[ 24 ][ 177 ],
   alphaCSR[ 24 ][ 178 ],
   alphaCSR[ 24 ][ 179 ],
   alphaCSR[ 24 ][ 180 ],
   alphaCSR[ 24 ][ 181 ],
   alphaCSR[ 24 ][ 182 ],
   alphaCSR[ 24 ][ 183 ],
   alphaCSR[ 24 ][ 184 ],
   alphaCSR[ 24 ][ 185 ],
   alphaCSR[ 24 ][ 186 ],
   alphaCSR[ 24 ][ 187 ],
   alphaCSR[ 24 ][ 188 ],
   alphaCSR[ 24 ][ 189 ],
   alphaCSR[ 24 ][ 190 ],
   alphaCSR[ 24 ][ 191 ],
   alphaCSR[ 24 ][ 192 ],
   alphaCSR[ 24 ][ 193 ],
   alphaCSR[ 24 ][ 194 ],
   alphaCSR[ 24 ][ 195 ],
   alphaCSR[ 24 ][ 196 ],
   alphaCSR[ 24 ][ 197 ],
   alphaCSR[ 24 ][ 198 ],
   alphaCSR[ 24 ][ 199 ],
   alphaCSR[ 24 ][ 200 ],
   alphaCSR[ 24 ][ 201 ],
   alphaCSR[ 24 ][ 202 ],
   alphaCSR[ 24 ][ 203 ],
   alphaCSR[ 24 ][ 204 ],
   alphaCSR[ 24 ][ 205 ],
   alphaCSR[ 24 ][ 206 ],
   alphaCSR[ 24 ][ 207 ],
   alphaCSR[ 24 ][ 208 ],
   alphaCSR[ 24 ][ 209 ],
   alphaCSR[ 24 ][ 210 ],
   alphaCSR[ 24 ][ 211 ],
   alphaCSR[ 24 ][ 212 ],
   alphaCSR[ 24 ][ 213 ],
   alphaCSR[ 24 ][ 214 ],
   alphaCSR[ 24 ][ 215 ],
   alphaCSR[ 24 ][ 216 ],
   alphaCSR[ 24 ][ 217 ],
   alphaCSR[ 24 ][ 218 ],
   alphaCSR[ 24 ][ 219 ],
   alphaCSR[ 24 ][ 220 ],
   alphaCSR[ 24 ][ 221 ],
   alphaCSR[ 24 ][ 222 ],
   alphaCSR[ 24 ][ 223 ],
   alphaCSR[ 24 ][ 224 ],
   alphaCSR[ 24 ][ 225 ],
   alphaCSR[ 24 ][ 226 ],
   alphaCSR[ 24 ][ 227 ],
   alphaCSR[ 24 ][ 228 ],
   alphaCSR[ 24 ][ 229 ],
   alphaCSR[ 24 ][ 230 ],
   alphaCSR[ 24 ][ 231 ],
   alphaCSR[ 24 ][ 232 ],
   alphaCSR[ 24 ][ 233 ],
   alphaCSR[ 24 ][ 234 ],
   alphaCSR[ 24 ][ 235 ],
   alphaCSR[ 24 ][ 236 ],
   alphaCSR[ 24 ][ 237 ],
   alphaCSR[ 24 ][ 238 ],
   alphaCSR[ 24 ][ 239 ],
   alphaCSR[ 24 ][ 240 ],
   alphaCSR[ 24 ][ 241 ],
   alphaCSR[ 24 ][ 242 ],
   alphaCSR[ 24 ][ 243 ],
   alphaCSR[ 24 ][ 244 ],
   alphaCSR[ 24 ][ 245 ],
   alphaCSR[ 24 ][ 246 ],
   alphaCSR[ 24 ][ 247 ],
   alphaCSR[ 24 ][ 248 ],
   alphaCSR[ 24 ][ 249 ],
   alphaCSR[ 24 ][ 250 ],
   alphaCSR[ 24 ][ 251 ],
   alphaCSR[ 24 ][ 252 ],
   alphaCSR[ 24 ][ 253 ],
   alphaCSR[ 24 ][ 254 ],
   alphaCSR[ 24 ][ 255 ],
   alphaCSR[ 24 ][ 256 ],
   alphaCSR[ 24 ][ 257 ],
   alphaCSR[ 24 ][ 258 ],
   alphaCSR[ 24 ][ 259 ],
   alphaCSR[ 24 ][ 260 ],
   alphaCSR[ 24 ][ 261 ],
   alphaCSR[ 24 ][ 262 ],
   alphaCSR[ 24 ][ 263 ],
   alphaCSR[ 24 ][ 264 ],
   alphaCSR[ 24 ][ 265 ],
   alphaCSR[ 24 ][ 266 ],
   alphaCSR[ 24 ][ 267 ],
   alphaCSR[ 24 ][ 268 ],
   alphaCSR[ 24 ][ 269 ],
   alphaCSR[ 24 ][ 270 ],
   alphaCSR[ 24 ][ 271 ],
   alphaCSR[ 24 ][ 272 ],
   alphaCSR[ 24 ][ 273 ],
   alphaCSR[ 24 ][ 274 ],
   alphaCSR[ 24 ][ 275 ],
   alphaCSR[ 24 ][ 276 ],
   alphaCSR[ 24 ][ 277 ],
   alphaCSR[ 24 ][ 278 ],
   alphaCSR[ 24 ][ 279 ],
   alphaCSR[ 24 ][ 280 ],
   alphaCSR[ 24 ][ 281 ],
   alphaCSR[ 24 ][ 282 ],
   alphaCSR[ 24 ][ 283 ],
   alphaCSR[ 24 ][ 284 ],
   alphaCSR[ 24 ][ 285 ],
   alphaCSR[ 24 ][ 286 ],
   alphaCSR[ 24 ][ 287 ],
   alphaCSR[ 24 ][ 288 ],
   alphaCSR[ 24 ][ 289 ],
   alphaCSR[ 24 ][ 290 ],
   alphaCSR[ 24 ][ 291 ],
   alphaCSR[ 24 ][ 292 ],
   alphaCSR[ 24 ][ 293 ],
   alphaCSR[ 24 ][ 294 ],
   alphaCSR[ 24 ][ 295 ],
   alphaCSR[ 24 ][ 296 ],
   alphaCSR[ 24 ][ 297 ],
   alphaCSR[ 24 ][ 298 ],
   alphaCSR[ 24 ][ 299 ],
   alphaCSR[ 24 ][ 300 ],
   alphaCSR[ 24 ][ 301 ],
   alphaCSR[ 24 ][ 302 ],
   alphaCSR[ 24 ][ 303 ],
   alphaCSR[ 24 ][ 304 ],
   alphaCSR[ 24 ][ 305 ],
   alphaCSR[ 24 ][ 306 ],
   alphaCSR[ 24 ][ 307 ],
   alphaCSR[ 24 ][ 308 ],
   alphaCSR[ 24 ][ 309 ],
   alphaCSR[ 24 ][ 310 ],
   alphaCSR[ 24 ][ 311 ],
   alphaCSR[ 24 ][ 312 ],
   alphaCSR[ 24 ][ 313 ],
   alphaCSR[ 24 ][ 314 ],
   alphaCSR[ 24 ][ 315 ],
   alphaCSR[ 24 ][ 316 ],
   alphaCSR[ 24 ][ 317 ],
   alphaCSR[ 24 ][ 318 ],
   alphaCSR[ 24 ][ 319 ],
   alphaCSR[ 24 ][ 320 ],
   alphaCSR[ 24 ][ 321 ],
   alphaCSR[ 24 ][ 322 ],
   alphaCSR[ 24 ][ 323 ],
   alphaCSR[ 24 ][ 324 ],
   alphaCSR[ 24 ][ 325 ],
   alphaCSR[ 24 ][ 326 ],
   alphaCSR[ 24 ][ 327 ],
   alphaCSR[ 24 ][ 328 ],
   alphaCSR[ 24 ][ 329 ],
   alphaCSR[ 24 ][ 330 ],
   alphaCSR[ 24 ][ 331 ],
   alphaCSR[ 24 ][ 332 ],
   alphaCSR[ 24 ][ 333 ],
   alphaCSR[ 24 ][ 334 ],
   alphaCSR[ 24 ][ 335 ],
   alphaCSR[ 24 ][ 336 ],
   alphaCSR[ 24 ][ 337 ],
   alphaCSR[ 24 ][ 338 ],
   alphaCSR[ 24 ][ 339 ],
   alphaCSR[ 24 ][ 340 ],
   alphaCSR[ 24 ][ 341 ],
   alphaCSR[ 24 ][ 342 ],
   alphaCSR[ 24 ][ 343 ],
   alphaCSR[ 24 ][ 344 ],
   alphaCSR[ 24 ][ 345 ],
   alphaCSR[ 24 ][ 346 ],
   alphaCSR[ 24 ][ 347 ],
   alphaCSR[ 24 ][ 348 ],
   alphaCSR[ 24 ][ 349 ],
   alphaCSR[ 24 ][ 350 ],
   alphaCSR[ 24 ][ 351 ],
   alphaCSR[ 24 ][ 352 ],
   alphaCSR[ 24 ][ 353 ],
   alphaCSR[ 24 ][ 354 ],
   alphaCSR[ 24 ][ 355 ],
   alphaCSR[ 24 ][ 356 ],
   alphaCSR[ 24 ][ 357 ],
   alphaCSR[ 24 ][ 358 ],
   alphaCSR[ 24 ][ 359 ],
   alphaCSR[ 24 ][ 360 ],
   alphaCSR[ 24 ][ 361 ],
   alphaCSR[ 24 ][ 362 ],
   alphaCSR[ 24 ][ 363 ],
   alphaCSR[ 24 ][ 364 ],
   alphaCSR[ 24 ][ 365 ],
   alphaCSR[ 24 ][ 366 ],
   alphaCSR[ 24 ][ 367 ],
   alphaCSR[ 24 ][ 368 ],
   alphaCSR[ 24 ][ 369 ],
   alphaCSR[ 24 ][ 370 ],
   alphaCSR[ 24 ][ 371 ],
   alphaCSR[ 24 ][ 372 ],
   alphaCSR[ 24 ][ 373 ],
   alphaCSR[ 24 ][ 374 ],
   alphaCSR[ 24 ][ 375 ],
   alphaCSR[ 24 ][ 376 ],
   alphaCSR[ 24 ][ 377 ],
   alphaCSR[ 24 ][ 378 ],
   alphaCSR[ 24 ][ 379 ],
   alphaCSR[ 24 ][ 380 ],
   alphaCSR[ 24 ][ 381 ],
   alphaCSR[ 24 ][ 382 ],
   alphaCSR[ 24 ][ 383 ],
   alphaCSR[ 25 ][ 0 ],
   alphaCSR[ 25 ][ 1 ],
   alphaCSR[ 25 ][ 2 ],
   alphaCSR[ 25 ][ 3 ],
   alphaCSR[ 25 ][ 4 ],
   alphaCSR[ 25 ][ 5 ],
   alphaCSR[ 25 ][ 6 ],
   alphaCSR[ 25 ][ 7 ],
   alphaCSR[ 25 ][ 8 ],
   alphaCSR[ 25 ][ 9 ],
   alphaCSR[ 25 ][ 10 ],
   alphaCSR[ 25 ][ 11 ],
   alphaCSR[ 25 ][ 12 ],
   alphaCSR[ 25 ][ 13 ],
   alphaCSR[ 25 ][ 14 ],
   alphaCSR[ 25 ][ 15 ],
   alphaCSR[ 25 ][ 16 ],
   alphaCSR[ 25 ][ 17 ],
   alphaCSR[ 25 ][ 18 ],
   alphaCSR[ 25 ][ 19 ],
   alphaCSR[ 25 ][ 20 ],
   alphaCSR[ 25 ][ 21 ],
   alphaCSR[ 25 ][ 22 ],
   alphaCSR[ 25 ][ 23 ],
   alphaCSR[ 25 ][ 24 ],
   alphaCSR[ 25 ][ 25 ],
   alphaCSR[ 25 ][ 26 ],
   alphaCSR[ 25 ][ 27 ],
   alphaCSR[ 25 ][ 28 ],
   alphaCSR[ 25 ][ 29 ],
   alphaCSR[ 25 ][ 30 ],
   alphaCSR[ 25 ][ 31 ],
   alphaCSR[ 25 ][ 32 ],
   alphaCSR[ 25 ][ 33 ],
   alphaCSR[ 25 ][ 34 ],
   alphaCSR[ 25 ][ 35 ],
   alphaCSR[ 25 ][ 36 ],
   alphaCSR[ 25 ][ 37 ],
   alphaCSR[ 25 ][ 38 ],
   alphaCSR[ 25 ][ 39 ],
   alphaCSR[ 25 ][ 40 ],
   alphaCSR[ 25 ][ 41 ],
   alphaCSR[ 25 ][ 42 ],
   alphaCSR[ 25 ][ 43 ],
   alphaCSR[ 25 ][ 44 ],
   alphaCSR[ 25 ][ 45 ],
   alphaCSR[ 25 ][ 46 ],
   alphaCSR[ 25 ][ 47 ],
   alphaCSR[ 25 ][ 48 ],
   alphaCSR[ 25 ][ 49 ],
   alphaCSR[ 25 ][ 50 ],
   alphaCSR[ 25 ][ 51 ],
   alphaCSR[ 25 ][ 52 ],
   alphaCSR[ 25 ][ 53 ],
   alphaCSR[ 25 ][ 54 ],
   alphaCSR[ 25 ][ 55 ],
   alphaCSR[ 25 ][ 56 ],
   alphaCSR[ 25 ][ 57 ],
   alphaCSR[ 25 ][ 58 ],
   alphaCSR[ 25 ][ 59 ],
   alphaCSR[ 25 ][ 60 ],
   alphaCSR[ 25 ][ 61 ],
   alphaCSR[ 25 ][ 62 ],
   alphaCSR[ 25 ][ 63 ],
   alphaCSR[ 25 ][ 64 ],
   alphaCSR[ 25 ][ 65 ],
   alphaCSR[ 25 ][ 66 ],
   alphaCSR[ 25 ][ 67 ],
   alphaCSR[ 25 ][ 68 ],
   alphaCSR[ 25 ][ 69 ],
   alphaCSR[ 25 ][ 70 ],
   alphaCSR[ 25 ][ 71 ],
   alphaCSR[ 25 ][ 72 ],
   alphaCSR[ 25 ][ 73 ],
   alphaCSR[ 25 ][ 74 ],
   alphaCSR[ 25 ][ 75 ],
   alphaCSR[ 25 ][ 76 ],
   alphaCSR[ 25 ][ 77 ],
   alphaCSR[ 25 ][ 78 ],
   alphaCSR[ 25 ][ 79 ],
   alphaCSR[ 25 ][ 80 ],
   alphaCSR[ 25 ][ 81 ],
   alphaCSR[ 25 ][ 82 ],
   alphaCSR[ 25 ][ 83 ],
   alphaCSR[ 25 ][ 84 ],
   alphaCSR[ 25 ][ 85 ],
   alphaCSR[ 25 ][ 86 ],
   alphaCSR[ 25 ][ 87 ],
   alphaCSR[ 25 ][ 88 ],
   alphaCSR[ 25 ][ 89 ],
   alphaCSR[ 25 ][ 90 ],
   alphaCSR[ 25 ][ 91 ],
   alphaCSR[ 25 ][ 92 ],
   alphaCSR[ 25 ][ 93 ],
   alphaCSR[ 25 ][ 94 ],
   alphaCSR[ 25 ][ 95 ],
   alphaCSR[ 25 ][ 96 ],
   alphaCSR[ 25 ][ 97 ],
   alphaCSR[ 25 ][ 98 ],
   alphaCSR[ 25 ][ 99 ],
   alphaCSR[ 25 ][ 100 ],
   alphaCSR[ 25 ][ 101 ],
   alphaCSR[ 25 ][ 102 ],
   alphaCSR[ 25 ][ 103 ],
   alphaCSR[ 25 ][ 104 ],
   alphaCSR[ 25 ][ 105 ],
   alphaCSR[ 25 ][ 106 ],
   alphaCSR[ 25 ][ 107 ],
   alphaCSR[ 25 ][ 108 ],
   alphaCSR[ 25 ][ 109 ],
   alphaCSR[ 25 ][ 110 ],
   alphaCSR[ 25 ][ 111 ],
   alphaCSR[ 25 ][ 112 ],
   alphaCSR[ 25 ][ 113 ],
   alphaCSR[ 25 ][ 114 ],
   alphaCSR[ 25 ][ 115 ],
   alphaCSR[ 25 ][ 116 ],
   alphaCSR[ 25 ][ 117 ],
   alphaCSR[ 25 ][ 118 ],
   alphaCSR[ 25 ][ 119 ],
   alphaCSR[ 25 ][ 120 ],
   alphaCSR[ 25 ][ 121 ],
   alphaCSR[ 25 ][ 122 ],
   alphaCSR[ 25 ][ 123 ],
   alphaCSR[ 25 ][ 124 ],
   alphaCSR[ 25 ][ 125 ],
   alphaCSR[ 25 ][ 126 ],
   alphaCSR[ 25 ][ 127 ],
   alphaCSR[ 25 ][ 128 ],
   alphaCSR[ 25 ][ 129 ],
   alphaCSR[ 25 ][ 130 ],
   alphaCSR[ 25 ][ 131 ],
   alphaCSR[ 25 ][ 132 ],
   alphaCSR[ 25 ][ 133 ],
   alphaCSR[ 25 ][ 134 ],
   alphaCSR[ 25 ][ 135 ],
   alphaCSR[ 25 ][ 136 ],
   alphaCSR[ 25 ][ 137 ],
   alphaCSR[ 25 ][ 138 ],
   alphaCSR[ 25 ][ 139 ],
   alphaCSR[ 25 ][ 140 ],
   alphaCSR[ 25 ][ 141 ],
   alphaCSR[ 25 ][ 142 ],
   alphaCSR[ 25 ][ 143 ],
   alphaCSR[ 25 ][ 144 ],
   alphaCSR[ 25 ][ 145 ],
   alphaCSR[ 25 ][ 146 ],
   alphaCSR[ 25 ][ 147 ],
   alphaCSR[ 25 ][ 148 ],
   alphaCSR[ 25 ][ 149 ],
   alphaCSR[ 25 ][ 150 ],
   alphaCSR[ 25 ][ 151 ],
   alphaCSR[ 25 ][ 152 ],
   alphaCSR[ 25 ][ 153 ],
   alphaCSR[ 25 ][ 154 ],
   alphaCSR[ 25 ][ 155 ],
   alphaCSR[ 25 ][ 156 ],
   alphaCSR[ 25 ][ 157 ],
   alphaCSR[ 25 ][ 158 ],
   alphaCSR[ 25 ][ 159 ],
   alphaCSR[ 25 ][ 160 ],
   alphaCSR[ 25 ][ 161 ],
   alphaCSR[ 25 ][ 162 ],
   alphaCSR[ 25 ][ 163 ],
   alphaCSR[ 25 ][ 164 ],
   alphaCSR[ 25 ][ 165 ],
   alphaCSR[ 25 ][ 166 ],
   alphaCSR[ 25 ][ 167 ],
   alphaCSR[ 25 ][ 168 ],
   alphaCSR[ 25 ][ 169 ],
   alphaCSR[ 25 ][ 170 ],
   alphaCSR[ 25 ][ 171 ],
   alphaCSR[ 25 ][ 172 ],
   alphaCSR[ 25 ][ 173 ],
   alphaCSR[ 25 ][ 174 ],
   alphaCSR[ 25 ][ 175 ],
   alphaCSR[ 25 ][ 176 ],
   alphaCSR[ 25 ][ 177 ],
   alphaCSR[ 25 ][ 178 ],
   alphaCSR[ 25 ][ 179 ],
   alphaCSR[ 25 ][ 180 ],
   alphaCSR[ 25 ][ 181 ],
   alphaCSR[ 25 ][ 182 ],
   alphaCSR[ 25 ][ 183 ],
   alphaCSR[ 25 ][ 184 ],
   alphaCSR[ 25 ][ 185 ],
   alphaCSR[ 25 ][ 186 ],
   alphaCSR[ 25 ][ 187 ],
   alphaCSR[ 25 ][ 188 ],
   alphaCSR[ 25 ][ 189 ],
   alphaCSR[ 25 ][ 190 ],
   alphaCSR[ 25 ][ 191 ],
   alphaCSR[ 25 ][ 192 ],
   alphaCSR[ 25 ][ 193 ],
   alphaCSR[ 25 ][ 194 ],
   alphaCSR[ 25 ][ 195 ],
   alphaCSR[ 25 ][ 196 ],
   alphaCSR[ 25 ][ 197 ],
   alphaCSR[ 25 ][ 198 ],
   alphaCSR[ 25 ][ 199 ],
   alphaCSR[ 25 ][ 200 ],
   alphaCSR[ 25 ][ 201 ],
   alphaCSR[ 25 ][ 202 ],
   alphaCSR[ 25 ][ 203 ],
   alphaCSR[ 25 ][ 204 ],
   alphaCSR[ 25 ][ 205 ],
   alphaCSR[ 25 ][ 206 ],
   alphaCSR[ 25 ][ 207 ],
   alphaCSR[ 25 ][ 208 ],
   alphaCSR[ 25 ][ 209 ],
   alphaCSR[ 25 ][ 210 ],
   alphaCSR[ 25 ][ 211 ],
   alphaCSR[ 25 ][ 212 ],
   alphaCSR[ 25 ][ 213 ],
   alphaCSR[ 25 ][ 214 ],
   alphaCSR[ 25 ][ 215 ],
   alphaCSR[ 25 ][ 216 ],
   alphaCSR[ 25 ][ 217 ],
   alphaCSR[ 25 ][ 218 ],
   alphaCSR[ 25 ][ 219 ],
   alphaCSR[ 25 ][ 220 ],
   alphaCSR[ 25 ][ 221 ],
   alphaCSR[ 25 ][ 222 ],
   alphaCSR[ 25 ][ 223 ],
   alphaCSR[ 25 ][ 224 ],
   alphaCSR[ 25 ][ 225 ],
   alphaCSR[ 25 ][ 226 ],
   alphaCSR[ 25 ][ 227 ],
   alphaCSR[ 25 ][ 228 ],
   alphaCSR[ 25 ][ 229 ],
   alphaCSR[ 25 ][ 230 ],
   alphaCSR[ 25 ][ 231 ],
   alphaCSR[ 25 ][ 232 ],
   alphaCSR[ 25 ][ 233 ],
   alphaCSR[ 25 ][ 234 ],
   alphaCSR[ 25 ][ 235 ],
   alphaCSR[ 25 ][ 236 ],
   alphaCSR[ 25 ][ 237 ],
   alphaCSR[ 25 ][ 238 ],
   alphaCSR[ 25 ][ 239 ],
   alphaCSR[ 25 ][ 240 ],
   alphaCSR[ 25 ][ 241 ],
   alphaCSR[ 25 ][ 242 ],
   alphaCSR[ 25 ][ 243 ],
   alphaCSR[ 25 ][ 244 ],
   alphaCSR[ 25 ][ 245 ],
   alphaCSR[ 25 ][ 246 ],
   alphaCSR[ 25 ][ 247 ],
   alphaCSR[ 25 ][ 248 ],
   alphaCSR[ 25 ][ 249 ],
   alphaCSR[ 25 ][ 250 ],
   alphaCSR[ 25 ][ 251 ],
   alphaCSR[ 25 ][ 252 ],
   alphaCSR[ 25 ][ 253 ],
   alphaCSR[ 25 ][ 254 ],
   alphaCSR[ 25 ][ 255 ],
   alphaCSR[ 25 ][ 256 ],
   alphaCSR[ 25 ][ 257 ],
   alphaCSR[ 25 ][ 258 ],
   alphaCSR[ 25 ][ 259 ],
   alphaCSR[ 25 ][ 260 ],
   alphaCSR[ 25 ][ 261 ],
   alphaCSR[ 25 ][ 262 ],
   alphaCSR[ 25 ][ 263 ],
   alphaCSR[ 25 ][ 264 ],
   alphaCSR[ 25 ][ 265 ],
   alphaCSR[ 25 ][ 266 ],
   alphaCSR[ 25 ][ 267 ],
   alphaCSR[ 25 ][ 268 ],
   alphaCSR[ 25 ][ 269 ],
   alphaCSR[ 25 ][ 270 ],
   alphaCSR[ 25 ][ 271 ],
   alphaCSR[ 25 ][ 272 ],
   alphaCSR[ 25 ][ 273 ],
   alphaCSR[ 25 ][ 274 ],
   alphaCSR[ 25 ][ 275 ],
   alphaCSR[ 25 ][ 276 ],
   alphaCSR[ 25 ][ 277 ],
   alphaCSR[ 25 ][ 278 ],
   alphaCSR[ 25 ][ 279 ],
   alphaCSR[ 25 ][ 280 ],
   alphaCSR[ 25 ][ 281 ],
   alphaCSR[ 25 ][ 282 ],
   alphaCSR[ 25 ][ 283 ],
   alphaCSR[ 25 ][ 284 ],
   alphaCSR[ 25 ][ 285 ],
   alphaCSR[ 25 ][ 286 ],
   alphaCSR[ 25 ][ 287 ],
   alphaCSR[ 25 ][ 288 ],
   alphaCSR[ 25 ][ 289 ],
   alphaCSR[ 25 ][ 290 ],
   alphaCSR[ 25 ][ 291 ],
   alphaCSR[ 25 ][ 292 ],
   alphaCSR[ 25 ][ 293 ],
   alphaCSR[ 25 ][ 294 ],
   alphaCSR[ 25 ][ 295 ],
   alphaCSR[ 25 ][ 296 ],
   alphaCSR[ 25 ][ 297 ],
   alphaCSR[ 25 ][ 298 ],
   alphaCSR[ 25 ][ 299 ],
   alphaCSR[ 25 ][ 300 ],
   alphaCSR[ 25 ][ 301 ],
   alphaCSR[ 25 ][ 302 ],
   alphaCSR[ 25 ][ 303 ],
   alphaCSR[ 25 ][ 304 ],
   alphaCSR[ 25 ][ 305 ],
   alphaCSR[ 25 ][ 306 ],
   alphaCSR[ 25 ][ 307 ],
   alphaCSR[ 25 ][ 308 ],
   alphaCSR[ 25 ][ 309 ],
   alphaCSR[ 25 ][ 310 ],
   alphaCSR[ 25 ][ 311 ],
   alphaCSR[ 25 ][ 312 ],
   alphaCSR[ 25 ][ 313 ],
   alphaCSR[ 25 ][ 314 ],
   alphaCSR[ 25 ][ 315 ],
   alphaCSR[ 25 ][ 316 ],
   alphaCSR[ 25 ][ 317 ],
   alphaCSR[ 25 ][ 318 ],
   alphaCSR[ 25 ][ 319 ],
   alphaCSR[ 25 ][ 320 ],
   alphaCSR[ 25 ][ 321 ],
   alphaCSR[ 25 ][ 322 ],
   alphaCSR[ 25 ][ 323 ],
   alphaCSR[ 25 ][ 324 ],
   alphaCSR[ 25 ][ 325 ],
   alphaCSR[ 25 ][ 326 ],
   alphaCSR[ 25 ][ 327 ],
   alphaCSR[ 25 ][ 328 ],
   alphaCSR[ 25 ][ 329 ],
   alphaCSR[ 25 ][ 330 ],
   alphaCSR[ 25 ][ 331 ],
   alphaCSR[ 25 ][ 332 ],
   alphaCSR[ 25 ][ 333 ],
   alphaCSR[ 25 ][ 334 ],
   alphaCSR[ 25 ][ 335 ],
   alphaCSR[ 25 ][ 336 ],
   alphaCSR[ 25 ][ 337 ],
   alphaCSR[ 25 ][ 338 ],
   alphaCSR[ 25 ][ 339 ],
   alphaCSR[ 25 ][ 340 ],
   alphaCSR[ 25 ][ 341 ],
   alphaCSR[ 25 ][ 342 ],
   alphaCSR[ 25 ][ 343 ],
   alphaCSR[ 25 ][ 344 ],
   alphaCSR[ 25 ][ 345 ],
   alphaCSR[ 25 ][ 346 ],
   alphaCSR[ 25 ][ 347 ],
   alphaCSR[ 25 ][ 348 ],
   alphaCSR[ 25 ][ 349 ],
   alphaCSR[ 25 ][ 350 ],
   alphaCSR[ 25 ][ 351 ],
   alphaCSR[ 25 ][ 352 ],
   alphaCSR[ 25 ][ 353 ],
   alphaCSR[ 25 ][ 354 ],
   alphaCSR[ 25 ][ 355 ],
   alphaCSR[ 25 ][ 356 ],
   alphaCSR[ 25 ][ 357 ],
   alphaCSR[ 25 ][ 358 ],
   alphaCSR[ 25 ][ 359 ],
   alphaCSR[ 25 ][ 360 ],
   alphaCSR[ 25 ][ 361 ],
   alphaCSR[ 25 ][ 362 ],
   alphaCSR[ 25 ][ 363 ],
   alphaCSR[ 25 ][ 364 ],
   alphaCSR[ 25 ][ 365 ],
   alphaCSR[ 25 ][ 366 ],
   alphaCSR[ 25 ][ 367 ],
   alphaCSR[ 25 ][ 368 ],
   alphaCSR[ 25 ][ 369 ],
   alphaCSR[ 25 ][ 370 ],
   alphaCSR[ 25 ][ 371 ],
   alphaCSR[ 25 ][ 372 ],
   alphaCSR[ 25 ][ 373 ],
   alphaCSR[ 25 ][ 374 ],
   alphaCSR[ 25 ][ 375 ],
   alphaCSR[ 25 ][ 376 ],
   alphaCSR[ 25 ][ 377 ],
   alphaCSR[ 25 ][ 378 ],
   alphaCSR[ 25 ][ 379 ],
   alphaCSR[ 25 ][ 380 ],
   alphaCSR[ 25 ][ 381 ],
   alphaCSR[ 25 ][ 382 ],
   alphaCSR[ 25 ][ 383 ],
   alphaCSR[ 26 ][ 0 ],
   alphaCSR[ 26 ][ 1 ],
   alphaCSR[ 26 ][ 2 ],
   alphaCSR[ 26 ][ 3 ],
   alphaCSR[ 26 ][ 4 ],
   alphaCSR[ 26 ][ 5 ],
   alphaCSR[ 26 ][ 6 ],
   alphaCSR[ 26 ][ 7 ],
   alphaCSR[ 26 ][ 8 ],
   alphaCSR[ 26 ][ 9 ],
   alphaCSR[ 26 ][ 10 ],
   alphaCSR[ 26 ][ 11 ],
   alphaCSR[ 26 ][ 12 ],
   alphaCSR[ 26 ][ 13 ],
   alphaCSR[ 26 ][ 14 ],
   alphaCSR[ 26 ][ 15 ],
   alphaCSR[ 26 ][ 16 ],
   alphaCSR[ 26 ][ 17 ],
   alphaCSR[ 26 ][ 18 ],
   alphaCSR[ 26 ][ 19 ],
   alphaCSR[ 26 ][ 20 ],
   alphaCSR[ 26 ][ 21 ],
   alphaCSR[ 26 ][ 22 ],
   alphaCSR[ 26 ][ 23 ],
   alphaCSR[ 26 ][ 24 ],
   alphaCSR[ 26 ][ 25 ],
   alphaCSR[ 26 ][ 26 ],
   alphaCSR[ 26 ][ 27 ],
   alphaCSR[ 26 ][ 28 ],
   alphaCSR[ 26 ][ 29 ],
   alphaCSR[ 26 ][ 30 ],
   alphaCSR[ 26 ][ 31 ],
   alphaCSR[ 26 ][ 32 ],
   alphaCSR[ 26 ][ 33 ],
   alphaCSR[ 26 ][ 34 ],
   alphaCSR[ 26 ][ 35 ],
   alphaCSR[ 26 ][ 36 ],
   alphaCSR[ 26 ][ 37 ],
   alphaCSR[ 26 ][ 38 ],
   alphaCSR[ 26 ][ 39 ],
   alphaCSR[ 26 ][ 40 ],
   alphaCSR[ 26 ][ 41 ],
   alphaCSR[ 26 ][ 42 ],
   alphaCSR[ 26 ][ 43 ],
   alphaCSR[ 26 ][ 44 ],
   alphaCSR[ 26 ][ 45 ],
   alphaCSR[ 26 ][ 46 ],
   alphaCSR[ 26 ][ 47 ],
   alphaCSR[ 26 ][ 48 ],
   alphaCSR[ 26 ][ 49 ],
   alphaCSR[ 26 ][ 50 ],
   alphaCSR[ 26 ][ 51 ],
   alphaCSR[ 26 ][ 52 ],
   alphaCSR[ 26 ][ 53 ],
   alphaCSR[ 26 ][ 54 ],
   alphaCSR[ 26 ][ 55 ],
   alphaCSR[ 26 ][ 56 ],
   alphaCSR[ 26 ][ 57 ],
   alphaCSR[ 26 ][ 58 ],
   alphaCSR[ 26 ][ 59 ],
   alphaCSR[ 26 ][ 60 ],
   alphaCSR[ 26 ][ 61 ],
   alphaCSR[ 26 ][ 62 ],
   alphaCSR[ 26 ][ 63 ],
   alphaCSR[ 26 ][ 64 ],
   alphaCSR[ 26 ][ 65 ],
   alphaCSR[ 26 ][ 66 ],
   alphaCSR[ 26 ][ 67 ],
   alphaCSR[ 26 ][ 68 ],
   alphaCSR[ 26 ][ 69 ],
   alphaCSR[ 26 ][ 70 ],
   alphaCSR[ 26 ][ 71 ],
   alphaCSR[ 26 ][ 72 ],
   alphaCSR[ 26 ][ 73 ],
   alphaCSR[ 26 ][ 74 ],
   alphaCSR[ 26 ][ 75 ],
   alphaCSR[ 26 ][ 76 ],
   alphaCSR[ 26 ][ 77 ],
   alphaCSR[ 26 ][ 78 ],
   alphaCSR[ 26 ][ 79 ],
   alphaCSR[ 26 ][ 80 ],
   alphaCSR[ 26 ][ 81 ],
   alphaCSR[ 26 ][ 82 ],
   alphaCSR[ 26 ][ 83 ],
   alphaCSR[ 26 ][ 84 ],
   alphaCSR[ 26 ][ 85 ],
   alphaCSR[ 26 ][ 86 ],
   alphaCSR[ 26 ][ 87 ],
   alphaCSR[ 26 ][ 88 ],
   alphaCSR[ 26 ][ 89 ],
   alphaCSR[ 26 ][ 90 ],
   alphaCSR[ 26 ][ 91 ],
   alphaCSR[ 26 ][ 92 ],
   alphaCSR[ 26 ][ 93 ],
   alphaCSR[ 26 ][ 94 ],
   alphaCSR[ 26 ][ 95 ],
   alphaCSR[ 26 ][ 96 ],
   alphaCSR[ 26 ][ 97 ],
   alphaCSR[ 26 ][ 98 ],
   alphaCSR[ 26 ][ 99 ],
   alphaCSR[ 26 ][ 100 ],
   alphaCSR[ 26 ][ 101 ],
   alphaCSR[ 26 ][ 102 ],
   alphaCSR[ 26 ][ 103 ],
   alphaCSR[ 26 ][ 104 ],
   alphaCSR[ 26 ][ 105 ],
   alphaCSR[ 26 ][ 106 ],
   alphaCSR[ 26 ][ 107 ],
   alphaCSR[ 26 ][ 108 ],
   alphaCSR[ 26 ][ 109 ],
   alphaCSR[ 26 ][ 110 ],
   alphaCSR[ 26 ][ 111 ],
   alphaCSR[ 26 ][ 112 ],
   alphaCSR[ 26 ][ 113 ],
   alphaCSR[ 26 ][ 114 ],
   alphaCSR[ 26 ][ 115 ],
   alphaCSR[ 26 ][ 116 ],
   alphaCSR[ 26 ][ 117 ],
   alphaCSR[ 26 ][ 118 ],
   alphaCSR[ 26 ][ 119 ],
   alphaCSR[ 26 ][ 120 ],
   alphaCSR[ 26 ][ 121 ],
   alphaCSR[ 26 ][ 122 ],
   alphaCSR[ 26 ][ 123 ],
   alphaCSR[ 26 ][ 124 ],
   alphaCSR[ 26 ][ 125 ],
   alphaCSR[ 26 ][ 126 ],
   alphaCSR[ 26 ][ 127 ],
   alphaCSR[ 26 ][ 128 ],
   alphaCSR[ 26 ][ 129 ],
   alphaCSR[ 26 ][ 130 ],
   alphaCSR[ 26 ][ 131 ],
   alphaCSR[ 26 ][ 132 ],
   alphaCSR[ 26 ][ 133 ],
   alphaCSR[ 26 ][ 134 ],
   alphaCSR[ 26 ][ 135 ],
   alphaCSR[ 26 ][ 136 ],
   alphaCSR[ 26 ][ 137 ],
   alphaCSR[ 26 ][ 138 ],
   alphaCSR[ 26 ][ 139 ],
   alphaCSR[ 26 ][ 140 ],
   alphaCSR[ 26 ][ 141 ],
   alphaCSR[ 26 ][ 142 ],
   alphaCSR[ 26 ][ 143 ],
   alphaCSR[ 26 ][ 144 ],
   alphaCSR[ 26 ][ 145 ],
   alphaCSR[ 26 ][ 146 ],
   alphaCSR[ 26 ][ 147 ],
   alphaCSR[ 26 ][ 148 ],
   alphaCSR[ 26 ][ 149 ],
   alphaCSR[ 26 ][ 150 ],
   alphaCSR[ 26 ][ 151 ],
   alphaCSR[ 26 ][ 152 ],
   alphaCSR[ 26 ][ 153 ],
   alphaCSR[ 26 ][ 154 ],
   alphaCSR[ 26 ][ 155 ],
   alphaCSR[ 26 ][ 156 ],
   alphaCSR[ 26 ][ 157 ],
   alphaCSR[ 26 ][ 158 ],
   alphaCSR[ 26 ][ 159 ],
   alphaCSR[ 26 ][ 160 ],
   alphaCSR[ 26 ][ 161 ],
   alphaCSR[ 26 ][ 162 ],
   alphaCSR[ 26 ][ 163 ],
   alphaCSR[ 26 ][ 164 ],
   alphaCSR[ 26 ][ 165 ],
   alphaCSR[ 26 ][ 166 ],
   alphaCSR[ 26 ][ 167 ],
   alphaCSR[ 26 ][ 168 ],
   alphaCSR[ 26 ][ 169 ],
   alphaCSR[ 26 ][ 170 ],
   alphaCSR[ 26 ][ 171 ],
   alphaCSR[ 26 ][ 172 ],
   alphaCSR[ 26 ][ 173 ],
   alphaCSR[ 26 ][ 174 ],
   alphaCSR[ 26 ][ 175 ],
   alphaCSR[ 26 ][ 176 ],
   alphaCSR[ 26 ][ 177 ],
   alphaCSR[ 26 ][ 178 ],
   alphaCSR[ 26 ][ 179 ],
   alphaCSR[ 26 ][ 180 ],
   alphaCSR[ 26 ][ 181 ],
   alphaCSR[ 26 ][ 182 ],
   alphaCSR[ 26 ][ 183 ],
   alphaCSR[ 26 ][ 184 ],
   alphaCSR[ 26 ][ 185 ],
   alphaCSR[ 26 ][ 186 ],
   alphaCSR[ 26 ][ 187 ],
   alphaCSR[ 26 ][ 188 ],
   alphaCSR[ 26 ][ 189 ],
   alphaCSR[ 26 ][ 190 ],
   alphaCSR[ 26 ][ 191 ],
   alphaCSR[ 26 ][ 192 ],
   alphaCSR[ 26 ][ 193 ],
   alphaCSR[ 26 ][ 194 ],
   alphaCSR[ 26 ][ 195 ],
   alphaCSR[ 26 ][ 196 ],
   alphaCSR[ 26 ][ 197 ],
   alphaCSR[ 26 ][ 198 ],
   alphaCSR[ 26 ][ 199 ],
   alphaCSR[ 26 ][ 200 ],
   alphaCSR[ 26 ][ 201 ],
   alphaCSR[ 26 ][ 202 ],
   alphaCSR[ 26 ][ 203 ],
   alphaCSR[ 26 ][ 204 ],
   alphaCSR[ 26 ][ 205 ],
   alphaCSR[ 26 ][ 206 ],
   alphaCSR[ 26 ][ 207 ],
   alphaCSR[ 26 ][ 208 ],
   alphaCSR[ 26 ][ 209 ],
   alphaCSR[ 26 ][ 210 ],
   alphaCSR[ 26 ][ 211 ],
   alphaCSR[ 26 ][ 212 ],
   alphaCSR[ 26 ][ 213 ],
   alphaCSR[ 26 ][ 214 ],
   alphaCSR[ 26 ][ 215 ],
   alphaCSR[ 26 ][ 216 ],
   alphaCSR[ 26 ][ 217 ],
   alphaCSR[ 26 ][ 218 ],
   alphaCSR[ 26 ][ 219 ],
   alphaCSR[ 26 ][ 220 ],
   alphaCSR[ 26 ][ 221 ],
   alphaCSR[ 26 ][ 222 ],
   alphaCSR[ 26 ][ 223 ],
   alphaCSR[ 26 ][ 224 ],
   alphaCSR[ 26 ][ 225 ],
   alphaCSR[ 26 ][ 226 ],
   alphaCSR[ 26 ][ 227 ],
   alphaCSR[ 26 ][ 228 ],
   alphaCSR[ 26 ][ 229 ],
   alphaCSR[ 26 ][ 230 ],
   alphaCSR[ 26 ][ 231 ],
   alphaCSR[ 26 ][ 232 ],
   alphaCSR[ 26 ][ 233 ],
   alphaCSR[ 26 ][ 234 ],
   alphaCSR[ 26 ][ 235 ],
   alphaCSR[ 26 ][ 236 ],
   alphaCSR[ 26 ][ 237 ],
   alphaCSR[ 26 ][ 238 ],
   alphaCSR[ 26 ][ 239 ],
   alphaCSR[ 26 ][ 240 ],
   alphaCSR[ 26 ][ 241 ],
   alphaCSR[ 26 ][ 242 ],
   alphaCSR[ 26 ][ 243 ],
   alphaCSR[ 26 ][ 244 ],
   alphaCSR[ 26 ][ 245 ],
   alphaCSR[ 26 ][ 246 ],
   alphaCSR[ 26 ][ 247 ],
   alphaCSR[ 26 ][ 248 ],
   alphaCSR[ 26 ][ 249 ],
   alphaCSR[ 26 ][ 250 ],
   alphaCSR[ 26 ][ 251 ],
   alphaCSR[ 26 ][ 252 ],
   alphaCSR[ 26 ][ 253 ],
   alphaCSR[ 26 ][ 254 ],
   alphaCSR[ 26 ][ 255 ],
   alphaCSR[ 26 ][ 256 ],
   alphaCSR[ 26 ][ 257 ],
   alphaCSR[ 26 ][ 258 ],
   alphaCSR[ 26 ][ 259 ],
   alphaCSR[ 26 ][ 260 ],
   alphaCSR[ 26 ][ 261 ],
   alphaCSR[ 26 ][ 262 ],
   alphaCSR[ 26 ][ 263 ],
   alphaCSR[ 26 ][ 264 ],
   alphaCSR[ 26 ][ 265 ],
   alphaCSR[ 26 ][ 266 ],
   alphaCSR[ 26 ][ 267 ],
   alphaCSR[ 26 ][ 268 ],
   alphaCSR[ 26 ][ 269 ],
   alphaCSR[ 26 ][ 270 ],
   alphaCSR[ 26 ][ 271 ],
   alphaCSR[ 26 ][ 272 ],
   alphaCSR[ 26 ][ 273 ],
   alphaCSR[ 26 ][ 274 ],
   alphaCSR[ 26 ][ 275 ],
   alphaCSR[ 26 ][ 276 ],
   alphaCSR[ 26 ][ 277 ],
   alphaCSR[ 26 ][ 278 ],
   alphaCSR[ 26 ][ 279 ],
   alphaCSR[ 26 ][ 280 ],
   alphaCSR[ 26 ][ 281 ],
   alphaCSR[ 26 ][ 282 ],
   alphaCSR[ 26 ][ 283 ],
   alphaCSR[ 26 ][ 284 ],
   alphaCSR[ 26 ][ 285 ],
   alphaCSR[ 26 ][ 286 ],
   alphaCSR[ 26 ][ 287 ],
   alphaCSR[ 26 ][ 288 ],
   alphaCSR[ 26 ][ 289 ],
   alphaCSR[ 26 ][ 290 ],
   alphaCSR[ 26 ][ 291 ],
   alphaCSR[ 26 ][ 292 ],
   alphaCSR[ 26 ][ 293 ],
   alphaCSR[ 26 ][ 294 ],
   alphaCSR[ 26 ][ 295 ],
   alphaCSR[ 26 ][ 296 ],
   alphaCSR[ 26 ][ 297 ],
   alphaCSR[ 26 ][ 298 ],
   alphaCSR[ 26 ][ 299 ],
   alphaCSR[ 26 ][ 300 ],
   alphaCSR[ 26 ][ 301 ],
   alphaCSR[ 26 ][ 302 ],
   alphaCSR[ 26 ][ 303 ],
   alphaCSR[ 26 ][ 304 ],
   alphaCSR[ 26 ][ 305 ],
   alphaCSR[ 26 ][ 306 ],
   alphaCSR[ 26 ][ 307 ],
   alphaCSR[ 26 ][ 308 ],
   alphaCSR[ 26 ][ 309 ],
   alphaCSR[ 26 ][ 310 ],
   alphaCSR[ 26 ][ 311 ],
   alphaCSR[ 26 ][ 312 ],
   alphaCSR[ 26 ][ 313 ],
   alphaCSR[ 26 ][ 314 ],
   alphaCSR[ 26 ][ 315 ],
   alphaCSR[ 26 ][ 316 ],
   alphaCSR[ 26 ][ 317 ],
   alphaCSR[ 26 ][ 318 ],
   alphaCSR[ 26 ][ 319 ],
   alphaCSR[ 26 ][ 320 ],
   alphaCSR[ 26 ][ 321 ],
   alphaCSR[ 26 ][ 322 ],
   alphaCSR[ 26 ][ 323 ],
   alphaCSR[ 26 ][ 324 ],
   alphaCSR[ 26 ][ 325 ],
   alphaCSR[ 26 ][ 326 ],
   alphaCSR[ 26 ][ 327 ],
   alphaCSR[ 26 ][ 328 ],
   alphaCSR[ 26 ][ 329 ],
   alphaCSR[ 26 ][ 330 ],
   alphaCSR[ 26 ][ 331 ],
   alphaCSR[ 26 ][ 332 ],
   alphaCSR[ 26 ][ 333 ],
   alphaCSR[ 26 ][ 334 ],
   alphaCSR[ 26 ][ 335 ],
   alphaCSR[ 26 ][ 336 ],
   alphaCSR[ 26 ][ 337 ],
   alphaCSR[ 26 ][ 338 ],
   alphaCSR[ 26 ][ 339 ],
   alphaCSR[ 26 ][ 340 ],
   alphaCSR[ 26 ][ 341 ],
   alphaCSR[ 26 ][ 342 ],
   alphaCSR[ 26 ][ 343 ],
   alphaCSR[ 26 ][ 344 ],
   alphaCSR[ 26 ][ 345 ],
   alphaCSR[ 26 ][ 346 ],
   alphaCSR[ 26 ][ 347 ],
   alphaCSR[ 26 ][ 348 ],
   alphaCSR[ 26 ][ 349 ],
   alphaCSR[ 26 ][ 350 ],
   alphaCSR[ 26 ][ 351 ],
   alphaCSR[ 26 ][ 352 ],
   alphaCSR[ 26 ][ 353 ],
   alphaCSR[ 26 ][ 354 ],
   alphaCSR[ 26 ][ 355 ],
   alphaCSR[ 26 ][ 356 ],
   alphaCSR[ 26 ][ 357 ],
   alphaCSR[ 26 ][ 358 ],
   alphaCSR[ 26 ][ 359 ],
   alphaCSR[ 26 ][ 360 ],
   alphaCSR[ 26 ][ 361 ],
   alphaCSR[ 26 ][ 362 ],
   alphaCSR[ 26 ][ 363 ],
   alphaCSR[ 26 ][ 364 ],
   alphaCSR[ 26 ][ 365 ],
   alphaCSR[ 26 ][ 366 ],
   alphaCSR[ 26 ][ 367 ],
   alphaCSR[ 26 ][ 368 ],
   alphaCSR[ 26 ][ 369 ],
   alphaCSR[ 26 ][ 370 ],
   alphaCSR[ 26 ][ 371 ],
   alphaCSR[ 26 ][ 372 ],
   alphaCSR[ 26 ][ 373 ],
   alphaCSR[ 26 ][ 374 ],
   alphaCSR[ 26 ][ 375 ],
   alphaCSR[ 26 ][ 376 ],
   alphaCSR[ 26 ][ 377 ],
   alphaCSR[ 26 ][ 378 ],
   alphaCSR[ 26 ][ 379 ],
   alphaCSR[ 26 ][ 380 ],
   alphaCSR[ 26 ][ 381 ],
   alphaCSR[ 26 ][ 382 ],
   alphaCSR[ 26 ][ 383 ],
   alphaCSR[ 27 ][ 0 ],
   alphaCSR[ 27 ][ 1 ],
   alphaCSR[ 27 ][ 2 ],
   alphaCSR[ 27 ][ 3 ],
   alphaCSR[ 27 ][ 4 ],
   alphaCSR[ 27 ][ 5 ],
   alphaCSR[ 27 ][ 6 ],
   alphaCSR[ 27 ][ 7 ],
   alphaCSR[ 27 ][ 8 ],
   alphaCSR[ 27 ][ 9 ],
   alphaCSR[ 27 ][ 10 ],
   alphaCSR[ 27 ][ 11 ],
   alphaCSR[ 27 ][ 12 ],
   alphaCSR[ 27 ][ 13 ],
   alphaCSR[ 27 ][ 14 ],
   alphaCSR[ 27 ][ 15 ],
   alphaCSR[ 27 ][ 16 ],
   alphaCSR[ 27 ][ 17 ],
   alphaCSR[ 27 ][ 18 ],
   alphaCSR[ 27 ][ 19 ],
   alphaCSR[ 27 ][ 20 ],
   alphaCSR[ 27 ][ 21 ],
   alphaCSR[ 27 ][ 22 ],
   alphaCSR[ 27 ][ 23 ],
   alphaCSR[ 27 ][ 24 ],
   alphaCSR[ 27 ][ 25 ],
   alphaCSR[ 27 ][ 26 ],
   alphaCSR[ 27 ][ 27 ],
   alphaCSR[ 27 ][ 28 ],
   alphaCSR[ 27 ][ 29 ],
   alphaCSR[ 27 ][ 30 ],
   alphaCSR[ 27 ][ 31 ],
   alphaCSR[ 27 ][ 32 ],
   alphaCSR[ 27 ][ 33 ],
   alphaCSR[ 27 ][ 34 ],
   alphaCSR[ 27 ][ 35 ],
   alphaCSR[ 27 ][ 36 ],
   alphaCSR[ 27 ][ 37 ],
   alphaCSR[ 27 ][ 38 ],
   alphaCSR[ 27 ][ 39 ],
   alphaCSR[ 27 ][ 40 ],
   alphaCSR[ 27 ][ 41 ],
   alphaCSR[ 27 ][ 42 ],
   alphaCSR[ 27 ][ 43 ],
   alphaCSR[ 27 ][ 44 ],
   alphaCSR[ 27 ][ 45 ],
   alphaCSR[ 27 ][ 46 ],
   alphaCSR[ 27 ][ 47 ],
   alphaCSR[ 27 ][ 48 ],
   alphaCSR[ 27 ][ 49 ],
   alphaCSR[ 27 ][ 50 ],
   alphaCSR[ 27 ][ 51 ],
   alphaCSR[ 27 ][ 52 ],
   alphaCSR[ 27 ][ 53 ],
   alphaCSR[ 27 ][ 54 ],
   alphaCSR[ 27 ][ 55 ],
   alphaCSR[ 27 ][ 56 ],
   alphaCSR[ 27 ][ 57 ],
   alphaCSR[ 27 ][ 58 ],
   alphaCSR[ 27 ][ 59 ],
   alphaCSR[ 27 ][ 60 ],
   alphaCSR[ 27 ][ 61 ],
   alphaCSR[ 27 ][ 62 ],
   alphaCSR[ 27 ][ 63 ],
   alphaCSR[ 27 ][ 64 ],
   alphaCSR[ 27 ][ 65 ],
   alphaCSR[ 27 ][ 66 ],
   alphaCSR[ 27 ][ 67 ],
   alphaCSR[ 27 ][ 68 ],
   alphaCSR[ 27 ][ 69 ],
   alphaCSR[ 27 ][ 70 ],
   alphaCSR[ 27 ][ 71 ],
   alphaCSR[ 27 ][ 72 ],
   alphaCSR[ 27 ][ 73 ],
   alphaCSR[ 27 ][ 74 ],
   alphaCSR[ 27 ][ 75 ],
   alphaCSR[ 27 ][ 76 ],
   alphaCSR[ 27 ][ 77 ],
   alphaCSR[ 27 ][ 78 ],
   alphaCSR[ 27 ][ 79 ],
   alphaCSR[ 27 ][ 80 ],
   alphaCSR[ 27 ][ 81 ],
   alphaCSR[ 27 ][ 82 ],
   alphaCSR[ 27 ][ 83 ],
   alphaCSR[ 27 ][ 84 ],
   alphaCSR[ 27 ][ 85 ],
   alphaCSR[ 27 ][ 86 ],
   alphaCSR[ 27 ][ 87 ],
   alphaCSR[ 27 ][ 88 ],
   alphaCSR[ 27 ][ 89 ],
   alphaCSR[ 27 ][ 90 ],
   alphaCSR[ 27 ][ 91 ],
   alphaCSR[ 27 ][ 92 ],
   alphaCSR[ 27 ][ 93 ],
   alphaCSR[ 27 ][ 94 ],
   alphaCSR[ 27 ][ 95 ],
   alphaCSR[ 27 ][ 96 ],
   alphaCSR[ 27 ][ 97 ],
   alphaCSR[ 27 ][ 98 ],
   alphaCSR[ 27 ][ 99 ],
   alphaCSR[ 27 ][ 100 ],
   alphaCSR[ 27 ][ 101 ],
   alphaCSR[ 27 ][ 102 ],
   alphaCSR[ 27 ][ 103 ],
   alphaCSR[ 27 ][ 104 ],
   alphaCSR[ 27 ][ 105 ],
   alphaCSR[ 27 ][ 106 ],
   alphaCSR[ 27 ][ 107 ],
   alphaCSR[ 27 ][ 108 ],
   alphaCSR[ 27 ][ 109 ],
   alphaCSR[ 27 ][ 110 ],
   alphaCSR[ 27 ][ 111 ],
   alphaCSR[ 27 ][ 112 ],
   alphaCSR[ 27 ][ 113 ],
   alphaCSR[ 27 ][ 114 ],
   alphaCSR[ 27 ][ 115 ],
   alphaCSR[ 27 ][ 116 ],
   alphaCSR[ 27 ][ 117 ],
   alphaCSR[ 27 ][ 118 ],
   alphaCSR[ 27 ][ 119 ],
   alphaCSR[ 27 ][ 120 ],
   alphaCSR[ 27 ][ 121 ],
   alphaCSR[ 27 ][ 122 ],
   alphaCSR[ 27 ][ 123 ],
   alphaCSR[ 27 ][ 124 ],
   alphaCSR[ 27 ][ 125 ],
   alphaCSR[ 27 ][ 126 ],
   alphaCSR[ 27 ][ 127 ],
   alphaCSR[ 27 ][ 128 ],
   alphaCSR[ 27 ][ 129 ],
   alphaCSR[ 27 ][ 130 ],
   alphaCSR[ 27 ][ 131 ],
   alphaCSR[ 27 ][ 132 ],
   alphaCSR[ 27 ][ 133 ],
   alphaCSR[ 27 ][ 134 ],
   alphaCSR[ 27 ][ 135 ],
   alphaCSR[ 27 ][ 136 ],
   alphaCSR[ 27 ][ 137 ],
   alphaCSR[ 27 ][ 138 ],
   alphaCSR[ 27 ][ 139 ],
   alphaCSR[ 27 ][ 140 ],
   alphaCSR[ 27 ][ 141 ],
   alphaCSR[ 27 ][ 142 ],
   alphaCSR[ 27 ][ 143 ],
   alphaCSR[ 27 ][ 144 ],
   alphaCSR[ 27 ][ 145 ],
   alphaCSR[ 27 ][ 146 ],
   alphaCSR[ 27 ][ 147 ],
   alphaCSR[ 27 ][ 148 ],
   alphaCSR[ 27 ][ 149 ],
   alphaCSR[ 27 ][ 150 ],
   alphaCSR[ 27 ][ 151 ],
   alphaCSR[ 27 ][ 152 ],
   alphaCSR[ 27 ][ 153 ],
   alphaCSR[ 27 ][ 154 ],
   alphaCSR[ 27 ][ 155 ],
   alphaCSR[ 27 ][ 156 ],
   alphaCSR[ 27 ][ 157 ],
   alphaCSR[ 27 ][ 158 ],
   alphaCSR[ 27 ][ 159 ],
   alphaCSR[ 27 ][ 160 ],
   alphaCSR[ 27 ][ 161 ],
   alphaCSR[ 27 ][ 162 ],
   alphaCSR[ 27 ][ 163 ],
   alphaCSR[ 27 ][ 164 ],
   alphaCSR[ 27 ][ 165 ],
   alphaCSR[ 27 ][ 166 ],
   alphaCSR[ 27 ][ 167 ],
   alphaCSR[ 27 ][ 168 ],
   alphaCSR[ 27 ][ 169 ],
   alphaCSR[ 27 ][ 170 ],
   alphaCSR[ 27 ][ 171 ],
   alphaCSR[ 27 ][ 172 ],
   alphaCSR[ 27 ][ 173 ],
   alphaCSR[ 27 ][ 174 ],
   alphaCSR[ 27 ][ 175 ],
   alphaCSR[ 27 ][ 176 ],
   alphaCSR[ 27 ][ 177 ],
   alphaCSR[ 27 ][ 178 ],
   alphaCSR[ 27 ][ 179 ],
   alphaCSR[ 27 ][ 180 ],
   alphaCSR[ 27 ][ 181 ],
   alphaCSR[ 27 ][ 182 ],
   alphaCSR[ 27 ][ 183 ],
   alphaCSR[ 27 ][ 184 ],
   alphaCSR[ 27 ][ 185 ],
   alphaCSR[ 27 ][ 186 ],
   alphaCSR[ 27 ][ 187 ],
   alphaCSR[ 27 ][ 188 ],
   alphaCSR[ 27 ][ 189 ],
   alphaCSR[ 27 ][ 190 ],
   alphaCSR[ 27 ][ 191 ],
   alphaCSR[ 27 ][ 192 ],
   alphaCSR[ 27 ][ 193 ],
   alphaCSR[ 27 ][ 194 ],
   alphaCSR[ 27 ][ 195 ],
   alphaCSR[ 27 ][ 196 ],
   alphaCSR[ 27 ][ 197 ],
   alphaCSR[ 27 ][ 198 ],
   alphaCSR[ 27 ][ 199 ],
   alphaCSR[ 27 ][ 200 ],
   alphaCSR[ 27 ][ 201 ],
   alphaCSR[ 27 ][ 202 ],
   alphaCSR[ 27 ][ 203 ],
   alphaCSR[ 27 ][ 204 ],
   alphaCSR[ 27 ][ 205 ],
   alphaCSR[ 27 ][ 206 ],
   alphaCSR[ 27 ][ 207 ],
   alphaCSR[ 27 ][ 208 ],
   alphaCSR[ 27 ][ 209 ],
   alphaCSR[ 27 ][ 210 ],
   alphaCSR[ 27 ][ 211 ],
   alphaCSR[ 27 ][ 212 ],
   alphaCSR[ 27 ][ 213 ],
   alphaCSR[ 27 ][ 214 ],
   alphaCSR[ 27 ][ 215 ],
   alphaCSR[ 27 ][ 216 ],
   alphaCSR[ 27 ][ 217 ],
   alphaCSR[ 27 ][ 218 ],
   alphaCSR[ 27 ][ 219 ],
   alphaCSR[ 27 ][ 220 ],
   alphaCSR[ 27 ][ 221 ],
   alphaCSR[ 27 ][ 222 ],
   alphaCSR[ 27 ][ 223 ],
   alphaCSR[ 27 ][ 224 ],
   alphaCSR[ 27 ][ 225 ],
   alphaCSR[ 27 ][ 226 ],
   alphaCSR[ 27 ][ 227 ],
   alphaCSR[ 27 ][ 228 ],
   alphaCSR[ 27 ][ 229 ],
   alphaCSR[ 27 ][ 230 ],
   alphaCSR[ 27 ][ 231 ],
   alphaCSR[ 27 ][ 232 ],
   alphaCSR[ 27 ][ 233 ],
   alphaCSR[ 27 ][ 234 ],
   alphaCSR[ 27 ][ 235 ],
   alphaCSR[ 27 ][ 236 ],
   alphaCSR[ 27 ][ 237 ],
   alphaCSR[ 27 ][ 238 ],
   alphaCSR[ 27 ][ 239 ],
   alphaCSR[ 27 ][ 240 ],
   alphaCSR[ 27 ][ 241 ],
   alphaCSR[ 27 ][ 242 ],
   alphaCSR[ 27 ][ 243 ],
   alphaCSR[ 27 ][ 244 ],
   alphaCSR[ 27 ][ 245 ],
   alphaCSR[ 27 ][ 246 ],
   alphaCSR[ 27 ][ 247 ],
   alphaCSR[ 27 ][ 248 ],
   alphaCSR[ 27 ][ 249 ],
   alphaCSR[ 27 ][ 250 ],
   alphaCSR[ 27 ][ 251 ],
   alphaCSR[ 27 ][ 252 ],
   alphaCSR[ 27 ][ 253 ],
   alphaCSR[ 27 ][ 254 ],
   alphaCSR[ 27 ][ 255 ],
   alphaCSR[ 27 ][ 256 ],
   alphaCSR[ 27 ][ 257 ],
   alphaCSR[ 27 ][ 258 ],
   alphaCSR[ 27 ][ 259 ],
   alphaCSR[ 27 ][ 260 ],
   alphaCSR[ 27 ][ 261 ],
   alphaCSR[ 27 ][ 262 ],
   alphaCSR[ 27 ][ 263 ],
   alphaCSR[ 27 ][ 264 ],
   alphaCSR[ 27 ][ 265 ],
   alphaCSR[ 27 ][ 266 ],
   alphaCSR[ 27 ][ 267 ],
   alphaCSR[ 27 ][ 268 ],
   alphaCSR[ 27 ][ 269 ],
   alphaCSR[ 27 ][ 270 ],
   alphaCSR[ 27 ][ 271 ],
   alphaCSR[ 27 ][ 272 ],
   alphaCSR[ 27 ][ 273 ],
   alphaCSR[ 27 ][ 274 ],
   alphaCSR[ 27 ][ 275 ],
   alphaCSR[ 27 ][ 276 ],
   alphaCSR[ 27 ][ 277 ],
   alphaCSR[ 27 ][ 278 ],
   alphaCSR[ 27 ][ 279 ],
   alphaCSR[ 27 ][ 280 ],
   alphaCSR[ 27 ][ 281 ],
   alphaCSR[ 27 ][ 282 ],
   alphaCSR[ 27 ][ 283 ],
   alphaCSR[ 27 ][ 284 ],
   alphaCSR[ 27 ][ 285 ],
   alphaCSR[ 27 ][ 286 ],
   alphaCSR[ 27 ][ 287 ],
   alphaCSR[ 27 ][ 288 ],
   alphaCSR[ 27 ][ 289 ],
   alphaCSR[ 27 ][ 290 ],
   alphaCSR[ 27 ][ 291 ],
   alphaCSR[ 27 ][ 292 ],
   alphaCSR[ 27 ][ 293 ],
   alphaCSR[ 27 ][ 294 ],
   alphaCSR[ 27 ][ 295 ],
   alphaCSR[ 27 ][ 296 ],
   alphaCSR[ 27 ][ 297 ],
   alphaCSR[ 27 ][ 298 ],
   alphaCSR[ 27 ][ 299 ],
   alphaCSR[ 27 ][ 300 ],
   alphaCSR[ 27 ][ 301 ],
   alphaCSR[ 27 ][ 302 ],
   alphaCSR[ 27 ][ 303 ],
   alphaCSR[ 27 ][ 304 ],
   alphaCSR[ 27 ][ 305 ],
   alphaCSR[ 27 ][ 306 ],
   alphaCSR[ 27 ][ 307 ],
   alphaCSR[ 27 ][ 308 ],
   alphaCSR[ 27 ][ 309 ],
   alphaCSR[ 27 ][ 310 ],
   alphaCSR[ 27 ][ 311 ],
   alphaCSR[ 27 ][ 312 ],
   alphaCSR[ 27 ][ 313 ],
   alphaCSR[ 27 ][ 314 ],
   alphaCSR[ 27 ][ 315 ],
   alphaCSR[ 27 ][ 316 ],
   alphaCSR[ 27 ][ 317 ],
   alphaCSR[ 27 ][ 318 ],
   alphaCSR[ 27 ][ 319 ],
   alphaCSR[ 27 ][ 320 ],
   alphaCSR[ 27 ][ 321 ],
   alphaCSR[ 27 ][ 322 ],
   alphaCSR[ 27 ][ 323 ],
   alphaCSR[ 27 ][ 324 ],
   alphaCSR[ 27 ][ 325 ],
   alphaCSR[ 27 ][ 326 ],
   alphaCSR[ 27 ][ 327 ],
   alphaCSR[ 27 ][ 328 ],
   alphaCSR[ 27 ][ 329 ],
   alphaCSR[ 27 ][ 330 ],
   alphaCSR[ 27 ][ 331 ],
   alphaCSR[ 27 ][ 332 ],
   alphaCSR[ 27 ][ 333 ],
   alphaCSR[ 27 ][ 334 ],
   alphaCSR[ 27 ][ 335 ],
   alphaCSR[ 27 ][ 336 ],
   alphaCSR[ 27 ][ 337 ],
   alphaCSR[ 27 ][ 338 ],
   alphaCSR[ 27 ][ 339 ],
   alphaCSR[ 27 ][ 340 ],
   alphaCSR[ 27 ][ 341 ],
   alphaCSR[ 27 ][ 342 ],
   alphaCSR[ 27 ][ 343 ],
   alphaCSR[ 27 ][ 344 ],
   alphaCSR[ 27 ][ 345 ],
   alphaCSR[ 27 ][ 346 ],
   alphaCSR[ 27 ][ 347 ],
   alphaCSR[ 27 ][ 348 ],
   alphaCSR[ 27 ][ 349 ],
   alphaCSR[ 27 ][ 350 ],
   alphaCSR[ 27 ][ 351 ],
   alphaCSR[ 27 ][ 352 ],
   alphaCSR[ 27 ][ 353 ],
   alphaCSR[ 27 ][ 354 ],
   alphaCSR[ 27 ][ 355 ],
   alphaCSR[ 27 ][ 356 ],
   alphaCSR[ 27 ][ 357 ],
   alphaCSR[ 27 ][ 358 ],
   alphaCSR[ 27 ][ 359 ],
   alphaCSR[ 27 ][ 360 ],
   alphaCSR[ 27 ][ 361 ],
   alphaCSR[ 27 ][ 362 ],
   alphaCSR[ 27 ][ 363 ],
   alphaCSR[ 27 ][ 364 ],
   alphaCSR[ 27 ][ 365 ],
   alphaCSR[ 27 ][ 366 ],
   alphaCSR[ 27 ][ 367 ],
   alphaCSR[ 27 ][ 368 ],
   alphaCSR[ 27 ][ 369 ],
   alphaCSR[ 27 ][ 370 ],
   alphaCSR[ 27 ][ 371 ],
   alphaCSR[ 27 ][ 372 ],
   alphaCSR[ 27 ][ 373 ],
   alphaCSR[ 27 ][ 374 ],
   alphaCSR[ 27 ][ 375 ],
   alphaCSR[ 27 ][ 376 ],
   alphaCSR[ 27 ][ 377 ],
   alphaCSR[ 27 ][ 378 ],
   alphaCSR[ 27 ][ 379 ],
   alphaCSR[ 27 ][ 380 ],
   alphaCSR[ 27 ][ 381 ],
   alphaCSR[ 27 ][ 382 ],
   alphaCSR[ 27 ][ 383 ],
   alphaCSR[ 28 ][ 0 ],
   alphaCSR[ 28 ][ 1 ],
   alphaCSR[ 28 ][ 2 ],
   alphaCSR[ 28 ][ 3 ],
   alphaCSR[ 28 ][ 4 ],
   alphaCSR[ 28 ][ 5 ],
   alphaCSR[ 28 ][ 6 ],
   alphaCSR[ 28 ][ 7 ],
   alphaCSR[ 28 ][ 8 ],
   alphaCSR[ 28 ][ 9 ],
   alphaCSR[ 28 ][ 10 ],
   alphaCSR[ 28 ][ 11 ],
   alphaCSR[ 28 ][ 12 ],
   alphaCSR[ 28 ][ 13 ],
   alphaCSR[ 28 ][ 14 ],
   alphaCSR[ 28 ][ 15 ],
   alphaCSR[ 28 ][ 16 ],
   alphaCSR[ 28 ][ 17 ],
   alphaCSR[ 28 ][ 18 ],
   alphaCSR[ 28 ][ 19 ],
   alphaCSR[ 28 ][ 20 ],
   alphaCSR[ 28 ][ 21 ],
   alphaCSR[ 28 ][ 22 ],
   alphaCSR[ 28 ][ 23 ],
   alphaCSR[ 28 ][ 24 ],
   alphaCSR[ 28 ][ 25 ],
   alphaCSR[ 28 ][ 26 ],
   alphaCSR[ 28 ][ 27 ],
   alphaCSR[ 28 ][ 28 ],
   alphaCSR[ 28 ][ 29 ],
   alphaCSR[ 28 ][ 30 ],
   alphaCSR[ 28 ][ 31 ],
   alphaCSR[ 28 ][ 32 ],
   alphaCSR[ 28 ][ 33 ],
   alphaCSR[ 28 ][ 34 ],
   alphaCSR[ 28 ][ 35 ],
   alphaCSR[ 28 ][ 36 ],
   alphaCSR[ 28 ][ 37 ],
   alphaCSR[ 28 ][ 38 ],
   alphaCSR[ 28 ][ 39 ],
   alphaCSR[ 28 ][ 40 ],
   alphaCSR[ 28 ][ 41 ],
   alphaCSR[ 28 ][ 42 ],
   alphaCSR[ 28 ][ 43 ],
   alphaCSR[ 28 ][ 44 ],
   alphaCSR[ 28 ][ 45 ],
   alphaCSR[ 28 ][ 46 ],
   alphaCSR[ 28 ][ 47 ],
   alphaCSR[ 28 ][ 48 ],
   alphaCSR[ 28 ][ 49 ],
   alphaCSR[ 28 ][ 50 ],
   alphaCSR[ 28 ][ 51 ],
   alphaCSR[ 28 ][ 52 ],
   alphaCSR[ 28 ][ 53 ],
   alphaCSR[ 28 ][ 54 ],
   alphaCSR[ 28 ][ 55 ],
   alphaCSR[ 28 ][ 56 ],
   alphaCSR[ 28 ][ 57 ],
   alphaCSR[ 28 ][ 58 ],
   alphaCSR[ 28 ][ 59 ],
   alphaCSR[ 28 ][ 60 ],
   alphaCSR[ 28 ][ 61 ],
   alphaCSR[ 28 ][ 62 ],
   alphaCSR[ 28 ][ 63 ],
   alphaCSR[ 28 ][ 64 ],
   alphaCSR[ 28 ][ 65 ],
   alphaCSR[ 28 ][ 66 ],
   alphaCSR[ 28 ][ 67 ],
   alphaCSR[ 28 ][ 68 ],
   alphaCSR[ 28 ][ 69 ],
   alphaCSR[ 28 ][ 70 ],
   alphaCSR[ 28 ][ 71 ],
   alphaCSR[ 28 ][ 72 ],
   alphaCSR[ 28 ][ 73 ],
   alphaCSR[ 28 ][ 74 ],
   alphaCSR[ 28 ][ 75 ],
   alphaCSR[ 28 ][ 76 ],
   alphaCSR[ 28 ][ 77 ],
   alphaCSR[ 28 ][ 78 ],
   alphaCSR[ 28 ][ 79 ],
   alphaCSR[ 28 ][ 80 ],
   alphaCSR[ 28 ][ 81 ],
   alphaCSR[ 28 ][ 82 ],
   alphaCSR[ 28 ][ 83 ],
   alphaCSR[ 28 ][ 84 ],
   alphaCSR[ 28 ][ 85 ],
   alphaCSR[ 28 ][ 86 ],
   alphaCSR[ 28 ][ 87 ],
   alphaCSR[ 28 ][ 88 ],
   alphaCSR[ 28 ][ 89 ],
   alphaCSR[ 28 ][ 90 ],
   alphaCSR[ 28 ][ 91 ],
   alphaCSR[ 28 ][ 92 ],
   alphaCSR[ 28 ][ 93 ],
   alphaCSR[ 28 ][ 94 ],
   alphaCSR[ 28 ][ 95 ],
   alphaCSR[ 28 ][ 96 ],
   alphaCSR[ 28 ][ 97 ],
   alphaCSR[ 28 ][ 98 ],
   alphaCSR[ 28 ][ 99 ],
   alphaCSR[ 28 ][ 100 ],
   alphaCSR[ 28 ][ 101 ],
   alphaCSR[ 28 ][ 102 ],
   alphaCSR[ 28 ][ 103 ],
   alphaCSR[ 28 ][ 104 ],
   alphaCSR[ 28 ][ 105 ],
   alphaCSR[ 28 ][ 106 ],
   alphaCSR[ 28 ][ 107 ],
   alphaCSR[ 28 ][ 108 ],
   alphaCSR[ 28 ][ 109 ],
   alphaCSR[ 28 ][ 110 ],
   alphaCSR[ 28 ][ 111 ],
   alphaCSR[ 28 ][ 112 ],
   alphaCSR[ 28 ][ 113 ],
   alphaCSR[ 28 ][ 114 ],
   alphaCSR[ 28 ][ 115 ],
   alphaCSR[ 28 ][ 116 ],
   alphaCSR[ 28 ][ 117 ],
   alphaCSR[ 28 ][ 118 ],
   alphaCSR[ 28 ][ 119 ],
   alphaCSR[ 28 ][ 120 ],
   alphaCSR[ 28 ][ 121 ],
   alphaCSR[ 28 ][ 122 ],
   alphaCSR[ 28 ][ 123 ],
   alphaCSR[ 28 ][ 124 ],
   alphaCSR[ 28 ][ 125 ],
   alphaCSR[ 28 ][ 126 ],
   alphaCSR[ 28 ][ 127 ],
   alphaCSR[ 28 ][ 128 ],
   alphaCSR[ 28 ][ 129 ],
   alphaCSR[ 28 ][ 130 ],
   alphaCSR[ 28 ][ 131 ],
   alphaCSR[ 28 ][ 132 ],
   alphaCSR[ 28 ][ 133 ],
   alphaCSR[ 28 ][ 134 ],
   alphaCSR[ 28 ][ 135 ],
   alphaCSR[ 28 ][ 136 ],
   alphaCSR[ 28 ][ 137 ],
   alphaCSR[ 28 ][ 138 ],
   alphaCSR[ 28 ][ 139 ],
   alphaCSR[ 28 ][ 140 ],
   alphaCSR[ 28 ][ 141 ],
   alphaCSR[ 28 ][ 142 ],
   alphaCSR[ 28 ][ 143 ],
   alphaCSR[ 28 ][ 144 ],
   alphaCSR[ 28 ][ 145 ],
   alphaCSR[ 28 ][ 146 ],
   alphaCSR[ 28 ][ 147 ],
   alphaCSR[ 28 ][ 148 ],
   alphaCSR[ 28 ][ 149 ],
   alphaCSR[ 28 ][ 150 ],
   alphaCSR[ 28 ][ 151 ],
   alphaCSR[ 28 ][ 152 ],
   alphaCSR[ 28 ][ 153 ],
   alphaCSR[ 28 ][ 154 ],
   alphaCSR[ 28 ][ 155 ],
   alphaCSR[ 28 ][ 156 ],
   alphaCSR[ 28 ][ 157 ],
   alphaCSR[ 28 ][ 158 ],
   alphaCSR[ 28 ][ 159 ],
   alphaCSR[ 28 ][ 160 ],
   alphaCSR[ 28 ][ 161 ],
   alphaCSR[ 28 ][ 162 ],
   alphaCSR[ 28 ][ 163 ],
   alphaCSR[ 28 ][ 164 ],
   alphaCSR[ 28 ][ 165 ],
   alphaCSR[ 28 ][ 166 ],
   alphaCSR[ 28 ][ 167 ],
   alphaCSR[ 28 ][ 168 ],
   alphaCSR[ 28 ][ 169 ],
   alphaCSR[ 28 ][ 170 ],
   alphaCSR[ 28 ][ 171 ],
   alphaCSR[ 28 ][ 172 ],
   alphaCSR[ 28 ][ 173 ],
   alphaCSR[ 28 ][ 174 ],
   alphaCSR[ 28 ][ 175 ],
   alphaCSR[ 28 ][ 176 ],
   alphaCSR[ 28 ][ 177 ],
   alphaCSR[ 28 ][ 178 ],
   alphaCSR[ 28 ][ 179 ],
   alphaCSR[ 28 ][ 180 ],
   alphaCSR[ 28 ][ 181 ],
   alphaCSR[ 28 ][ 182 ],
   alphaCSR[ 28 ][ 183 ],
   alphaCSR[ 28 ][ 184 ],
   alphaCSR[ 28 ][ 185 ],
   alphaCSR[ 28 ][ 186 ],
   alphaCSR[ 28 ][ 187 ],
   alphaCSR[ 28 ][ 188 ],
   alphaCSR[ 28 ][ 189 ],
   alphaCSR[ 28 ][ 190 ],
   alphaCSR[ 28 ][ 191 ],
   alphaCSR[ 28 ][ 192 ],
   alphaCSR[ 28 ][ 193 ],
   alphaCSR[ 28 ][ 194 ],
   alphaCSR[ 28 ][ 195 ],
   alphaCSR[ 28 ][ 196 ],
   alphaCSR[ 28 ][ 197 ],
   alphaCSR[ 28 ][ 198 ],
   alphaCSR[ 28 ][ 199 ],
   alphaCSR[ 28 ][ 200 ],
   alphaCSR[ 28 ][ 201 ],
   alphaCSR[ 28 ][ 202 ],
   alphaCSR[ 28 ][ 203 ],
   alphaCSR[ 28 ][ 204 ],
   alphaCSR[ 28 ][ 205 ],
   alphaCSR[ 28 ][ 206 ],
   alphaCSR[ 28 ][ 207 ],
   alphaCSR[ 28 ][ 208 ],
   alphaCSR[ 28 ][ 209 ],
   alphaCSR[ 28 ][ 210 ],
   alphaCSR[ 28 ][ 211 ],
   alphaCSR[ 28 ][ 212 ],
   alphaCSR[ 28 ][ 213 ],
   alphaCSR[ 28 ][ 214 ],
   alphaCSR[ 28 ][ 215 ],
   alphaCSR[ 28 ][ 216 ],
   alphaCSR[ 28 ][ 217 ],
   alphaCSR[ 28 ][ 218 ],
   alphaCSR[ 28 ][ 219 ],
   alphaCSR[ 28 ][ 220 ],
   alphaCSR[ 28 ][ 221 ],
   alphaCSR[ 28 ][ 222 ],
   alphaCSR[ 28 ][ 223 ],
   alphaCSR[ 28 ][ 224 ],
   alphaCSR[ 28 ][ 225 ],
   alphaCSR[ 28 ][ 226 ],
   alphaCSR[ 28 ][ 227 ],
   alphaCSR[ 28 ][ 228 ],
   alphaCSR[ 28 ][ 229 ],
   alphaCSR[ 28 ][ 230 ],
   alphaCSR[ 28 ][ 231 ],
   alphaCSR[ 28 ][ 232 ],
   alphaCSR[ 28 ][ 233 ],
   alphaCSR[ 28 ][ 234 ],
   alphaCSR[ 28 ][ 235 ],
   alphaCSR[ 28 ][ 236 ],
   alphaCSR[ 28 ][ 237 ],
   alphaCSR[ 28 ][ 238 ],
   alphaCSR[ 28 ][ 239 ],
   alphaCSR[ 28 ][ 240 ],
   alphaCSR[ 28 ][ 241 ],
   alphaCSR[ 28 ][ 242 ],
   alphaCSR[ 28 ][ 243 ],
   alphaCSR[ 28 ][ 244 ],
   alphaCSR[ 28 ][ 245 ],
   alphaCSR[ 28 ][ 246 ],
   alphaCSR[ 28 ][ 247 ],
   alphaCSR[ 28 ][ 248 ],
   alphaCSR[ 28 ][ 249 ],
   alphaCSR[ 28 ][ 250 ],
   alphaCSR[ 28 ][ 251 ],
   alphaCSR[ 28 ][ 252 ],
   alphaCSR[ 28 ][ 253 ],
   alphaCSR[ 28 ][ 254 ],
   alphaCSR[ 28 ][ 255 ],
   alphaCSR[ 28 ][ 256 ],
   alphaCSR[ 28 ][ 257 ],
   alphaCSR[ 28 ][ 258 ],
   alphaCSR[ 28 ][ 259 ],
   alphaCSR[ 28 ][ 260 ],
   alphaCSR[ 28 ][ 261 ],
   alphaCSR[ 28 ][ 262 ],
   alphaCSR[ 28 ][ 263 ],
   alphaCSR[ 28 ][ 264 ],
   alphaCSR[ 28 ][ 265 ],
   alphaCSR[ 28 ][ 266 ],
   alphaCSR[ 28 ][ 267 ],
   alphaCSR[ 28 ][ 268 ],
   alphaCSR[ 28 ][ 269 ],
   alphaCSR[ 28 ][ 270 ],
   alphaCSR[ 28 ][ 271 ],
   alphaCSR[ 28 ][ 272 ],
   alphaCSR[ 28 ][ 273 ],
   alphaCSR[ 28 ][ 274 ],
   alphaCSR[ 28 ][ 275 ],
   alphaCSR[ 28 ][ 276 ],
   alphaCSR[ 28 ][ 277 ],
   alphaCSR[ 28 ][ 278 ],
   alphaCSR[ 28 ][ 279 ],
   alphaCSR[ 28 ][ 280 ],
   alphaCSR[ 28 ][ 281 ],
   alphaCSR[ 28 ][ 282 ],
   alphaCSR[ 28 ][ 283 ],
   alphaCSR[ 28 ][ 284 ],
   alphaCSR[ 28 ][ 285 ],
   alphaCSR[ 28 ][ 286 ],
   alphaCSR[ 28 ][ 287 ],
   alphaCSR[ 28 ][ 288 ],
   alphaCSR[ 28 ][ 289 ],
   alphaCSR[ 28 ][ 290 ],
   alphaCSR[ 28 ][ 291 ],
   alphaCSR[ 28 ][ 292 ],
   alphaCSR[ 28 ][ 293 ],
   alphaCSR[ 28 ][ 294 ],
   alphaCSR[ 28 ][ 295 ],
   alphaCSR[ 28 ][ 296 ],
   alphaCSR[ 28 ][ 297 ],
   alphaCSR[ 28 ][ 298 ],
   alphaCSR[ 28 ][ 299 ],
   alphaCSR[ 28 ][ 300 ],
   alphaCSR[ 28 ][ 301 ],
   alphaCSR[ 28 ][ 302 ],
   alphaCSR[ 28 ][ 303 ],
   alphaCSR[ 28 ][ 304 ],
   alphaCSR[ 28 ][ 305 ],
   alphaCSR[ 28 ][ 306 ],
   alphaCSR[ 28 ][ 307 ],
   alphaCSR[ 28 ][ 308 ],
   alphaCSR[ 28 ][ 309 ],
   alphaCSR[ 28 ][ 310 ],
   alphaCSR[ 28 ][ 311 ],
   alphaCSR[ 28 ][ 312 ],
   alphaCSR[ 28 ][ 313 ],
   alphaCSR[ 28 ][ 314 ],
   alphaCSR[ 28 ][ 315 ],
   alphaCSR[ 28 ][ 316 ],
   alphaCSR[ 28 ][ 317 ],
   alphaCSR[ 28 ][ 318 ],
   alphaCSR[ 28 ][ 319 ],
   alphaCSR[ 28 ][ 320 ],
   alphaCSR[ 28 ][ 321 ],
   alphaCSR[ 28 ][ 322 ],
   alphaCSR[ 28 ][ 323 ],
   alphaCSR[ 28 ][ 324 ],
   alphaCSR[ 28 ][ 325 ],
   alphaCSR[ 28 ][ 326 ],
   alphaCSR[ 28 ][ 327 ],
   alphaCSR[ 28 ][ 328 ],
   alphaCSR[ 28 ][ 329 ],
   alphaCSR[ 28 ][ 330 ],
   alphaCSR[ 28 ][ 331 ],
   alphaCSR[ 28 ][ 332 ],
   alphaCSR[ 28 ][ 333 ],
   alphaCSR[ 28 ][ 334 ],
   alphaCSR[ 28 ][ 335 ],
   alphaCSR[ 28 ][ 336 ],
   alphaCSR[ 28 ][ 337 ],
   alphaCSR[ 28 ][ 338 ],
   alphaCSR[ 28 ][ 339 ],
   alphaCSR[ 28 ][ 340 ],
   alphaCSR[ 28 ][ 341 ],
   alphaCSR[ 28 ][ 342 ],
   alphaCSR[ 28 ][ 343 ],
   alphaCSR[ 28 ][ 344 ],
   alphaCSR[ 28 ][ 345 ],
   alphaCSR[ 28 ][ 346 ],
   alphaCSR[ 28 ][ 347 ],
   alphaCSR[ 28 ][ 348 ],
   alphaCSR[ 28 ][ 349 ],
   alphaCSR[ 28 ][ 350 ],
   alphaCSR[ 28 ][ 351 ],
   alphaCSR[ 28 ][ 352 ],
   alphaCSR[ 28 ][ 353 ],
   alphaCSR[ 28 ][ 354 ],
   alphaCSR[ 28 ][ 355 ],
   alphaCSR[ 28 ][ 356 ],
   alphaCSR[ 28 ][ 357 ],
   alphaCSR[ 28 ][ 358 ],
   alphaCSR[ 28 ][ 359 ],
   alphaCSR[ 28 ][ 360 ],
   alphaCSR[ 28 ][ 361 ],
   alphaCSR[ 28 ][ 362 ],
   alphaCSR[ 28 ][ 363 ],
   alphaCSR[ 28 ][ 364 ],
   alphaCSR[ 28 ][ 365 ],
   alphaCSR[ 28 ][ 366 ],
   alphaCSR[ 28 ][ 367 ],
   alphaCSR[ 28 ][ 368 ],
   alphaCSR[ 28 ][ 369 ],
   alphaCSR[ 28 ][ 370 ],
   alphaCSR[ 28 ][ 371 ],
   alphaCSR[ 28 ][ 372 ],
   alphaCSR[ 28 ][ 373 ],
   alphaCSR[ 28 ][ 374 ],
   alphaCSR[ 28 ][ 375 ],
   alphaCSR[ 28 ][ 376 ],
   alphaCSR[ 28 ][ 377 ],
   alphaCSR[ 28 ][ 378 ],
   alphaCSR[ 28 ][ 379 ],
   alphaCSR[ 28 ][ 380 ],
   alphaCSR[ 28 ][ 381 ],
   alphaCSR[ 28 ][ 382 ],
   alphaCSR[ 28 ][ 383 ],
   alphaCSR[ 29 ][ 0 ],
   alphaCSR[ 29 ][ 1 ],
   alphaCSR[ 29 ][ 2 ],
   alphaCSR[ 29 ][ 3 ],
   alphaCSR[ 29 ][ 4 ],
   alphaCSR[ 29 ][ 5 ],
   alphaCSR[ 29 ][ 6 ],
   alphaCSR[ 29 ][ 7 ],
   alphaCSR[ 29 ][ 8 ],
   alphaCSR[ 29 ][ 9 ],
   alphaCSR[ 29 ][ 10 ],
   alphaCSR[ 29 ][ 11 ],
   alphaCSR[ 29 ][ 12 ],
   alphaCSR[ 29 ][ 13 ],
   alphaCSR[ 29 ][ 14 ],
   alphaCSR[ 29 ][ 15 ],
   alphaCSR[ 29 ][ 16 ],
   alphaCSR[ 29 ][ 17 ],
   alphaCSR[ 29 ][ 18 ],
   alphaCSR[ 29 ][ 19 ],
   alphaCSR[ 29 ][ 20 ],
   alphaCSR[ 29 ][ 21 ],
   alphaCSR[ 29 ][ 22 ],
   alphaCSR[ 29 ][ 23 ],
   alphaCSR[ 29 ][ 24 ],
   alphaCSR[ 29 ][ 25 ],
   alphaCSR[ 29 ][ 26 ],
   alphaCSR[ 29 ][ 27 ],
   alphaCSR[ 29 ][ 28 ],
   alphaCSR[ 29 ][ 29 ],
   alphaCSR[ 29 ][ 30 ],
   alphaCSR[ 29 ][ 31 ],
   alphaCSR[ 29 ][ 32 ],
   alphaCSR[ 29 ][ 33 ],
   alphaCSR[ 29 ][ 34 ],
   alphaCSR[ 29 ][ 35 ],
   alphaCSR[ 29 ][ 36 ],
   alphaCSR[ 29 ][ 37 ],
   alphaCSR[ 29 ][ 38 ],
   alphaCSR[ 29 ][ 39 ],
   alphaCSR[ 29 ][ 40 ],
   alphaCSR[ 29 ][ 41 ],
   alphaCSR[ 29 ][ 42 ],
   alphaCSR[ 29 ][ 43 ],
   alphaCSR[ 29 ][ 44 ],
   alphaCSR[ 29 ][ 45 ],
   alphaCSR[ 29 ][ 46 ],
   alphaCSR[ 29 ][ 47 ],
   alphaCSR[ 29 ][ 48 ],
   alphaCSR[ 29 ][ 49 ],
   alphaCSR[ 29 ][ 50 ],
   alphaCSR[ 29 ][ 51 ],
   alphaCSR[ 29 ][ 52 ],
   alphaCSR[ 29 ][ 53 ],
   alphaCSR[ 29 ][ 54 ],
   alphaCSR[ 29 ][ 55 ],
   alphaCSR[ 29 ][ 56 ],
   alphaCSR[ 29 ][ 57 ],
   alphaCSR[ 29 ][ 58 ],
   alphaCSR[ 29 ][ 59 ],
   alphaCSR[ 29 ][ 60 ],
   alphaCSR[ 29 ][ 61 ],
   alphaCSR[ 29 ][ 62 ],
   alphaCSR[ 29 ][ 63 ],
   alphaCSR[ 29 ][ 64 ],
   alphaCSR[ 29 ][ 65 ],
   alphaCSR[ 29 ][ 66 ],
   alphaCSR[ 29 ][ 67 ],
   alphaCSR[ 29 ][ 68 ],
   alphaCSR[ 29 ][ 69 ],
   alphaCSR[ 29 ][ 70 ],
   alphaCSR[ 29 ][ 71 ],
   alphaCSR[ 29 ][ 72 ],
   alphaCSR[ 29 ][ 73 ],
   alphaCSR[ 29 ][ 74 ],
   alphaCSR[ 29 ][ 75 ],
   alphaCSR[ 29 ][ 76 ],
   alphaCSR[ 29 ][ 77 ],
   alphaCSR[ 29 ][ 78 ],
   alphaCSR[ 29 ][ 79 ],
   alphaCSR[ 29 ][ 80 ],
   alphaCSR[ 29 ][ 81 ],
   alphaCSR[ 29 ][ 82 ],
   alphaCSR[ 29 ][ 83 ],
   alphaCSR[ 29 ][ 84 ],
   alphaCSR[ 29 ][ 85 ],
   alphaCSR[ 29 ][ 86 ],
   alphaCSR[ 29 ][ 87 ],
   alphaCSR[ 29 ][ 88 ],
   alphaCSR[ 29 ][ 89 ],
   alphaCSR[ 29 ][ 90 ],
   alphaCSR[ 29 ][ 91 ],
   alphaCSR[ 29 ][ 92 ],
   alphaCSR[ 29 ][ 93 ],
   alphaCSR[ 29 ][ 94 ],
   alphaCSR[ 29 ][ 95 ],
   alphaCSR[ 29 ][ 96 ],
   alphaCSR[ 29 ][ 97 ],
   alphaCSR[ 29 ][ 98 ],
   alphaCSR[ 29 ][ 99 ],
   alphaCSR[ 29 ][ 100 ],
   alphaCSR[ 29 ][ 101 ],
   alphaCSR[ 29 ][ 102 ],
   alphaCSR[ 29 ][ 103 ],
   alphaCSR[ 29 ][ 104 ],
   alphaCSR[ 29 ][ 105 ],
   alphaCSR[ 29 ][ 106 ],
   alphaCSR[ 29 ][ 107 ],
   alphaCSR[ 29 ][ 108 ],
   alphaCSR[ 29 ][ 109 ],
   alphaCSR[ 29 ][ 110 ],
   alphaCSR[ 29 ][ 111 ],
   alphaCSR[ 29 ][ 112 ],
   alphaCSR[ 29 ][ 113 ],
   alphaCSR[ 29 ][ 114 ],
   alphaCSR[ 29 ][ 115 ],
   alphaCSR[ 29 ][ 116 ],
   alphaCSR[ 29 ][ 117 ],
   alphaCSR[ 29 ][ 118 ],
   alphaCSR[ 29 ][ 119 ],
   alphaCSR[ 29 ][ 120 ],
   alphaCSR[ 29 ][ 121 ],
   alphaCSR[ 29 ][ 122 ],
   alphaCSR[ 29 ][ 123 ],
   alphaCSR[ 29 ][ 124 ],
   alphaCSR[ 29 ][ 125 ],
   alphaCSR[ 29 ][ 126 ],
   alphaCSR[ 29 ][ 127 ],
   alphaCSR[ 29 ][ 128 ],
   alphaCSR[ 29 ][ 129 ],
   alphaCSR[ 29 ][ 130 ],
   alphaCSR[ 29 ][ 131 ],
   alphaCSR[ 29 ][ 132 ],
   alphaCSR[ 29 ][ 133 ],
   alphaCSR[ 29 ][ 134 ],
   alphaCSR[ 29 ][ 135 ],
   alphaCSR[ 29 ][ 136 ],
   alphaCSR[ 29 ][ 137 ],
   alphaCSR[ 29 ][ 138 ],
   alphaCSR[ 29 ][ 139 ],
   alphaCSR[ 29 ][ 140 ],
   alphaCSR[ 29 ][ 141 ],
   alphaCSR[ 29 ][ 142 ],
   alphaCSR[ 29 ][ 143 ],
   alphaCSR[ 29 ][ 144 ],
   alphaCSR[ 29 ][ 145 ],
   alphaCSR[ 29 ][ 146 ],
   alphaCSR[ 29 ][ 147 ],
   alphaCSR[ 29 ][ 148 ],
   alphaCSR[ 29 ][ 149 ],
   alphaCSR[ 29 ][ 150 ],
   alphaCSR[ 29 ][ 151 ],
   alphaCSR[ 29 ][ 152 ],
   alphaCSR[ 29 ][ 153 ],
   alphaCSR[ 29 ][ 154 ],
   alphaCSR[ 29 ][ 155 ],
   alphaCSR[ 29 ][ 156 ],
   alphaCSR[ 29 ][ 157 ],
   alphaCSR[ 29 ][ 158 ],
   alphaCSR[ 29 ][ 159 ],
   alphaCSR[ 29 ][ 160 ],
   alphaCSR[ 29 ][ 161 ],
   alphaCSR[ 29 ][ 162 ],
   alphaCSR[ 29 ][ 163 ],
   alphaCSR[ 29 ][ 164 ],
   alphaCSR[ 29 ][ 165 ],
   alphaCSR[ 29 ][ 166 ],
   alphaCSR[ 29 ][ 167 ],
   alphaCSR[ 29 ][ 168 ],
   alphaCSR[ 29 ][ 169 ],
   alphaCSR[ 29 ][ 170 ],
   alphaCSR[ 29 ][ 171 ],
   alphaCSR[ 29 ][ 172 ],
   alphaCSR[ 29 ][ 173 ],
   alphaCSR[ 29 ][ 174 ],
   alphaCSR[ 29 ][ 175 ],
   alphaCSR[ 29 ][ 176 ],
   alphaCSR[ 29 ][ 177 ],
   alphaCSR[ 29 ][ 178 ],
   alphaCSR[ 29 ][ 179 ],
   alphaCSR[ 29 ][ 180 ],
   alphaCSR[ 29 ][ 181 ],
   alphaCSR[ 29 ][ 182 ],
   alphaCSR[ 29 ][ 183 ],
   alphaCSR[ 29 ][ 184 ],
   alphaCSR[ 29 ][ 185 ],
   alphaCSR[ 29 ][ 186 ],
   alphaCSR[ 29 ][ 187 ],
   alphaCSR[ 29 ][ 188 ],
   alphaCSR[ 29 ][ 189 ],
   alphaCSR[ 29 ][ 190 ],
   alphaCSR[ 29 ][ 191 ],
   alphaCSR[ 29 ][ 192 ],
   alphaCSR[ 29 ][ 193 ],
   alphaCSR[ 29 ][ 194 ],
   alphaCSR[ 29 ][ 195 ],
   alphaCSR[ 29 ][ 196 ],
   alphaCSR[ 29 ][ 197 ],
   alphaCSR[ 29 ][ 198 ],
   alphaCSR[ 29 ][ 199 ],
   alphaCSR[ 29 ][ 200 ],
   alphaCSR[ 29 ][ 201 ],
   alphaCSR[ 29 ][ 202 ],
   alphaCSR[ 29 ][ 203 ],
   alphaCSR[ 29 ][ 204 ],
   alphaCSR[ 29 ][ 205 ],
   alphaCSR[ 29 ][ 206 ],
   alphaCSR[ 29 ][ 207 ],
   alphaCSR[ 29 ][ 208 ],
   alphaCSR[ 29 ][ 209 ],
   alphaCSR[ 29 ][ 210 ],
   alphaCSR[ 29 ][ 211 ],
   alphaCSR[ 29 ][ 212 ],
   alphaCSR[ 29 ][ 213 ],
   alphaCSR[ 29 ][ 214 ],
   alphaCSR[ 29 ][ 215 ],
   alphaCSR[ 29 ][ 216 ],
   alphaCSR[ 29 ][ 217 ],
   alphaCSR[ 29 ][ 218 ],
   alphaCSR[ 29 ][ 219 ],
   alphaCSR[ 29 ][ 220 ],
   alphaCSR[ 29 ][ 221 ],
   alphaCSR[ 29 ][ 222 ],
   alphaCSR[ 29 ][ 223 ],
   alphaCSR[ 29 ][ 224 ],
   alphaCSR[ 29 ][ 225 ],
   alphaCSR[ 29 ][ 226 ],
   alphaCSR[ 29 ][ 227 ],
   alphaCSR[ 29 ][ 228 ],
   alphaCSR[ 29 ][ 229 ],
   alphaCSR[ 29 ][ 230 ],
   alphaCSR[ 29 ][ 231 ],
   alphaCSR[ 29 ][ 232 ],
   alphaCSR[ 29 ][ 233 ],
   alphaCSR[ 29 ][ 234 ],
   alphaCSR[ 29 ][ 235 ],
   alphaCSR[ 29 ][ 236 ],
   alphaCSR[ 29 ][ 237 ],
   alphaCSR[ 29 ][ 238 ],
   alphaCSR[ 29 ][ 239 ],
   alphaCSR[ 29 ][ 240 ],
   alphaCSR[ 29 ][ 241 ],
   alphaCSR[ 29 ][ 242 ],
   alphaCSR[ 29 ][ 243 ],
   alphaCSR[ 29 ][ 244 ],
   alphaCSR[ 29 ][ 245 ],
   alphaCSR[ 29 ][ 246 ],
   alphaCSR[ 29 ][ 247 ],
   alphaCSR[ 29 ][ 248 ],
   alphaCSR[ 29 ][ 249 ],
   alphaCSR[ 29 ][ 250 ],
   alphaCSR[ 29 ][ 251 ],
   alphaCSR[ 29 ][ 252 ],
   alphaCSR[ 29 ][ 253 ],
   alphaCSR[ 29 ][ 254 ],
   alphaCSR[ 29 ][ 255 ],
   alphaCSR[ 29 ][ 256 ],
   alphaCSR[ 29 ][ 257 ],
   alphaCSR[ 29 ][ 258 ],
   alphaCSR[ 29 ][ 259 ],
   alphaCSR[ 29 ][ 260 ],
   alphaCSR[ 29 ][ 261 ],
   alphaCSR[ 29 ][ 262 ],
   alphaCSR[ 29 ][ 263 ],
   alphaCSR[ 29 ][ 264 ],
   alphaCSR[ 29 ][ 265 ],
   alphaCSR[ 29 ][ 266 ],
   alphaCSR[ 29 ][ 267 ],
   alphaCSR[ 29 ][ 268 ],
   alphaCSR[ 29 ][ 269 ],
   alphaCSR[ 29 ][ 270 ],
   alphaCSR[ 29 ][ 271 ],
   alphaCSR[ 29 ][ 272 ],
   alphaCSR[ 29 ][ 273 ],
   alphaCSR[ 29 ][ 274 ],
   alphaCSR[ 29 ][ 275 ],
   alphaCSR[ 29 ][ 276 ],
   alphaCSR[ 29 ][ 277 ],
   alphaCSR[ 29 ][ 278 ],
   alphaCSR[ 29 ][ 279 ],
   alphaCSR[ 29 ][ 280 ],
   alphaCSR[ 29 ][ 281 ],
   alphaCSR[ 29 ][ 282 ],
   alphaCSR[ 29 ][ 283 ],
   alphaCSR[ 29 ][ 284 ],
   alphaCSR[ 29 ][ 285 ],
   alphaCSR[ 29 ][ 286 ],
   alphaCSR[ 29 ][ 287 ],
   alphaCSR[ 29 ][ 288 ],
   alphaCSR[ 29 ][ 289 ],
   alphaCSR[ 29 ][ 290 ],
   alphaCSR[ 29 ][ 291 ],
   alphaCSR[ 29 ][ 292 ],
   alphaCSR[ 29 ][ 293 ],
   alphaCSR[ 29 ][ 294 ],
   alphaCSR[ 29 ][ 295 ],
   alphaCSR[ 29 ][ 296 ],
   alphaCSR[ 29 ][ 297 ],
   alphaCSR[ 29 ][ 298 ],
   alphaCSR[ 29 ][ 299 ],
   alphaCSR[ 29 ][ 300 ],
   alphaCSR[ 29 ][ 301 ],
   alphaCSR[ 29 ][ 302 ],
   alphaCSR[ 29 ][ 303 ],
   alphaCSR[ 29 ][ 304 ],
   alphaCSR[ 29 ][ 305 ],
   alphaCSR[ 29 ][ 306 ],
   alphaCSR[ 29 ][ 307 ],
   alphaCSR[ 29 ][ 308 ],
   alphaCSR[ 29 ][ 309 ],
   alphaCSR[ 29 ][ 310 ],
   alphaCSR[ 29 ][ 311 ],
   alphaCSR[ 29 ][ 312 ],
   alphaCSR[ 29 ][ 313 ],
   alphaCSR[ 29 ][ 314 ],
   alphaCSR[ 29 ][ 315 ],
   alphaCSR[ 29 ][ 316 ],
   alphaCSR[ 29 ][ 317 ],
   alphaCSR[ 29 ][ 318 ],
   alphaCSR[ 29 ][ 319 ],
   alphaCSR[ 29 ][ 320 ],
   alphaCSR[ 29 ][ 321 ],
   alphaCSR[ 29 ][ 322 ],
   alphaCSR[ 29 ][ 323 ],
   alphaCSR[ 29 ][ 324 ],
   alphaCSR[ 29 ][ 325 ],
   alphaCSR[ 29 ][ 326 ],
   alphaCSR[ 29 ][ 327 ],
   alphaCSR[ 29 ][ 328 ],
   alphaCSR[ 29 ][ 329 ],
   alphaCSR[ 29 ][ 330 ],
   alphaCSR[ 29 ][ 331 ],
   alphaCSR[ 29 ][ 332 ],
   alphaCSR[ 29 ][ 333 ],
   alphaCSR[ 29 ][ 334 ],
   alphaCSR[ 29 ][ 335 ],
   alphaCSR[ 29 ][ 336 ],
   alphaCSR[ 29 ][ 337 ],
   alphaCSR[ 29 ][ 338 ],
   alphaCSR[ 29 ][ 339 ],
   alphaCSR[ 29 ][ 340 ],
   alphaCSR[ 29 ][ 341 ],
   alphaCSR[ 29 ][ 342 ],
   alphaCSR[ 29 ][ 343 ],
   alphaCSR[ 29 ][ 344 ],
   alphaCSR[ 29 ][ 345 ],
   alphaCSR[ 29 ][ 346 ],
   alphaCSR[ 29 ][ 347 ],
   alphaCSR[ 29 ][ 348 ],
   alphaCSR[ 29 ][ 349 ],
   alphaCSR[ 29 ][ 350 ],
   alphaCSR[ 29 ][ 351 ],
   alphaCSR[ 29 ][ 352 ],
   alphaCSR[ 29 ][ 353 ],
   alphaCSR[ 29 ][ 354 ],
   alphaCSR[ 29 ][ 355 ],
   alphaCSR[ 29 ][ 356 ],
   alphaCSR[ 29 ][ 357 ],
   alphaCSR[ 29 ][ 358 ],
   alphaCSR[ 29 ][ 359 ],
   alphaCSR[ 29 ][ 360 ],
   alphaCSR[ 29 ][ 361 ],
   alphaCSR[ 29 ][ 362 ],
   alphaCSR[ 29 ][ 363 ],
   alphaCSR[ 29 ][ 364 ],
   alphaCSR[ 29 ][ 365 ],
   alphaCSR[ 29 ][ 366 ],
   alphaCSR[ 29 ][ 367 ],
   alphaCSR[ 29 ][ 368 ],
   alphaCSR[ 29 ][ 369 ],
   alphaCSR[ 29 ][ 370 ],
   alphaCSR[ 29 ][ 371 ],
   alphaCSR[ 29 ][ 372 ],
   alphaCSR[ 29 ][ 373 ],
   alphaCSR[ 29 ][ 374 ],
   alphaCSR[ 29 ][ 375 ],
   alphaCSR[ 29 ][ 376 ],
   alphaCSR[ 29 ][ 377 ],
   alphaCSR[ 29 ][ 378 ],
   alphaCSR[ 29 ][ 379 ],
   alphaCSR[ 29 ][ 380 ],
   alphaCSR[ 29 ][ 381 ],
   alphaCSR[ 29 ][ 382 ],
   alphaCSR[ 29 ][ 383 ],
   alphaCSR[ 30 ][ 0 ],
   alphaCSR[ 30 ][ 1 ],
   alphaCSR[ 30 ][ 2 ],
   alphaCSR[ 30 ][ 3 ],
   alphaCSR[ 30 ][ 4 ],
   alphaCSR[ 30 ][ 5 ],
   alphaCSR[ 30 ][ 6 ],
   alphaCSR[ 30 ][ 7 ],
   alphaCSR[ 30 ][ 8 ],
   alphaCSR[ 30 ][ 9 ],
   alphaCSR[ 30 ][ 10 ],
   alphaCSR[ 30 ][ 11 ],
   alphaCSR[ 30 ][ 12 ],
   alphaCSR[ 30 ][ 13 ],
   alphaCSR[ 30 ][ 14 ],
   alphaCSR[ 30 ][ 15 ],
   alphaCSR[ 30 ][ 16 ],
   alphaCSR[ 30 ][ 17 ],
   alphaCSR[ 30 ][ 18 ],
   alphaCSR[ 30 ][ 19 ],
   alphaCSR[ 30 ][ 20 ],
   alphaCSR[ 30 ][ 21 ],
   alphaCSR[ 30 ][ 22 ],
   alphaCSR[ 30 ][ 23 ],
   alphaCSR[ 30 ][ 24 ],
   alphaCSR[ 30 ][ 25 ],
   alphaCSR[ 30 ][ 26 ],
   alphaCSR[ 30 ][ 27 ],
   alphaCSR[ 30 ][ 28 ],
   alphaCSR[ 30 ][ 29 ],
   alphaCSR[ 30 ][ 30 ],
   alphaCSR[ 30 ][ 31 ],
   alphaCSR[ 30 ][ 32 ],
   alphaCSR[ 30 ][ 33 ],
   alphaCSR[ 30 ][ 34 ],
   alphaCSR[ 30 ][ 35 ],
   alphaCSR[ 30 ][ 36 ],
   alphaCSR[ 30 ][ 37 ],
   alphaCSR[ 30 ][ 38 ],
   alphaCSR[ 30 ][ 39 ],
   alphaCSR[ 30 ][ 40 ],
   alphaCSR[ 30 ][ 41 ],
   alphaCSR[ 30 ][ 42 ],
   alphaCSR[ 30 ][ 43 ],
   alphaCSR[ 30 ][ 44 ],
   alphaCSR[ 30 ][ 45 ],
   alphaCSR[ 30 ][ 46 ],
   alphaCSR[ 30 ][ 47 ],
   alphaCSR[ 30 ][ 48 ],
   alphaCSR[ 30 ][ 49 ],
   alphaCSR[ 30 ][ 50 ],
   alphaCSR[ 30 ][ 51 ],
   alphaCSR[ 30 ][ 52 ],
   alphaCSR[ 30 ][ 53 ],
   alphaCSR[ 30 ][ 54 ],
   alphaCSR[ 30 ][ 55 ],
   alphaCSR[ 30 ][ 56 ],
   alphaCSR[ 30 ][ 57 ],
   alphaCSR[ 30 ][ 58 ],
   alphaCSR[ 30 ][ 59 ],
   alphaCSR[ 30 ][ 60 ],
   alphaCSR[ 30 ][ 61 ],
   alphaCSR[ 30 ][ 62 ],
   alphaCSR[ 30 ][ 63 ],
   alphaCSR[ 30 ][ 64 ],
   alphaCSR[ 30 ][ 65 ],
   alphaCSR[ 30 ][ 66 ],
   alphaCSR[ 30 ][ 67 ],
   alphaCSR[ 30 ][ 68 ],
   alphaCSR[ 30 ][ 69 ],
   alphaCSR[ 30 ][ 70 ],
   alphaCSR[ 30 ][ 71 ],
   alphaCSR[ 30 ][ 72 ],
   alphaCSR[ 30 ][ 73 ],
   alphaCSR[ 30 ][ 74 ],
   alphaCSR[ 30 ][ 75 ],
   alphaCSR[ 30 ][ 76 ],
   alphaCSR[ 30 ][ 77 ],
   alphaCSR[ 30 ][ 78 ],
   alphaCSR[ 30 ][ 79 ],
   alphaCSR[ 30 ][ 80 ],
   alphaCSR[ 30 ][ 81 ],
   alphaCSR[ 30 ][ 82 ],
   alphaCSR[ 30 ][ 83 ],
   alphaCSR[ 30 ][ 84 ],
   alphaCSR[ 30 ][ 85 ],
   alphaCSR[ 30 ][ 86 ],
   alphaCSR[ 30 ][ 87 ],
   alphaCSR[ 30 ][ 88 ],
   alphaCSR[ 30 ][ 89 ],
   alphaCSR[ 30 ][ 90 ],
   alphaCSR[ 30 ][ 91 ],
   alphaCSR[ 30 ][ 92 ],
   alphaCSR[ 30 ][ 93 ],
   alphaCSR[ 30 ][ 94 ],
   alphaCSR[ 30 ][ 95 ],
   alphaCSR[ 30 ][ 96 ],
   alphaCSR[ 30 ][ 97 ],
   alphaCSR[ 30 ][ 98 ],
   alphaCSR[ 30 ][ 99 ],
   alphaCSR[ 30 ][ 100 ],
   alphaCSR[ 30 ][ 101 ],
   alphaCSR[ 30 ][ 102 ],
   alphaCSR[ 30 ][ 103 ],
   alphaCSR[ 30 ][ 104 ],
   alphaCSR[ 30 ][ 105 ],
   alphaCSR[ 30 ][ 106 ],
   alphaCSR[ 30 ][ 107 ],
   alphaCSR[ 30 ][ 108 ],
   alphaCSR[ 30 ][ 109 ],
   alphaCSR[ 30 ][ 110 ],
   alphaCSR[ 30 ][ 111 ],
   alphaCSR[ 30 ][ 112 ],
   alphaCSR[ 30 ][ 113 ],
   alphaCSR[ 30 ][ 114 ],
   alphaCSR[ 30 ][ 115 ],
   alphaCSR[ 30 ][ 116 ],
   alphaCSR[ 30 ][ 117 ],
   alphaCSR[ 30 ][ 118 ],
   alphaCSR[ 30 ][ 119 ],
   alphaCSR[ 30 ][ 120 ],
   alphaCSR[ 30 ][ 121 ],
   alphaCSR[ 30 ][ 122 ],
   alphaCSR[ 30 ][ 123 ],
   alphaCSR[ 30 ][ 124 ],
   alphaCSR[ 30 ][ 125 ],
   alphaCSR[ 30 ][ 126 ],
   alphaCSR[ 30 ][ 127 ],
   alphaCSR[ 30 ][ 128 ],
   alphaCSR[ 30 ][ 129 ],
   alphaCSR[ 30 ][ 130 ],
   alphaCSR[ 30 ][ 131 ],
   alphaCSR[ 30 ][ 132 ],
   alphaCSR[ 30 ][ 133 ],
   alphaCSR[ 30 ][ 134 ],
   alphaCSR[ 30 ][ 135 ],
   alphaCSR[ 30 ][ 136 ],
   alphaCSR[ 30 ][ 137 ],
   alphaCSR[ 30 ][ 138 ],
   alphaCSR[ 30 ][ 139 ],
   alphaCSR[ 30 ][ 140 ],
   alphaCSR[ 30 ][ 141 ],
   alphaCSR[ 30 ][ 142 ],
   alphaCSR[ 30 ][ 143 ],
   alphaCSR[ 30 ][ 144 ],
   alphaCSR[ 30 ][ 145 ],
   alphaCSR[ 30 ][ 146 ],
   alphaCSR[ 30 ][ 147 ],
   alphaCSR[ 30 ][ 148 ],
   alphaCSR[ 30 ][ 149 ],
   alphaCSR[ 30 ][ 150 ],
   alphaCSR[ 30 ][ 151 ],
   alphaCSR[ 30 ][ 152 ],
   alphaCSR[ 30 ][ 153 ],
   alphaCSR[ 30 ][ 154 ],
   alphaCSR[ 30 ][ 155 ],
   alphaCSR[ 30 ][ 156 ],
   alphaCSR[ 30 ][ 157 ],
   alphaCSR[ 30 ][ 158 ],
   alphaCSR[ 30 ][ 159 ],
   alphaCSR[ 30 ][ 160 ],
   alphaCSR[ 30 ][ 161 ],
   alphaCSR[ 30 ][ 162 ],
   alphaCSR[ 30 ][ 163 ],
   alphaCSR[ 30 ][ 164 ],
   alphaCSR[ 30 ][ 165 ],
   alphaCSR[ 30 ][ 166 ],
   alphaCSR[ 30 ][ 167 ],
   alphaCSR[ 30 ][ 168 ],
   alphaCSR[ 30 ][ 169 ],
   alphaCSR[ 30 ][ 170 ],
   alphaCSR[ 30 ][ 171 ],
   alphaCSR[ 30 ][ 172 ],
   alphaCSR[ 30 ][ 173 ],
   alphaCSR[ 30 ][ 174 ],
   alphaCSR[ 30 ][ 175 ],
   alphaCSR[ 30 ][ 176 ],
   alphaCSR[ 30 ][ 177 ],
   alphaCSR[ 30 ][ 178 ],
   alphaCSR[ 30 ][ 179 ],
   alphaCSR[ 30 ][ 180 ],
   alphaCSR[ 30 ][ 181 ],
   alphaCSR[ 30 ][ 182 ],
   alphaCSR[ 30 ][ 183 ],
   alphaCSR[ 30 ][ 184 ],
   alphaCSR[ 30 ][ 185 ],
   alphaCSR[ 30 ][ 186 ],
   alphaCSR[ 30 ][ 187 ],
   alphaCSR[ 30 ][ 188 ],
   alphaCSR[ 30 ][ 189 ],
   alphaCSR[ 30 ][ 190 ],
   alphaCSR[ 30 ][ 191 ],
   alphaCSR[ 30 ][ 192 ],
   alphaCSR[ 30 ][ 193 ],
   alphaCSR[ 30 ][ 194 ],
   alphaCSR[ 30 ][ 195 ],
   alphaCSR[ 30 ][ 196 ],
   alphaCSR[ 30 ][ 197 ],
   alphaCSR[ 30 ][ 198 ],
   alphaCSR[ 30 ][ 199 ],
   alphaCSR[ 30 ][ 200 ],
   alphaCSR[ 30 ][ 201 ],
   alphaCSR[ 30 ][ 202 ],
   alphaCSR[ 30 ][ 203 ],
   alphaCSR[ 30 ][ 204 ],
   alphaCSR[ 30 ][ 205 ],
   alphaCSR[ 30 ][ 206 ],
   alphaCSR[ 30 ][ 207 ],
   alphaCSR[ 30 ][ 208 ],
   alphaCSR[ 30 ][ 209 ],
   alphaCSR[ 30 ][ 210 ],
   alphaCSR[ 30 ][ 211 ],
   alphaCSR[ 30 ][ 212 ],
   alphaCSR[ 30 ][ 213 ],
   alphaCSR[ 30 ][ 214 ],
   alphaCSR[ 30 ][ 215 ],
   alphaCSR[ 30 ][ 216 ],
   alphaCSR[ 30 ][ 217 ],
   alphaCSR[ 30 ][ 218 ],
   alphaCSR[ 30 ][ 219 ],
   alphaCSR[ 30 ][ 220 ],
   alphaCSR[ 30 ][ 221 ],
   alphaCSR[ 30 ][ 222 ],
   alphaCSR[ 30 ][ 223 ],
   alphaCSR[ 30 ][ 224 ],
   alphaCSR[ 30 ][ 225 ],
   alphaCSR[ 30 ][ 226 ],
   alphaCSR[ 30 ][ 227 ],
   alphaCSR[ 30 ][ 228 ],
   alphaCSR[ 30 ][ 229 ],
   alphaCSR[ 30 ][ 230 ],
   alphaCSR[ 30 ][ 231 ],
   alphaCSR[ 30 ][ 232 ],
   alphaCSR[ 30 ][ 233 ],
   alphaCSR[ 30 ][ 234 ],
   alphaCSR[ 30 ][ 235 ],
   alphaCSR[ 30 ][ 236 ],
   alphaCSR[ 30 ][ 237 ],
   alphaCSR[ 30 ][ 238 ],
   alphaCSR[ 30 ][ 239 ],
   alphaCSR[ 30 ][ 240 ],
   alphaCSR[ 30 ][ 241 ],
   alphaCSR[ 30 ][ 242 ],
   alphaCSR[ 30 ][ 243 ],
   alphaCSR[ 30 ][ 244 ],
   alphaCSR[ 30 ][ 245 ],
   alphaCSR[ 30 ][ 246 ],
   alphaCSR[ 30 ][ 247 ],
   alphaCSR[ 30 ][ 248 ],
   alphaCSR[ 30 ][ 249 ],
   alphaCSR[ 30 ][ 250 ],
   alphaCSR[ 30 ][ 251 ],
   alphaCSR[ 30 ][ 252 ],
   alphaCSR[ 30 ][ 253 ],
   alphaCSR[ 30 ][ 254 ],
   alphaCSR[ 30 ][ 255 ],
   alphaCSR[ 30 ][ 256 ],
   alphaCSR[ 30 ][ 257 ],
   alphaCSR[ 30 ][ 258 ],
   alphaCSR[ 30 ][ 259 ],
   alphaCSR[ 30 ][ 260 ],
   alphaCSR[ 30 ][ 261 ],
   alphaCSR[ 30 ][ 262 ],
   alphaCSR[ 30 ][ 263 ],
   alphaCSR[ 30 ][ 264 ],
   alphaCSR[ 30 ][ 265 ],
   alphaCSR[ 30 ][ 266 ],
   alphaCSR[ 30 ][ 267 ],
   alphaCSR[ 30 ][ 268 ],
   alphaCSR[ 30 ][ 269 ],
   alphaCSR[ 30 ][ 270 ],
   alphaCSR[ 30 ][ 271 ],
   alphaCSR[ 30 ][ 272 ],
   alphaCSR[ 30 ][ 273 ],
   alphaCSR[ 30 ][ 274 ],
   alphaCSR[ 30 ][ 275 ],
   alphaCSR[ 30 ][ 276 ],
   alphaCSR[ 30 ][ 277 ],
   alphaCSR[ 30 ][ 278 ],
   alphaCSR[ 30 ][ 279 ],
   alphaCSR[ 30 ][ 280 ],
   alphaCSR[ 30 ][ 281 ],
   alphaCSR[ 30 ][ 282 ],
   alphaCSR[ 30 ][ 283 ],
   alphaCSR[ 30 ][ 284 ],
   alphaCSR[ 30 ][ 285 ],
   alphaCSR[ 30 ][ 286 ],
   alphaCSR[ 30 ][ 287 ],
   alphaCSR[ 30 ][ 288 ],
   alphaCSR[ 30 ][ 289 ],
   alphaCSR[ 30 ][ 290 ],
   alphaCSR[ 30 ][ 291 ],
   alphaCSR[ 30 ][ 292 ],
   alphaCSR[ 30 ][ 293 ],
   alphaCSR[ 30 ][ 294 ],
   alphaCSR[ 30 ][ 295 ],
   alphaCSR[ 30 ][ 296 ],
   alphaCSR[ 30 ][ 297 ],
   alphaCSR[ 30 ][ 298 ],
   alphaCSR[ 30 ][ 299 ],
   alphaCSR[ 30 ][ 300 ],
   alphaCSR[ 30 ][ 301 ],
   alphaCSR[ 30 ][ 302 ],
   alphaCSR[ 30 ][ 303 ],
   alphaCSR[ 30 ][ 304 ],
   alphaCSR[ 30 ][ 305 ],
   alphaCSR[ 30 ][ 306 ],
   alphaCSR[ 30 ][ 307 ],
   alphaCSR[ 30 ][ 308 ],
   alphaCSR[ 30 ][ 309 ],
   alphaCSR[ 30 ][ 310 ],
   alphaCSR[ 30 ][ 311 ],
   alphaCSR[ 30 ][ 312 ],
   alphaCSR[ 30 ][ 313 ],
   alphaCSR[ 30 ][ 314 ],
   alphaCSR[ 30 ][ 315 ],
   alphaCSR[ 30 ][ 316 ],
   alphaCSR[ 30 ][ 317 ],
   alphaCSR[ 30 ][ 318 ],
   alphaCSR[ 30 ][ 319 ],
   alphaCSR[ 30 ][ 320 ],
   alphaCSR[ 30 ][ 321 ],
   alphaCSR[ 30 ][ 322 ],
   alphaCSR[ 30 ][ 323 ],
   alphaCSR[ 30 ][ 324 ],
   alphaCSR[ 30 ][ 325 ],
   alphaCSR[ 30 ][ 326 ],
   alphaCSR[ 30 ][ 327 ],
   alphaCSR[ 30 ][ 328 ],
   alphaCSR[ 30 ][ 329 ],
   alphaCSR[ 30 ][ 330 ],
   alphaCSR[ 30 ][ 331 ],
   alphaCSR[ 30 ][ 332 ],
   alphaCSR[ 30 ][ 333 ],
   alphaCSR[ 30 ][ 334 ],
   alphaCSR[ 30 ][ 335 ],
   alphaCSR[ 30 ][ 336 ],
   alphaCSR[ 30 ][ 337 ],
   alphaCSR[ 30 ][ 338 ],
   alphaCSR[ 30 ][ 339 ],
   alphaCSR[ 30 ][ 340 ],
   alphaCSR[ 30 ][ 341 ],
   alphaCSR[ 30 ][ 342 ],
   alphaCSR[ 30 ][ 343 ],
   alphaCSR[ 30 ][ 344 ],
   alphaCSR[ 30 ][ 345 ],
   alphaCSR[ 30 ][ 346 ],
   alphaCSR[ 30 ][ 347 ],
   alphaCSR[ 30 ][ 348 ],
   alphaCSR[ 30 ][ 349 ],
   alphaCSR[ 30 ][ 350 ],
   alphaCSR[ 30 ][ 351 ],
   alphaCSR[ 30 ][ 352 ],
   alphaCSR[ 30 ][ 353 ],
   alphaCSR[ 30 ][ 354 ],
   alphaCSR[ 30 ][ 355 ],
   alphaCSR[ 30 ][ 356 ],
   alphaCSR[ 30 ][ 357 ],
   alphaCSR[ 30 ][ 358 ],
   alphaCSR[ 30 ][ 359 ],
   alphaCSR[ 30 ][ 360 ],
   alphaCSR[ 30 ][ 361 ],
   alphaCSR[ 30 ][ 362 ],
   alphaCSR[ 30 ][ 363 ],
   alphaCSR[ 30 ][ 364 ],
   alphaCSR[ 30 ][ 365 ],
   alphaCSR[ 30 ][ 366 ],
   alphaCSR[ 30 ][ 367 ],
   alphaCSR[ 30 ][ 368 ],
   alphaCSR[ 30 ][ 369 ],
   alphaCSR[ 30 ][ 370 ],
   alphaCSR[ 30 ][ 371 ],
   alphaCSR[ 30 ][ 372 ],
   alphaCSR[ 30 ][ 373 ],
   alphaCSR[ 30 ][ 374 ],
   alphaCSR[ 30 ][ 375 ],
   alphaCSR[ 30 ][ 376 ],
   alphaCSR[ 30 ][ 377 ],
   alphaCSR[ 30 ][ 378 ],
   alphaCSR[ 30 ][ 379 ],
   alphaCSR[ 30 ][ 380 ],
   alphaCSR[ 30 ][ 381 ],
   alphaCSR[ 30 ][ 382 ],
   alphaCSR[ 30 ][ 383 ],
   alphaCSR[ 31 ][ 0 ],
   alphaCSR[ 31 ][ 1 ],
   alphaCSR[ 31 ][ 2 ],
   alphaCSR[ 31 ][ 3 ],
   alphaCSR[ 31 ][ 4 ],
   alphaCSR[ 31 ][ 5 ],
   alphaCSR[ 31 ][ 6 ],
   alphaCSR[ 31 ][ 7 ],
   alphaCSR[ 31 ][ 8 ],
   alphaCSR[ 31 ][ 9 ],
   alphaCSR[ 31 ][ 10 ],
   alphaCSR[ 31 ][ 11 ],
   alphaCSR[ 31 ][ 12 ],
   alphaCSR[ 31 ][ 13 ],
   alphaCSR[ 31 ][ 14 ],
   alphaCSR[ 31 ][ 15 ],
   alphaCSR[ 31 ][ 16 ],
   alphaCSR[ 31 ][ 17 ],
   alphaCSR[ 31 ][ 18 ],
   alphaCSR[ 31 ][ 19 ],
   alphaCSR[ 31 ][ 20 ],
   alphaCSR[ 31 ][ 21 ],
   alphaCSR[ 31 ][ 22 ],
   alphaCSR[ 31 ][ 23 ],
   alphaCSR[ 31 ][ 24 ],
   alphaCSR[ 31 ][ 25 ],
   alphaCSR[ 31 ][ 26 ],
   alphaCSR[ 31 ][ 27 ],
   alphaCSR[ 31 ][ 28 ],
   alphaCSR[ 31 ][ 29 ],
   alphaCSR[ 31 ][ 30 ],
   alphaCSR[ 31 ][ 31 ],
   alphaCSR[ 31 ][ 32 ],
   alphaCSR[ 31 ][ 33 ],
   alphaCSR[ 31 ][ 34 ],
   alphaCSR[ 31 ][ 35 ],
   alphaCSR[ 31 ][ 36 ],
   alphaCSR[ 31 ][ 37 ],
   alphaCSR[ 31 ][ 38 ],
   alphaCSR[ 31 ][ 39 ],
   alphaCSR[ 31 ][ 40 ],
   alphaCSR[ 31 ][ 41 ],
   alphaCSR[ 31 ][ 42 ],
   alphaCSR[ 31 ][ 43 ],
   alphaCSR[ 31 ][ 44 ],
   alphaCSR[ 31 ][ 45 ],
   alphaCSR[ 31 ][ 46 ],
   alphaCSR[ 31 ][ 47 ],
   alphaCSR[ 31 ][ 48 ],
   alphaCSR[ 31 ][ 49 ],
   alphaCSR[ 31 ][ 50 ],
   alphaCSR[ 31 ][ 51 ],
   alphaCSR[ 31 ][ 52 ],
   alphaCSR[ 31 ][ 53 ],
   alphaCSR[ 31 ][ 54 ],
   alphaCSR[ 31 ][ 55 ],
   alphaCSR[ 31 ][ 56 ],
   alphaCSR[ 31 ][ 57 ],
   alphaCSR[ 31 ][ 58 ],
   alphaCSR[ 31 ][ 59 ],
   alphaCSR[ 31 ][ 60 ],
   alphaCSR[ 31 ][ 61 ],
   alphaCSR[ 31 ][ 62 ],
   alphaCSR[ 31 ][ 63 ],
   alphaCSR[ 31 ][ 64 ],
   alphaCSR[ 31 ][ 65 ],
   alphaCSR[ 31 ][ 66 ],
   alphaCSR[ 31 ][ 67 ],
   alphaCSR[ 31 ][ 68 ],
   alphaCSR[ 31 ][ 69 ],
   alphaCSR[ 31 ][ 70 ],
   alphaCSR[ 31 ][ 71 ],
   alphaCSR[ 31 ][ 72 ],
   alphaCSR[ 31 ][ 73 ],
   alphaCSR[ 31 ][ 74 ],
   alphaCSR[ 31 ][ 75 ],
   alphaCSR[ 31 ][ 76 ],
   alphaCSR[ 31 ][ 77 ],
   alphaCSR[ 31 ][ 78 ],
   alphaCSR[ 31 ][ 79 ],
   alphaCSR[ 31 ][ 80 ],
   alphaCSR[ 31 ][ 81 ],
   alphaCSR[ 31 ][ 82 ],
   alphaCSR[ 31 ][ 83 ],
   alphaCSR[ 31 ][ 84 ],
   alphaCSR[ 31 ][ 85 ],
   alphaCSR[ 31 ][ 86 ],
   alphaCSR[ 31 ][ 87 ],
   alphaCSR[ 31 ][ 88 ],
   alphaCSR[ 31 ][ 89 ],
   alphaCSR[ 31 ][ 90 ],
   alphaCSR[ 31 ][ 91 ],
   alphaCSR[ 31 ][ 92 ],
   alphaCSR[ 31 ][ 93 ],
   alphaCSR[ 31 ][ 94 ],
   alphaCSR[ 31 ][ 95 ],
   alphaCSR[ 31 ][ 96 ],
   alphaCSR[ 31 ][ 97 ],
   alphaCSR[ 31 ][ 98 ],
   alphaCSR[ 31 ][ 99 ],
   alphaCSR[ 31 ][ 100 ],
   alphaCSR[ 31 ][ 101 ],
   alphaCSR[ 31 ][ 102 ],
   alphaCSR[ 31 ][ 103 ],
   alphaCSR[ 31 ][ 104 ],
   alphaCSR[ 31 ][ 105 ],
   alphaCSR[ 31 ][ 106 ],
   alphaCSR[ 31 ][ 107 ],
   alphaCSR[ 31 ][ 108 ],
   alphaCSR[ 31 ][ 109 ],
   alphaCSR[ 31 ][ 110 ],
   alphaCSR[ 31 ][ 111 ],
   alphaCSR[ 31 ][ 112 ],
   alphaCSR[ 31 ][ 113 ],
   alphaCSR[ 31 ][ 114 ],
   alphaCSR[ 31 ][ 115 ],
   alphaCSR[ 31 ][ 116 ],
   alphaCSR[ 31 ][ 117 ],
   alphaCSR[ 31 ][ 118 ],
   alphaCSR[ 31 ][ 119 ],
   alphaCSR[ 31 ][ 120 ],
   alphaCSR[ 31 ][ 121 ],
   alphaCSR[ 31 ][ 122 ],
   alphaCSR[ 31 ][ 123 ],
   alphaCSR[ 31 ][ 124 ],
   alphaCSR[ 31 ][ 125 ],
   alphaCSR[ 31 ][ 126 ],
   alphaCSR[ 31 ][ 127 ],
   alphaCSR[ 31 ][ 128 ],
   alphaCSR[ 31 ][ 129 ],
   alphaCSR[ 31 ][ 130 ],
   alphaCSR[ 31 ][ 131 ],
   alphaCSR[ 31 ][ 132 ],
   alphaCSR[ 31 ][ 133 ],
   alphaCSR[ 31 ][ 134 ],
   alphaCSR[ 31 ][ 135 ],
   alphaCSR[ 31 ][ 136 ],
   alphaCSR[ 31 ][ 137 ],
   alphaCSR[ 31 ][ 138 ],
   alphaCSR[ 31 ][ 139 ],
   alphaCSR[ 31 ][ 140 ],
   alphaCSR[ 31 ][ 141 ],
   alphaCSR[ 31 ][ 142 ],
   alphaCSR[ 31 ][ 143 ],
   alphaCSR[ 31 ][ 144 ],
   alphaCSR[ 31 ][ 145 ],
   alphaCSR[ 31 ][ 146 ],
   alphaCSR[ 31 ][ 147 ],
   alphaCSR[ 31 ][ 148 ],
   alphaCSR[ 31 ][ 149 ],
   alphaCSR[ 31 ][ 150 ],
   alphaCSR[ 31 ][ 151 ],
   alphaCSR[ 31 ][ 152 ],
   alphaCSR[ 31 ][ 153 ],
   alphaCSR[ 31 ][ 154 ],
   alphaCSR[ 31 ][ 155 ],
   alphaCSR[ 31 ][ 156 ],
   alphaCSR[ 31 ][ 157 ],
   alphaCSR[ 31 ][ 158 ],
   alphaCSR[ 31 ][ 159 ],
   alphaCSR[ 31 ][ 160 ],
   alphaCSR[ 31 ][ 161 ],
   alphaCSR[ 31 ][ 162 ],
   alphaCSR[ 31 ][ 163 ],
   alphaCSR[ 31 ][ 164 ],
   alphaCSR[ 31 ][ 165 ],
   alphaCSR[ 31 ][ 166 ],
   alphaCSR[ 31 ][ 167 ],
   alphaCSR[ 31 ][ 168 ],
   alphaCSR[ 31 ][ 169 ],
   alphaCSR[ 31 ][ 170 ],
   alphaCSR[ 31 ][ 171 ],
   alphaCSR[ 31 ][ 172 ],
   alphaCSR[ 31 ][ 173 ],
   alphaCSR[ 31 ][ 174 ],
   alphaCSR[ 31 ][ 175 ],
   alphaCSR[ 31 ][ 176 ],
   alphaCSR[ 31 ][ 177 ],
   alphaCSR[ 31 ][ 178 ],
   alphaCSR[ 31 ][ 179 ],
   alphaCSR[ 31 ][ 180 ],
   alphaCSR[ 31 ][ 181 ],
   alphaCSR[ 31 ][ 182 ],
   alphaCSR[ 31 ][ 183 ],
   alphaCSR[ 31 ][ 184 ],
   alphaCSR[ 31 ][ 185 ],
   alphaCSR[ 31 ][ 186 ],
   alphaCSR[ 31 ][ 187 ],
   alphaCSR[ 31 ][ 188 ],
   alphaCSR[ 31 ][ 189 ],
   alphaCSR[ 31 ][ 190 ],
   alphaCSR[ 31 ][ 191 ],
   alphaCSR[ 31 ][ 192 ],
   alphaCSR[ 31 ][ 193 ],
   alphaCSR[ 31 ][ 194 ],
   alphaCSR[ 31 ][ 195 ],
   alphaCSR[ 31 ][ 196 ],
   alphaCSR[ 31 ][ 197 ],
   alphaCSR[ 31 ][ 198 ],
   alphaCSR[ 31 ][ 199 ],
   alphaCSR[ 31 ][ 200 ],
   alphaCSR[ 31 ][ 201 ],
   alphaCSR[ 31 ][ 202 ],
   alphaCSR[ 31 ][ 203 ],
   alphaCSR[ 31 ][ 204 ],
   alphaCSR[ 31 ][ 205 ],
   alphaCSR[ 31 ][ 206 ],
   alphaCSR[ 31 ][ 207 ],
   alphaCSR[ 31 ][ 208 ],
   alphaCSR[ 31 ][ 209 ],
   alphaCSR[ 31 ][ 210 ],
   alphaCSR[ 31 ][ 211 ],
   alphaCSR[ 31 ][ 212 ],
   alphaCSR[ 31 ][ 213 ],
   alphaCSR[ 31 ][ 214 ],
   alphaCSR[ 31 ][ 215 ],
   alphaCSR[ 31 ][ 216 ],
   alphaCSR[ 31 ][ 217 ],
   alphaCSR[ 31 ][ 218 ],
   alphaCSR[ 31 ][ 219 ],
   alphaCSR[ 31 ][ 220 ],
   alphaCSR[ 31 ][ 221 ],
   alphaCSR[ 31 ][ 222 ],
   alphaCSR[ 31 ][ 223 ],
   alphaCSR[ 31 ][ 224 ],
   alphaCSR[ 31 ][ 225 ],
   alphaCSR[ 31 ][ 226 ],
   alphaCSR[ 31 ][ 227 ],
   alphaCSR[ 31 ][ 228 ],
   alphaCSR[ 31 ][ 229 ],
   alphaCSR[ 31 ][ 230 ],
   alphaCSR[ 31 ][ 231 ],
   alphaCSR[ 31 ][ 232 ],
   alphaCSR[ 31 ][ 233 ],
   alphaCSR[ 31 ][ 234 ],
   alphaCSR[ 31 ][ 235 ],
   alphaCSR[ 31 ][ 236 ],
   alphaCSR[ 31 ][ 237 ],
   alphaCSR[ 31 ][ 238 ],
   alphaCSR[ 31 ][ 239 ],
   alphaCSR[ 31 ][ 240 ],
   alphaCSR[ 31 ][ 241 ],
   alphaCSR[ 31 ][ 242 ],
   alphaCSR[ 31 ][ 243 ],
   alphaCSR[ 31 ][ 244 ],
   alphaCSR[ 31 ][ 245 ],
   alphaCSR[ 31 ][ 246 ],
   alphaCSR[ 31 ][ 247 ],
   alphaCSR[ 31 ][ 248 ],
   alphaCSR[ 31 ][ 249 ],
   alphaCSR[ 31 ][ 250 ],
   alphaCSR[ 31 ][ 251 ],
   alphaCSR[ 31 ][ 252 ],
   alphaCSR[ 31 ][ 253 ],
   alphaCSR[ 31 ][ 254 ],
   alphaCSR[ 31 ][ 255 ],
   alphaCSR[ 31 ][ 256 ],
   alphaCSR[ 31 ][ 257 ],
   alphaCSR[ 31 ][ 258 ],
   alphaCSR[ 31 ][ 259 ],
   alphaCSR[ 31 ][ 260 ],
   alphaCSR[ 31 ][ 261 ],
   alphaCSR[ 31 ][ 262 ],
   alphaCSR[ 31 ][ 263 ],
   alphaCSR[ 31 ][ 264 ],
   alphaCSR[ 31 ][ 265 ],
   alphaCSR[ 31 ][ 266 ],
   alphaCSR[ 31 ][ 267 ],
   alphaCSR[ 31 ][ 268 ],
   alphaCSR[ 31 ][ 269 ],
   alphaCSR[ 31 ][ 270 ],
   alphaCSR[ 31 ][ 271 ],
   alphaCSR[ 31 ][ 272 ],
   alphaCSR[ 31 ][ 273 ],
   alphaCSR[ 31 ][ 274 ],
   alphaCSR[ 31 ][ 275 ],
   alphaCSR[ 31 ][ 276 ],
   alphaCSR[ 31 ][ 277 ],
   alphaCSR[ 31 ][ 278 ],
   alphaCSR[ 31 ][ 279 ],
   alphaCSR[ 31 ][ 280 ],
   alphaCSR[ 31 ][ 281 ],
   alphaCSR[ 31 ][ 282 ],
   alphaCSR[ 31 ][ 283 ],
   alphaCSR[ 31 ][ 284 ],
   alphaCSR[ 31 ][ 285 ],
   alphaCSR[ 31 ][ 286 ],
   alphaCSR[ 31 ][ 287 ],
   alphaCSR[ 31 ][ 288 ],
   alphaCSR[ 31 ][ 289 ],
   alphaCSR[ 31 ][ 290 ],
   alphaCSR[ 31 ][ 291 ],
   alphaCSR[ 31 ][ 292 ],
   alphaCSR[ 31 ][ 293 ],
   alphaCSR[ 31 ][ 294 ],
   alphaCSR[ 31 ][ 295 ],
   alphaCSR[ 31 ][ 296 ],
   alphaCSR[ 31 ][ 297 ],
   alphaCSR[ 31 ][ 298 ],
   alphaCSR[ 31 ][ 299 ],
   alphaCSR[ 31 ][ 300 ],
   alphaCSR[ 31 ][ 301 ],
   alphaCSR[ 31 ][ 302 ],
   alphaCSR[ 31 ][ 303 ],
   alphaCSR[ 31 ][ 304 ],
   alphaCSR[ 31 ][ 305 ],
   alphaCSR[ 31 ][ 306 ],
   alphaCSR[ 31 ][ 307 ],
   alphaCSR[ 31 ][ 308 ],
   alphaCSR[ 31 ][ 309 ],
   alphaCSR[ 31 ][ 310 ],
   alphaCSR[ 31 ][ 311 ],
   alphaCSR[ 31 ][ 312 ],
   alphaCSR[ 31 ][ 313 ],
   alphaCSR[ 31 ][ 314 ],
   alphaCSR[ 31 ][ 315 ],
   alphaCSR[ 31 ][ 316 ],
   alphaCSR[ 31 ][ 317 ],
   alphaCSR[ 31 ][ 318 ],
   alphaCSR[ 31 ][ 319 ],
   alphaCSR[ 31 ][ 320 ],
   alphaCSR[ 31 ][ 321 ],
   alphaCSR[ 31 ][ 322 ],
   alphaCSR[ 31 ][ 323 ],
   alphaCSR[ 31 ][ 324 ],
   alphaCSR[ 31 ][ 325 ],
   alphaCSR[ 31 ][ 326 ],
   alphaCSR[ 31 ][ 327 ],
   alphaCSR[ 31 ][ 328 ],
   alphaCSR[ 31 ][ 329 ],
   alphaCSR[ 31 ][ 330 ],
   alphaCSR[ 31 ][ 331 ],
   alphaCSR[ 31 ][ 332 ],
   alphaCSR[ 31 ][ 333 ],
   alphaCSR[ 31 ][ 334 ],
   alphaCSR[ 31 ][ 335 ],
   alphaCSR[ 31 ][ 336 ],
   alphaCSR[ 31 ][ 337 ],
   alphaCSR[ 31 ][ 338 ],
   alphaCSR[ 31 ][ 339 ],
   alphaCSR[ 31 ][ 340 ],
   alphaCSR[ 31 ][ 341 ],
   alphaCSR[ 31 ][ 342 ],
   alphaCSR[ 31 ][ 343 ],
   alphaCSR[ 31 ][ 344 ],
   alphaCSR[ 31 ][ 345 ],
   alphaCSR[ 31 ][ 346 ],
   alphaCSR[ 31 ][ 347 ],
   alphaCSR[ 31 ][ 348 ],
   alphaCSR[ 31 ][ 349 ],
   alphaCSR[ 31 ][ 350 ],
   alphaCSR[ 31 ][ 351 ],
   alphaCSR[ 31 ][ 352 ],
   alphaCSR[ 31 ][ 353 ],
   alphaCSR[ 31 ][ 354 ],
   alphaCSR[ 31 ][ 355 ],
   alphaCSR[ 31 ][ 356 ],
   alphaCSR[ 31 ][ 357 ],
   alphaCSR[ 31 ][ 358 ],
   alphaCSR[ 31 ][ 359 ],
   alphaCSR[ 31 ][ 360 ],
   alphaCSR[ 31 ][ 361 ],
   alphaCSR[ 31 ][ 362 ],
   alphaCSR[ 31 ][ 363 ],
   alphaCSR[ 31 ][ 364 ],
   alphaCSR[ 31 ][ 365 ],
   alphaCSR[ 31 ][ 366 ],
   alphaCSR[ 31 ][ 367 ],
   alphaCSR[ 31 ][ 368 ],
   alphaCSR[ 31 ][ 369 ],
   alphaCSR[ 31 ][ 370 ],
   alphaCSR[ 31 ][ 371 ],
   alphaCSR[ 31 ][ 372 ],
   alphaCSR[ 31 ][ 373 ],
   alphaCSR[ 31 ][ 374 ],
   alphaCSR[ 31 ][ 375 ],
   alphaCSR[ 31 ][ 376 ],
   alphaCSR[ 31 ][ 377 ],
   alphaCSR[ 31 ][ 378 ],
   alphaCSR[ 31 ][ 379 ],
   alphaCSR[ 31 ][ 380 ],
   alphaCSR[ 31 ][ 381 ],
   alphaCSR[ 31 ][ 382 ],
   alphaCSR[ 31 ][ 383 ],
   alphaCSR[ 32 ][ 0 ],
   alphaCSR[ 32 ][ 1 ],
   alphaCSR[ 32 ][ 2 ],
   alphaCSR[ 32 ][ 3 ],
   alphaCSR[ 32 ][ 4 ],
   alphaCSR[ 32 ][ 5 ],
   alphaCSR[ 32 ][ 6 ],
   alphaCSR[ 32 ][ 7 ],
   alphaCSR[ 32 ][ 8 ],
   alphaCSR[ 32 ][ 9 ],
   alphaCSR[ 32 ][ 10 ],
   alphaCSR[ 32 ][ 11 ],
   alphaCSR[ 32 ][ 12 ],
   alphaCSR[ 32 ][ 13 ],
   alphaCSR[ 32 ][ 14 ],
   alphaCSR[ 32 ][ 15 ],
   alphaCSR[ 32 ][ 16 ],
   alphaCSR[ 32 ][ 17 ],
   alphaCSR[ 32 ][ 18 ],
   alphaCSR[ 32 ][ 19 ],
   alphaCSR[ 32 ][ 20 ],
   alphaCSR[ 32 ][ 21 ],
   alphaCSR[ 32 ][ 22 ],
   alphaCSR[ 32 ][ 23 ],
   alphaCSR[ 32 ][ 24 ],
   alphaCSR[ 32 ][ 25 ],
   alphaCSR[ 32 ][ 26 ],
   alphaCSR[ 32 ][ 27 ],
   alphaCSR[ 32 ][ 28 ],
   alphaCSR[ 32 ][ 29 ],
   alphaCSR[ 32 ][ 30 ],
   alphaCSR[ 32 ][ 31 ],
   alphaCSR[ 32 ][ 32 ],
   alphaCSR[ 32 ][ 33 ],
   alphaCSR[ 32 ][ 34 ],
   alphaCSR[ 32 ][ 35 ],
   alphaCSR[ 32 ][ 36 ],
   alphaCSR[ 32 ][ 37 ],
   alphaCSR[ 32 ][ 38 ],
   alphaCSR[ 32 ][ 39 ],
   alphaCSR[ 32 ][ 40 ],
   alphaCSR[ 32 ][ 41 ],
   alphaCSR[ 32 ][ 42 ],
   alphaCSR[ 32 ][ 43 ],
   alphaCSR[ 32 ][ 44 ],
   alphaCSR[ 32 ][ 45 ],
   alphaCSR[ 32 ][ 46 ],
   alphaCSR[ 32 ][ 47 ],
   alphaCSR[ 32 ][ 48 ],
   alphaCSR[ 32 ][ 49 ],
   alphaCSR[ 32 ][ 50 ],
   alphaCSR[ 32 ][ 51 ],
   alphaCSR[ 32 ][ 52 ],
   alphaCSR[ 32 ][ 53 ],
   alphaCSR[ 32 ][ 54 ],
   alphaCSR[ 32 ][ 55 ],
   alphaCSR[ 32 ][ 56 ],
   alphaCSR[ 32 ][ 57 ],
   alphaCSR[ 32 ][ 58 ],
   alphaCSR[ 32 ][ 59 ],
   alphaCSR[ 32 ][ 60 ],
   alphaCSR[ 32 ][ 61 ],
   alphaCSR[ 32 ][ 62 ],
   alphaCSR[ 32 ][ 63 ],
   alphaCSR[ 32 ][ 64 ],
   alphaCSR[ 32 ][ 65 ],
   alphaCSR[ 32 ][ 66 ],
   alphaCSR[ 32 ][ 67 ],
   alphaCSR[ 32 ][ 68 ],
   alphaCSR[ 32 ][ 69 ],
   alphaCSR[ 32 ][ 70 ],
   alphaCSR[ 32 ][ 71 ],
   alphaCSR[ 32 ][ 72 ],
   alphaCSR[ 32 ][ 73 ],
   alphaCSR[ 32 ][ 74 ],
   alphaCSR[ 32 ][ 75 ],
   alphaCSR[ 32 ][ 76 ],
   alphaCSR[ 32 ][ 77 ],
   alphaCSR[ 32 ][ 78 ],
   alphaCSR[ 32 ][ 79 ],
   alphaCSR[ 32 ][ 80 ],
   alphaCSR[ 32 ][ 81 ],
   alphaCSR[ 32 ][ 82 ],
   alphaCSR[ 32 ][ 83 ],
   alphaCSR[ 32 ][ 84 ],
   alphaCSR[ 32 ][ 85 ],
   alphaCSR[ 32 ][ 86 ],
   alphaCSR[ 32 ][ 87 ],
   alphaCSR[ 32 ][ 88 ],
   alphaCSR[ 32 ][ 89 ],
   alphaCSR[ 32 ][ 90 ],
   alphaCSR[ 32 ][ 91 ],
   alphaCSR[ 32 ][ 92 ],
   alphaCSR[ 32 ][ 93 ],
   alphaCSR[ 32 ][ 94 ],
   alphaCSR[ 32 ][ 95 ],
   alphaCSR[ 32 ][ 96 ],
   alphaCSR[ 32 ][ 97 ],
   alphaCSR[ 32 ][ 98 ],
   alphaCSR[ 32 ][ 99 ],
   alphaCSR[ 32 ][ 100 ],
   alphaCSR[ 32 ][ 101 ],
   alphaCSR[ 32 ][ 102 ],
   alphaCSR[ 32 ][ 103 ],
   alphaCSR[ 32 ][ 104 ],
   alphaCSR[ 32 ][ 105 ],
   alphaCSR[ 32 ][ 106 ],
   alphaCSR[ 32 ][ 107 ],
   alphaCSR[ 32 ][ 108 ],
   alphaCSR[ 32 ][ 109 ],
   alphaCSR[ 32 ][ 110 ],
   alphaCSR[ 32 ][ 111 ],
   alphaCSR[ 32 ][ 112 ],
   alphaCSR[ 32 ][ 113 ],
   alphaCSR[ 32 ][ 114 ],
   alphaCSR[ 32 ][ 115 ],
   alphaCSR[ 32 ][ 116 ],
   alphaCSR[ 32 ][ 117 ],
   alphaCSR[ 32 ][ 118 ],
   alphaCSR[ 32 ][ 119 ],
   alphaCSR[ 32 ][ 120 ],
   alphaCSR[ 32 ][ 121 ],
   alphaCSR[ 32 ][ 122 ],
   alphaCSR[ 32 ][ 123 ],
   alphaCSR[ 32 ][ 124 ],
   alphaCSR[ 32 ][ 125 ],
   alphaCSR[ 32 ][ 126 ],
   alphaCSR[ 32 ][ 127 ],
   alphaCSR[ 32 ][ 128 ],
   alphaCSR[ 32 ][ 129 ],
   alphaCSR[ 32 ][ 130 ],
   alphaCSR[ 32 ][ 131 ],
   alphaCSR[ 32 ][ 132 ],
   alphaCSR[ 32 ][ 133 ],
   alphaCSR[ 32 ][ 134 ],
   alphaCSR[ 32 ][ 135 ],
   alphaCSR[ 32 ][ 136 ],
   alphaCSR[ 32 ][ 137 ],
   alphaCSR[ 32 ][ 138 ],
   alphaCSR[ 32 ][ 139 ],
   alphaCSR[ 32 ][ 140 ],
   alphaCSR[ 32 ][ 141 ],
   alphaCSR[ 32 ][ 142 ],
   alphaCSR[ 32 ][ 143 ],
   alphaCSR[ 32 ][ 144 ],
   alphaCSR[ 32 ][ 145 ],
   alphaCSR[ 32 ][ 146 ],
   alphaCSR[ 32 ][ 147 ],
   alphaCSR[ 32 ][ 148 ],
   alphaCSR[ 32 ][ 149 ],
   alphaCSR[ 32 ][ 150 ],
   alphaCSR[ 32 ][ 151 ],
   alphaCSR[ 32 ][ 152 ],
   alphaCSR[ 32 ][ 153 ],
   alphaCSR[ 32 ][ 154 ],
   alphaCSR[ 32 ][ 155 ],
   alphaCSR[ 32 ][ 156 ],
   alphaCSR[ 32 ][ 157 ],
   alphaCSR[ 32 ][ 158 ],
   alphaCSR[ 32 ][ 159 ],
   alphaCSR[ 32 ][ 160 ],
   alphaCSR[ 32 ][ 161 ],
   alphaCSR[ 32 ][ 162 ],
   alphaCSR[ 32 ][ 163 ],
   alphaCSR[ 32 ][ 164 ],
   alphaCSR[ 32 ][ 165 ],
   alphaCSR[ 32 ][ 166 ],
   alphaCSR[ 32 ][ 167 ],
   alphaCSR[ 32 ][ 168 ],
   alphaCSR[ 32 ][ 169 ],
   alphaCSR[ 32 ][ 170 ],
   alphaCSR[ 32 ][ 171 ],
   alphaCSR[ 32 ][ 172 ],
   alphaCSR[ 32 ][ 173 ],
   alphaCSR[ 32 ][ 174 ],
   alphaCSR[ 32 ][ 175 ],
   alphaCSR[ 32 ][ 176 ],
   alphaCSR[ 32 ][ 177 ],
   alphaCSR[ 32 ][ 178 ],
   alphaCSR[ 32 ][ 179 ],
   alphaCSR[ 32 ][ 180 ],
   alphaCSR[ 32 ][ 181 ],
   alphaCSR[ 32 ][ 182 ],
   alphaCSR[ 32 ][ 183 ],
   alphaCSR[ 32 ][ 184 ],
   alphaCSR[ 32 ][ 185 ],
   alphaCSR[ 32 ][ 186 ],
   alphaCSR[ 32 ][ 187 ],
   alphaCSR[ 32 ][ 188 ],
   alphaCSR[ 32 ][ 189 ],
   alphaCSR[ 32 ][ 190 ],
   alphaCSR[ 32 ][ 191 ],
   alphaCSR[ 32 ][ 192 ],
   alphaCSR[ 32 ][ 193 ],
   alphaCSR[ 32 ][ 194 ],
   alphaCSR[ 32 ][ 195 ],
   alphaCSR[ 32 ][ 196 ],
   alphaCSR[ 32 ][ 197 ],
   alphaCSR[ 32 ][ 198 ],
   alphaCSR[ 32 ][ 199 ],
   alphaCSR[ 32 ][ 200 ],
   alphaCSR[ 32 ][ 201 ],
   alphaCSR[ 32 ][ 202 ],
   alphaCSR[ 32 ][ 203 ],
   alphaCSR[ 32 ][ 204 ],
   alphaCSR[ 32 ][ 205 ],
   alphaCSR[ 32 ][ 206 ],
   alphaCSR[ 32 ][ 207 ],
   alphaCSR[ 32 ][ 208 ],
   alphaCSR[ 32 ][ 209 ],
   alphaCSR[ 32 ][ 210 ],
   alphaCSR[ 32 ][ 211 ],
   alphaCSR[ 32 ][ 212 ],
   alphaCSR[ 32 ][ 213 ],
   alphaCSR[ 32 ][ 214 ],
   alphaCSR[ 32 ][ 215 ],
   alphaCSR[ 32 ][ 216 ],
   alphaCSR[ 32 ][ 217 ],
   alphaCSR[ 32 ][ 218 ],
   alphaCSR[ 32 ][ 219 ],
   alphaCSR[ 32 ][ 220 ],
   alphaCSR[ 32 ][ 221 ],
   alphaCSR[ 32 ][ 222 ],
   alphaCSR[ 32 ][ 223 ],
   alphaCSR[ 32 ][ 224 ],
   alphaCSR[ 32 ][ 225 ],
   alphaCSR[ 32 ][ 226 ],
   alphaCSR[ 32 ][ 227 ],
   alphaCSR[ 32 ][ 228 ],
   alphaCSR[ 32 ][ 229 ],
   alphaCSR[ 32 ][ 230 ],
   alphaCSR[ 32 ][ 231 ],
   alphaCSR[ 32 ][ 232 ],
   alphaCSR[ 32 ][ 233 ],
   alphaCSR[ 32 ][ 234 ],
   alphaCSR[ 32 ][ 235 ],
   alphaCSR[ 32 ][ 236 ],
   alphaCSR[ 32 ][ 237 ],
   alphaCSR[ 32 ][ 238 ],
   alphaCSR[ 32 ][ 239 ],
   alphaCSR[ 32 ][ 240 ],
   alphaCSR[ 32 ][ 241 ],
   alphaCSR[ 32 ][ 242 ],
   alphaCSR[ 32 ][ 243 ],
   alphaCSR[ 32 ][ 244 ],
   alphaCSR[ 32 ][ 245 ],
   alphaCSR[ 32 ][ 246 ],
   alphaCSR[ 32 ][ 247 ],
   alphaCSR[ 32 ][ 248 ],
   alphaCSR[ 32 ][ 249 ],
   alphaCSR[ 32 ][ 250 ],
   alphaCSR[ 32 ][ 251 ],
   alphaCSR[ 32 ][ 252 ],
   alphaCSR[ 32 ][ 253 ],
   alphaCSR[ 32 ][ 254 ],
   alphaCSR[ 32 ][ 255 ],
   alphaCSR[ 32 ][ 256 ],
   alphaCSR[ 32 ][ 257 ],
   alphaCSR[ 32 ][ 258 ],
   alphaCSR[ 32 ][ 259 ],
   alphaCSR[ 32 ][ 260 ],
   alphaCSR[ 32 ][ 261 ],
   alphaCSR[ 32 ][ 262 ],
   alphaCSR[ 32 ][ 263 ],
   alphaCSR[ 32 ][ 264 ],
   alphaCSR[ 32 ][ 265 ],
   alphaCSR[ 32 ][ 266 ],
   alphaCSR[ 32 ][ 267 ],
   alphaCSR[ 32 ][ 268 ],
   alphaCSR[ 32 ][ 269 ],
   alphaCSR[ 32 ][ 270 ],
   alphaCSR[ 32 ][ 271 ],
   alphaCSR[ 32 ][ 272 ],
   alphaCSR[ 32 ][ 273 ],
   alphaCSR[ 32 ][ 274 ],
   alphaCSR[ 32 ][ 275 ],
   alphaCSR[ 32 ][ 276 ],
   alphaCSR[ 32 ][ 277 ],
   alphaCSR[ 32 ][ 278 ],
   alphaCSR[ 32 ][ 279 ],
   alphaCSR[ 32 ][ 280 ],
   alphaCSR[ 32 ][ 281 ],
   alphaCSR[ 32 ][ 282 ],
   alphaCSR[ 32 ][ 283 ],
   alphaCSR[ 32 ][ 284 ],
   alphaCSR[ 32 ][ 285 ],
   alphaCSR[ 32 ][ 286 ],
   alphaCSR[ 32 ][ 287 ],
   alphaCSR[ 32 ][ 288 ],
   alphaCSR[ 32 ][ 289 ],
   alphaCSR[ 32 ][ 290 ],
   alphaCSR[ 32 ][ 291 ],
   alphaCSR[ 32 ][ 292 ],
   alphaCSR[ 32 ][ 293 ],
   alphaCSR[ 32 ][ 294 ],
   alphaCSR[ 32 ][ 295 ],
   alphaCSR[ 32 ][ 296 ],
   alphaCSR[ 32 ][ 297 ],
   alphaCSR[ 32 ][ 298 ],
   alphaCSR[ 32 ][ 299 ],
   alphaCSR[ 32 ][ 300 ],
   alphaCSR[ 32 ][ 301 ],
   alphaCSR[ 32 ][ 302 ],
   alphaCSR[ 32 ][ 303 ],
   alphaCSR[ 32 ][ 304 ],
   alphaCSR[ 32 ][ 305 ],
   alphaCSR[ 32 ][ 306 ],
   alphaCSR[ 32 ][ 307 ],
   alphaCSR[ 32 ][ 308 ],
   alphaCSR[ 32 ][ 309 ],
   alphaCSR[ 32 ][ 310 ],
   alphaCSR[ 32 ][ 311 ],
   alphaCSR[ 32 ][ 312 ],
   alphaCSR[ 32 ][ 313 ],
   alphaCSR[ 32 ][ 314 ],
   alphaCSR[ 32 ][ 315 ],
   alphaCSR[ 32 ][ 316 ],
   alphaCSR[ 32 ][ 317 ],
   alphaCSR[ 32 ][ 318 ],
   alphaCSR[ 32 ][ 319 ],
   alphaCSR[ 32 ][ 320 ],
   alphaCSR[ 32 ][ 321 ],
   alphaCSR[ 32 ][ 322 ],
   alphaCSR[ 32 ][ 323 ],
   alphaCSR[ 32 ][ 324 ],
   alphaCSR[ 32 ][ 325 ],
   alphaCSR[ 32 ][ 326 ],
   alphaCSR[ 32 ][ 327 ],
   alphaCSR[ 32 ][ 328 ],
   alphaCSR[ 32 ][ 329 ],
   alphaCSR[ 32 ][ 330 ],
   alphaCSR[ 32 ][ 331 ],
   alphaCSR[ 32 ][ 332 ],
   alphaCSR[ 32 ][ 333 ],
   alphaCSR[ 32 ][ 334 ],
   alphaCSR[ 32 ][ 335 ],
   alphaCSR[ 32 ][ 336 ],
   alphaCSR[ 32 ][ 337 ],
   alphaCSR[ 32 ][ 338 ],
   alphaCSR[ 32 ][ 339 ],
   alphaCSR[ 32 ][ 340 ],
   alphaCSR[ 32 ][ 341 ],
   alphaCSR[ 32 ][ 342 ],
   alphaCSR[ 32 ][ 343 ],
   alphaCSR[ 32 ][ 344 ],
   alphaCSR[ 32 ][ 345 ],
   alphaCSR[ 32 ][ 346 ],
   alphaCSR[ 32 ][ 347 ],
   alphaCSR[ 32 ][ 348 ],
   alphaCSR[ 32 ][ 349 ],
   alphaCSR[ 32 ][ 350 ],
   alphaCSR[ 32 ][ 351 ],
   alphaCSR[ 32 ][ 352 ],
   alphaCSR[ 32 ][ 353 ],
   alphaCSR[ 32 ][ 354 ],
   alphaCSR[ 32 ][ 355 ],
   alphaCSR[ 32 ][ 356 ],
   alphaCSR[ 32 ][ 357 ],
   alphaCSR[ 32 ][ 358 ],
   alphaCSR[ 32 ][ 359 ],
   alphaCSR[ 32 ][ 360 ],
   alphaCSR[ 32 ][ 361 ],
   alphaCSR[ 32 ][ 362 ],
   alphaCSR[ 32 ][ 363 ],
   alphaCSR[ 32 ][ 364 ],
   alphaCSR[ 32 ][ 365 ],
   alphaCSR[ 32 ][ 366 ],
   alphaCSR[ 32 ][ 367 ],
   alphaCSR[ 32 ][ 368 ],
   alphaCSR[ 32 ][ 369 ],
   alphaCSR[ 32 ][ 370 ],
   alphaCSR[ 32 ][ 371 ],
   alphaCSR[ 32 ][ 372 ],
   alphaCSR[ 32 ][ 373 ],
   alphaCSR[ 32 ][ 374 ],
   alphaCSR[ 32 ][ 375 ],
   alphaCSR[ 32 ][ 376 ],
   alphaCSR[ 32 ][ 377 ],
   alphaCSR[ 32 ][ 378 ],
   alphaCSR[ 32 ][ 379 ],
   alphaCSR[ 32 ][ 380 ],
   alphaCSR[ 32 ][ 381 ],
   alphaCSR[ 32 ][ 382 ],
   alphaCSR[ 32 ][ 383 ],
   alphaCSR[ 33 ][ 0 ],
   alphaCSR[ 33 ][ 1 ],
   alphaCSR[ 33 ][ 2 ],
   alphaCSR[ 33 ][ 3 ],
   alphaCSR[ 33 ][ 4 ],
   alphaCSR[ 33 ][ 5 ],
   alphaCSR[ 33 ][ 6 ],
   alphaCSR[ 33 ][ 7 ],
   alphaCSR[ 33 ][ 8 ],
   alphaCSR[ 33 ][ 9 ],
   alphaCSR[ 33 ][ 10 ],
   alphaCSR[ 33 ][ 11 ],
   alphaCSR[ 33 ][ 12 ],
   alphaCSR[ 33 ][ 13 ],
   alphaCSR[ 33 ][ 14 ],
   alphaCSR[ 33 ][ 15 ],
   alphaCSR[ 33 ][ 16 ],
   alphaCSR[ 33 ][ 17 ],
   alphaCSR[ 33 ][ 18 ],
   alphaCSR[ 33 ][ 19 ],
   alphaCSR[ 33 ][ 20 ],
   alphaCSR[ 33 ][ 21 ],
   alphaCSR[ 33 ][ 22 ],
   alphaCSR[ 33 ][ 23 ],
   alphaCSR[ 33 ][ 24 ],
   alphaCSR[ 33 ][ 25 ],
   alphaCSR[ 33 ][ 26 ],
   alphaCSR[ 33 ][ 27 ],
   alphaCSR[ 33 ][ 28 ],
   alphaCSR[ 33 ][ 29 ],
   alphaCSR[ 33 ][ 30 ],
   alphaCSR[ 33 ][ 31 ],
   alphaCSR[ 33 ][ 32 ],
   alphaCSR[ 33 ][ 33 ],
   alphaCSR[ 33 ][ 34 ],
   alphaCSR[ 33 ][ 35 ],
   alphaCSR[ 33 ][ 36 ],
   alphaCSR[ 33 ][ 37 ],
   alphaCSR[ 33 ][ 38 ],
   alphaCSR[ 33 ][ 39 ],
   alphaCSR[ 33 ][ 40 ],
   alphaCSR[ 33 ][ 41 ],
   alphaCSR[ 33 ][ 42 ],
   alphaCSR[ 33 ][ 43 ],
   alphaCSR[ 33 ][ 44 ],
   alphaCSR[ 33 ][ 45 ],
   alphaCSR[ 33 ][ 46 ],
   alphaCSR[ 33 ][ 47 ],
   alphaCSR[ 33 ][ 48 ],
   alphaCSR[ 33 ][ 49 ],
   alphaCSR[ 33 ][ 50 ],
   alphaCSR[ 33 ][ 51 ],
   alphaCSR[ 33 ][ 52 ],
   alphaCSR[ 33 ][ 53 ],
   alphaCSR[ 33 ][ 54 ],
   alphaCSR[ 33 ][ 55 ],
   alphaCSR[ 33 ][ 56 ],
   alphaCSR[ 33 ][ 57 ],
   alphaCSR[ 33 ][ 58 ],
   alphaCSR[ 33 ][ 59 ],
   alphaCSR[ 33 ][ 60 ],
   alphaCSR[ 33 ][ 61 ],
   alphaCSR[ 33 ][ 62 ],
   alphaCSR[ 33 ][ 63 ],
   alphaCSR[ 33 ][ 64 ],
   alphaCSR[ 33 ][ 65 ],
   alphaCSR[ 33 ][ 66 ],
   alphaCSR[ 33 ][ 67 ],
   alphaCSR[ 33 ][ 68 ],
   alphaCSR[ 33 ][ 69 ],
   alphaCSR[ 33 ][ 70 ],
   alphaCSR[ 33 ][ 71 ],
   alphaCSR[ 33 ][ 72 ],
   alphaCSR[ 33 ][ 73 ],
   alphaCSR[ 33 ][ 74 ],
   alphaCSR[ 33 ][ 75 ],
   alphaCSR[ 33 ][ 76 ],
   alphaCSR[ 33 ][ 77 ],
   alphaCSR[ 33 ][ 78 ],
   alphaCSR[ 33 ][ 79 ],
   alphaCSR[ 33 ][ 80 ],
   alphaCSR[ 33 ][ 81 ],
   alphaCSR[ 33 ][ 82 ],
   alphaCSR[ 33 ][ 83 ],
   alphaCSR[ 33 ][ 84 ],
   alphaCSR[ 33 ][ 85 ],
   alphaCSR[ 33 ][ 86 ],
   alphaCSR[ 33 ][ 87 ],
   alphaCSR[ 33 ][ 88 ],
   alphaCSR[ 33 ][ 89 ],
   alphaCSR[ 33 ][ 90 ],
   alphaCSR[ 33 ][ 91 ],
   alphaCSR[ 33 ][ 92 ],
   alphaCSR[ 33 ][ 93 ],
   alphaCSR[ 33 ][ 94 ],
   alphaCSR[ 33 ][ 95 ],
   alphaCSR[ 33 ][ 96 ],
   alphaCSR[ 33 ][ 97 ],
   alphaCSR[ 33 ][ 98 ],
   alphaCSR[ 33 ][ 99 ],
   alphaCSR[ 33 ][ 100 ],
   alphaCSR[ 33 ][ 101 ],
   alphaCSR[ 33 ][ 102 ],
   alphaCSR[ 33 ][ 103 ],
   alphaCSR[ 33 ][ 104 ],
   alphaCSR[ 33 ][ 105 ],
   alphaCSR[ 33 ][ 106 ],
   alphaCSR[ 33 ][ 107 ],
   alphaCSR[ 33 ][ 108 ],
   alphaCSR[ 33 ][ 109 ],
   alphaCSR[ 33 ][ 110 ],
   alphaCSR[ 33 ][ 111 ],
   alphaCSR[ 33 ][ 112 ],
   alphaCSR[ 33 ][ 113 ],
   alphaCSR[ 33 ][ 114 ],
   alphaCSR[ 33 ][ 115 ],
   alphaCSR[ 33 ][ 116 ],
   alphaCSR[ 33 ][ 117 ],
   alphaCSR[ 33 ][ 118 ],
   alphaCSR[ 33 ][ 119 ],
   alphaCSR[ 33 ][ 120 ],
   alphaCSR[ 33 ][ 121 ],
   alphaCSR[ 33 ][ 122 ],
   alphaCSR[ 33 ][ 123 ],
   alphaCSR[ 33 ][ 124 ],
   alphaCSR[ 33 ][ 125 ],
   alphaCSR[ 33 ][ 126 ],
   alphaCSR[ 33 ][ 127 ],
   alphaCSR[ 33 ][ 128 ],
   alphaCSR[ 33 ][ 129 ],
   alphaCSR[ 33 ][ 130 ],
   alphaCSR[ 33 ][ 131 ],
   alphaCSR[ 33 ][ 132 ],
   alphaCSR[ 33 ][ 133 ],
   alphaCSR[ 33 ][ 134 ],
   alphaCSR[ 33 ][ 135 ],
   alphaCSR[ 33 ][ 136 ],
   alphaCSR[ 33 ][ 137 ],
   alphaCSR[ 33 ][ 138 ],
   alphaCSR[ 33 ][ 139 ],
   alphaCSR[ 33 ][ 140 ],
   alphaCSR[ 33 ][ 141 ],
   alphaCSR[ 33 ][ 142 ],
   alphaCSR[ 33 ][ 143 ],
   alphaCSR[ 33 ][ 144 ],
   alphaCSR[ 33 ][ 145 ],
   alphaCSR[ 33 ][ 146 ],
   alphaCSR[ 33 ][ 147 ],
   alphaCSR[ 33 ][ 148 ],
   alphaCSR[ 33 ][ 149 ],
   alphaCSR[ 33 ][ 150 ],
   alphaCSR[ 33 ][ 151 ],
   alphaCSR[ 33 ][ 152 ],
   alphaCSR[ 33 ][ 153 ],
   alphaCSR[ 33 ][ 154 ],
   alphaCSR[ 33 ][ 155 ],
   alphaCSR[ 33 ][ 156 ],
   alphaCSR[ 33 ][ 157 ],
   alphaCSR[ 33 ][ 158 ],
   alphaCSR[ 33 ][ 159 ],
   alphaCSR[ 33 ][ 160 ],
   alphaCSR[ 33 ][ 161 ],
   alphaCSR[ 33 ][ 162 ],
   alphaCSR[ 33 ][ 163 ],
   alphaCSR[ 33 ][ 164 ],
   alphaCSR[ 33 ][ 165 ],
   alphaCSR[ 33 ][ 166 ],
   alphaCSR[ 33 ][ 167 ],
   alphaCSR[ 33 ][ 168 ],
   alphaCSR[ 33 ][ 169 ],
   alphaCSR[ 33 ][ 170 ],
   alphaCSR[ 33 ][ 171 ],
   alphaCSR[ 33 ][ 172 ],
   alphaCSR[ 33 ][ 173 ],
   alphaCSR[ 33 ][ 174 ],
   alphaCSR[ 33 ][ 175 ],
   alphaCSR[ 33 ][ 176 ],
   alphaCSR[ 33 ][ 177 ],
   alphaCSR[ 33 ][ 178 ],
   alphaCSR[ 33 ][ 179 ],
   alphaCSR[ 33 ][ 180 ],
   alphaCSR[ 33 ][ 181 ],
   alphaCSR[ 33 ][ 182 ],
   alphaCSR[ 33 ][ 183 ],
   alphaCSR[ 33 ][ 184 ],
   alphaCSR[ 33 ][ 185 ],
   alphaCSR[ 33 ][ 186 ],
   alphaCSR[ 33 ][ 187 ],
   alphaCSR[ 33 ][ 188 ],
   alphaCSR[ 33 ][ 189 ],
   alphaCSR[ 33 ][ 190 ],
   alphaCSR[ 33 ][ 191 ],
   alphaCSR[ 33 ][ 192 ],
   alphaCSR[ 33 ][ 193 ],
   alphaCSR[ 33 ][ 194 ],
   alphaCSR[ 33 ][ 195 ],
   alphaCSR[ 33 ][ 196 ],
   alphaCSR[ 33 ][ 197 ],
   alphaCSR[ 33 ][ 198 ],
   alphaCSR[ 33 ][ 199 ],
   alphaCSR[ 33 ][ 200 ],
   alphaCSR[ 33 ][ 201 ],
   alphaCSR[ 33 ][ 202 ],
   alphaCSR[ 33 ][ 203 ],
   alphaCSR[ 33 ][ 204 ],
   alphaCSR[ 33 ][ 205 ],
   alphaCSR[ 33 ][ 206 ],
   alphaCSR[ 33 ][ 207 ],
   alphaCSR[ 33 ][ 208 ],
   alphaCSR[ 33 ][ 209 ],
   alphaCSR[ 33 ][ 210 ],
   alphaCSR[ 33 ][ 211 ],
   alphaCSR[ 33 ][ 212 ],
   alphaCSR[ 33 ][ 213 ],
   alphaCSR[ 33 ][ 214 ],
   alphaCSR[ 33 ][ 215 ],
   alphaCSR[ 33 ][ 216 ],
   alphaCSR[ 33 ][ 217 ],
   alphaCSR[ 33 ][ 218 ],
   alphaCSR[ 33 ][ 219 ],
   alphaCSR[ 33 ][ 220 ],
   alphaCSR[ 33 ][ 221 ],
   alphaCSR[ 33 ][ 222 ],
   alphaCSR[ 33 ][ 223 ],
   alphaCSR[ 33 ][ 224 ],
   alphaCSR[ 33 ][ 225 ],
   alphaCSR[ 33 ][ 226 ],
   alphaCSR[ 33 ][ 227 ],
   alphaCSR[ 33 ][ 228 ],
   alphaCSR[ 33 ][ 229 ],
   alphaCSR[ 33 ][ 230 ],
   alphaCSR[ 33 ][ 231 ],
   alphaCSR[ 33 ][ 232 ],
   alphaCSR[ 33 ][ 233 ],
   alphaCSR[ 33 ][ 234 ],
   alphaCSR[ 33 ][ 235 ],
   alphaCSR[ 33 ][ 236 ],
   alphaCSR[ 33 ][ 237 ],
   alphaCSR[ 33 ][ 238 ],
   alphaCSR[ 33 ][ 239 ],
   alphaCSR[ 33 ][ 240 ],
   alphaCSR[ 33 ][ 241 ],
   alphaCSR[ 33 ][ 242 ],
   alphaCSR[ 33 ][ 243 ],
   alphaCSR[ 33 ][ 244 ],
   alphaCSR[ 33 ][ 245 ],
   alphaCSR[ 33 ][ 246 ],
   alphaCSR[ 33 ][ 247 ],
   alphaCSR[ 33 ][ 248 ],
   alphaCSR[ 33 ][ 249 ],
   alphaCSR[ 33 ][ 250 ],
   alphaCSR[ 33 ][ 251 ],
   alphaCSR[ 33 ][ 252 ],
   alphaCSR[ 33 ][ 253 ],
   alphaCSR[ 33 ][ 254 ],
   alphaCSR[ 33 ][ 255 ],
   alphaCSR[ 33 ][ 256 ],
   alphaCSR[ 33 ][ 257 ],
   alphaCSR[ 33 ][ 258 ],
   alphaCSR[ 33 ][ 259 ],
   alphaCSR[ 33 ][ 260 ],
   alphaCSR[ 33 ][ 261 ],
   alphaCSR[ 33 ][ 262 ],
   alphaCSR[ 33 ][ 263 ],
   alphaCSR[ 33 ][ 264 ],
   alphaCSR[ 33 ][ 265 ],
   alphaCSR[ 33 ][ 266 ],
   alphaCSR[ 33 ][ 267 ],
   alphaCSR[ 33 ][ 268 ],
   alphaCSR[ 33 ][ 269 ],
   alphaCSR[ 33 ][ 270 ],
   alphaCSR[ 33 ][ 271 ],
   alphaCSR[ 33 ][ 272 ],
   alphaCSR[ 33 ][ 273 ],
   alphaCSR[ 33 ][ 274 ],
   alphaCSR[ 33 ][ 275 ],
   alphaCSR[ 33 ][ 276 ],
   alphaCSR[ 33 ][ 277 ],
   alphaCSR[ 33 ][ 278 ],
   alphaCSR[ 33 ][ 279 ],
   alphaCSR[ 33 ][ 280 ],
   alphaCSR[ 33 ][ 281 ],
   alphaCSR[ 33 ][ 282 ],
   alphaCSR[ 33 ][ 283 ],
   alphaCSR[ 33 ][ 284 ],
   alphaCSR[ 33 ][ 285 ],
   alphaCSR[ 33 ][ 286 ],
   alphaCSR[ 33 ][ 287 ],
   alphaCSR[ 33 ][ 288 ],
   alphaCSR[ 33 ][ 289 ],
   alphaCSR[ 33 ][ 290 ],
   alphaCSR[ 33 ][ 291 ],
   alphaCSR[ 33 ][ 292 ],
   alphaCSR[ 33 ][ 293 ],
   alphaCSR[ 33 ][ 294 ],
   alphaCSR[ 33 ][ 295 ],
   alphaCSR[ 33 ][ 296 ],
   alphaCSR[ 33 ][ 297 ],
   alphaCSR[ 33 ][ 298 ],
   alphaCSR[ 33 ][ 299 ],
   alphaCSR[ 33 ][ 300 ],
   alphaCSR[ 33 ][ 301 ],
   alphaCSR[ 33 ][ 302 ],
   alphaCSR[ 33 ][ 303 ],
   alphaCSR[ 33 ][ 304 ],
   alphaCSR[ 33 ][ 305 ],
   alphaCSR[ 33 ][ 306 ],
   alphaCSR[ 33 ][ 307 ],
   alphaCSR[ 33 ][ 308 ],
   alphaCSR[ 33 ][ 309 ],
   alphaCSR[ 33 ][ 310 ],
   alphaCSR[ 33 ][ 311 ],
   alphaCSR[ 33 ][ 312 ],
   alphaCSR[ 33 ][ 313 ],
   alphaCSR[ 33 ][ 314 ],
   alphaCSR[ 33 ][ 315 ],
   alphaCSR[ 33 ][ 316 ],
   alphaCSR[ 33 ][ 317 ],
   alphaCSR[ 33 ][ 318 ],
   alphaCSR[ 33 ][ 319 ],
   alphaCSR[ 33 ][ 320 ],
   alphaCSR[ 33 ][ 321 ],
   alphaCSR[ 33 ][ 322 ],
   alphaCSR[ 33 ][ 323 ],
   alphaCSR[ 33 ][ 324 ],
   alphaCSR[ 33 ][ 325 ],
   alphaCSR[ 33 ][ 326 ],
   alphaCSR[ 33 ][ 327 ],
   alphaCSR[ 33 ][ 328 ],
   alphaCSR[ 33 ][ 329 ],
   alphaCSR[ 33 ][ 330 ],
   alphaCSR[ 33 ][ 331 ],
   alphaCSR[ 33 ][ 332 ],
   alphaCSR[ 33 ][ 333 ],
   alphaCSR[ 33 ][ 334 ],
   alphaCSR[ 33 ][ 335 ],
   alphaCSR[ 33 ][ 336 ],
   alphaCSR[ 33 ][ 337 ],
   alphaCSR[ 33 ][ 338 ],
   alphaCSR[ 33 ][ 339 ],
   alphaCSR[ 33 ][ 340 ],
   alphaCSR[ 33 ][ 341 ],
   alphaCSR[ 33 ][ 342 ],
   alphaCSR[ 33 ][ 343 ],
   alphaCSR[ 33 ][ 344 ],
   alphaCSR[ 33 ][ 345 ],
   alphaCSR[ 33 ][ 346 ],
   alphaCSR[ 33 ][ 347 ],
   alphaCSR[ 33 ][ 348 ],
   alphaCSR[ 33 ][ 349 ],
   alphaCSR[ 33 ][ 350 ],
   alphaCSR[ 33 ][ 351 ],
   alphaCSR[ 33 ][ 352 ],
   alphaCSR[ 33 ][ 353 ],
   alphaCSR[ 33 ][ 354 ],
   alphaCSR[ 33 ][ 355 ],
   alphaCSR[ 33 ][ 356 ],
   alphaCSR[ 33 ][ 357 ],
   alphaCSR[ 33 ][ 358 ],
   alphaCSR[ 33 ][ 359 ],
   alphaCSR[ 33 ][ 360 ],
   alphaCSR[ 33 ][ 361 ],
   alphaCSR[ 33 ][ 362 ],
   alphaCSR[ 33 ][ 363 ],
   alphaCSR[ 33 ][ 364 ],
   alphaCSR[ 33 ][ 365 ],
   alphaCSR[ 33 ][ 366 ],
   alphaCSR[ 33 ][ 367 ],
   alphaCSR[ 33 ][ 368 ],
   alphaCSR[ 33 ][ 369 ],
   alphaCSR[ 33 ][ 370 ],
   alphaCSR[ 33 ][ 371 ],
   alphaCSR[ 33 ][ 372 ],
   alphaCSR[ 33 ][ 373 ],
   alphaCSR[ 33 ][ 374 ],
   alphaCSR[ 33 ][ 375 ],
   alphaCSR[ 33 ][ 376 ],
   alphaCSR[ 33 ][ 377 ],
   alphaCSR[ 33 ][ 378 ],
   alphaCSR[ 33 ][ 379 ],
   alphaCSR[ 33 ][ 380 ],
   alphaCSR[ 33 ][ 381 ],
   alphaCSR[ 33 ][ 382 ],
   alphaCSR[ 33 ][ 383 ],
   alphaCSR[ 34 ][ 0 ],
   alphaCSR[ 34 ][ 1 ],
   alphaCSR[ 34 ][ 2 ],
   alphaCSR[ 34 ][ 3 ],
   alphaCSR[ 34 ][ 4 ],
   alphaCSR[ 34 ][ 5 ],
   alphaCSR[ 34 ][ 6 ],
   alphaCSR[ 34 ][ 7 ],
   alphaCSR[ 34 ][ 8 ],
   alphaCSR[ 34 ][ 9 ],
   alphaCSR[ 34 ][ 10 ],
   alphaCSR[ 34 ][ 11 ],
   alphaCSR[ 34 ][ 12 ],
   alphaCSR[ 34 ][ 13 ],
   alphaCSR[ 34 ][ 14 ],
   alphaCSR[ 34 ][ 15 ],
   alphaCSR[ 34 ][ 16 ],
   alphaCSR[ 34 ][ 17 ],
   alphaCSR[ 34 ][ 18 ],
   alphaCSR[ 34 ][ 19 ],
   alphaCSR[ 34 ][ 20 ],
   alphaCSR[ 34 ][ 21 ],
   alphaCSR[ 34 ][ 22 ],
   alphaCSR[ 34 ][ 23 ],
   alphaCSR[ 34 ][ 24 ],
   alphaCSR[ 34 ][ 25 ],
   alphaCSR[ 34 ][ 26 ],
   alphaCSR[ 34 ][ 27 ],
   alphaCSR[ 34 ][ 28 ],
   alphaCSR[ 34 ][ 29 ],
   alphaCSR[ 34 ][ 30 ],
   alphaCSR[ 34 ][ 31 ],
   alphaCSR[ 34 ][ 32 ],
   alphaCSR[ 34 ][ 33 ],
   alphaCSR[ 34 ][ 34 ],
   alphaCSR[ 34 ][ 35 ],
   alphaCSR[ 34 ][ 36 ],
   alphaCSR[ 34 ][ 37 ],
   alphaCSR[ 34 ][ 38 ],
   alphaCSR[ 34 ][ 39 ],
   alphaCSR[ 34 ][ 40 ],
   alphaCSR[ 34 ][ 41 ],
   alphaCSR[ 34 ][ 42 ],
   alphaCSR[ 34 ][ 43 ],
   alphaCSR[ 34 ][ 44 ],
   alphaCSR[ 34 ][ 45 ],
   alphaCSR[ 34 ][ 46 ],
   alphaCSR[ 34 ][ 47 ],
   alphaCSR[ 34 ][ 48 ],
   alphaCSR[ 34 ][ 49 ],
   alphaCSR[ 34 ][ 50 ],
   alphaCSR[ 34 ][ 51 ],
   alphaCSR[ 34 ][ 52 ],
   alphaCSR[ 34 ][ 53 ],
   alphaCSR[ 34 ][ 54 ],
   alphaCSR[ 34 ][ 55 ],
   alphaCSR[ 34 ][ 56 ],
   alphaCSR[ 34 ][ 57 ],
   alphaCSR[ 34 ][ 58 ],
   alphaCSR[ 34 ][ 59 ],
   alphaCSR[ 34 ][ 60 ],
   alphaCSR[ 34 ][ 61 ],
   alphaCSR[ 34 ][ 62 ],
   alphaCSR[ 34 ][ 63 ],
   alphaCSR[ 34 ][ 64 ],
   alphaCSR[ 34 ][ 65 ],
   alphaCSR[ 34 ][ 66 ],
   alphaCSR[ 34 ][ 67 ],
   alphaCSR[ 34 ][ 68 ],
   alphaCSR[ 34 ][ 69 ],
   alphaCSR[ 34 ][ 70 ],
   alphaCSR[ 34 ][ 71 ],
   alphaCSR[ 34 ][ 72 ],
   alphaCSR[ 34 ][ 73 ],
   alphaCSR[ 34 ][ 74 ],
   alphaCSR[ 34 ][ 75 ],
   alphaCSR[ 34 ][ 76 ],
   alphaCSR[ 34 ][ 77 ],
   alphaCSR[ 34 ][ 78 ],
   alphaCSR[ 34 ][ 79 ],
   alphaCSR[ 34 ][ 80 ],
   alphaCSR[ 34 ][ 81 ],
   alphaCSR[ 34 ][ 82 ],
   alphaCSR[ 34 ][ 83 ],
   alphaCSR[ 34 ][ 84 ],
   alphaCSR[ 34 ][ 85 ],
   alphaCSR[ 34 ][ 86 ],
   alphaCSR[ 34 ][ 87 ],
   alphaCSR[ 34 ][ 88 ],
   alphaCSR[ 34 ][ 89 ],
   alphaCSR[ 34 ][ 90 ],
   alphaCSR[ 34 ][ 91 ],
   alphaCSR[ 34 ][ 92 ],
   alphaCSR[ 34 ][ 93 ],
   alphaCSR[ 34 ][ 94 ],
   alphaCSR[ 34 ][ 95 ],
   alphaCSR[ 34 ][ 96 ],
   alphaCSR[ 34 ][ 97 ],
   alphaCSR[ 34 ][ 98 ],
   alphaCSR[ 34 ][ 99 ],
   alphaCSR[ 34 ][ 100 ],
   alphaCSR[ 34 ][ 101 ],
   alphaCSR[ 34 ][ 102 ],
   alphaCSR[ 34 ][ 103 ],
   alphaCSR[ 34 ][ 104 ],
   alphaCSR[ 34 ][ 105 ],
   alphaCSR[ 34 ][ 106 ],
   alphaCSR[ 34 ][ 107 ],
   alphaCSR[ 34 ][ 108 ],
   alphaCSR[ 34 ][ 109 ],
   alphaCSR[ 34 ][ 110 ],
   alphaCSR[ 34 ][ 111 ],
   alphaCSR[ 34 ][ 112 ],
   alphaCSR[ 34 ][ 113 ],
   alphaCSR[ 34 ][ 114 ],
   alphaCSR[ 34 ][ 115 ],
   alphaCSR[ 34 ][ 116 ],
   alphaCSR[ 34 ][ 117 ],
   alphaCSR[ 34 ][ 118 ],
   alphaCSR[ 34 ][ 119 ],
   alphaCSR[ 34 ][ 120 ],
   alphaCSR[ 34 ][ 121 ],
   alphaCSR[ 34 ][ 122 ],
   alphaCSR[ 34 ][ 123 ],
   alphaCSR[ 34 ][ 124 ],
   alphaCSR[ 34 ][ 125 ],
   alphaCSR[ 34 ][ 126 ],
   alphaCSR[ 34 ][ 127 ],
   alphaCSR[ 34 ][ 128 ],
   alphaCSR[ 34 ][ 129 ],
   alphaCSR[ 34 ][ 130 ],
   alphaCSR[ 34 ][ 131 ],
   alphaCSR[ 34 ][ 132 ],
   alphaCSR[ 34 ][ 133 ],
   alphaCSR[ 34 ][ 134 ],
   alphaCSR[ 34 ][ 135 ],
   alphaCSR[ 34 ][ 136 ],
   alphaCSR[ 34 ][ 137 ],
   alphaCSR[ 34 ][ 138 ],
   alphaCSR[ 34 ][ 139 ],
   alphaCSR[ 34 ][ 140 ],
   alphaCSR[ 34 ][ 141 ],
   alphaCSR[ 34 ][ 142 ],
   alphaCSR[ 34 ][ 143 ],
   alphaCSR[ 34 ][ 144 ],
   alphaCSR[ 34 ][ 145 ],
   alphaCSR[ 34 ][ 146 ],
   alphaCSR[ 34 ][ 147 ],
   alphaCSR[ 34 ][ 148 ],
   alphaCSR[ 34 ][ 149 ],
   alphaCSR[ 34 ][ 150 ],
   alphaCSR[ 34 ][ 151 ],
   alphaCSR[ 34 ][ 152 ],
   alphaCSR[ 34 ][ 153 ],
   alphaCSR[ 34 ][ 154 ],
   alphaCSR[ 34 ][ 155 ],
   alphaCSR[ 34 ][ 156 ],
   alphaCSR[ 34 ][ 157 ],
   alphaCSR[ 34 ][ 158 ],
   alphaCSR[ 34 ][ 159 ],
   alphaCSR[ 34 ][ 160 ],
   alphaCSR[ 34 ][ 161 ],
   alphaCSR[ 34 ][ 162 ],
   alphaCSR[ 34 ][ 163 ],
   alphaCSR[ 34 ][ 164 ],
   alphaCSR[ 34 ][ 165 ],
   alphaCSR[ 34 ][ 166 ],
   alphaCSR[ 34 ][ 167 ],
   alphaCSR[ 34 ][ 168 ],
   alphaCSR[ 34 ][ 169 ],
   alphaCSR[ 34 ][ 170 ],
   alphaCSR[ 34 ][ 171 ],
   alphaCSR[ 34 ][ 172 ],
   alphaCSR[ 34 ][ 173 ],
   alphaCSR[ 34 ][ 174 ],
   alphaCSR[ 34 ][ 175 ],
   alphaCSR[ 34 ][ 176 ],
   alphaCSR[ 34 ][ 177 ],
   alphaCSR[ 34 ][ 178 ],
   alphaCSR[ 34 ][ 179 ],
   alphaCSR[ 34 ][ 180 ],
   alphaCSR[ 34 ][ 181 ],
   alphaCSR[ 34 ][ 182 ],
   alphaCSR[ 34 ][ 183 ],
   alphaCSR[ 34 ][ 184 ],
   alphaCSR[ 34 ][ 185 ],
   alphaCSR[ 34 ][ 186 ],
   alphaCSR[ 34 ][ 187 ],
   alphaCSR[ 34 ][ 188 ],
   alphaCSR[ 34 ][ 189 ],
   alphaCSR[ 34 ][ 190 ],
   alphaCSR[ 34 ][ 191 ],
   alphaCSR[ 34 ][ 192 ],
   alphaCSR[ 34 ][ 193 ],
   alphaCSR[ 34 ][ 194 ],
   alphaCSR[ 34 ][ 195 ],
   alphaCSR[ 34 ][ 196 ],
   alphaCSR[ 34 ][ 197 ],
   alphaCSR[ 34 ][ 198 ],
   alphaCSR[ 34 ][ 199 ],
   alphaCSR[ 34 ][ 200 ],
   alphaCSR[ 34 ][ 201 ],
   alphaCSR[ 34 ][ 202 ],
   alphaCSR[ 34 ][ 203 ],
   alphaCSR[ 34 ][ 204 ],
   alphaCSR[ 34 ][ 205 ],
   alphaCSR[ 34 ][ 206 ],
   alphaCSR[ 34 ][ 207 ],
   alphaCSR[ 34 ][ 208 ],
   alphaCSR[ 34 ][ 209 ],
   alphaCSR[ 34 ][ 210 ],
   alphaCSR[ 34 ][ 211 ],
   alphaCSR[ 34 ][ 212 ],
   alphaCSR[ 34 ][ 213 ],
   alphaCSR[ 34 ][ 214 ],
   alphaCSR[ 34 ][ 215 ],
   alphaCSR[ 34 ][ 216 ],
   alphaCSR[ 34 ][ 217 ],
   alphaCSR[ 34 ][ 218 ],
   alphaCSR[ 34 ][ 219 ],
   alphaCSR[ 34 ][ 220 ],
   alphaCSR[ 34 ][ 221 ],
   alphaCSR[ 34 ][ 222 ],
   alphaCSR[ 34 ][ 223 ],
   alphaCSR[ 34 ][ 224 ],
   alphaCSR[ 34 ][ 225 ],
   alphaCSR[ 34 ][ 226 ],
   alphaCSR[ 34 ][ 227 ],
   alphaCSR[ 34 ][ 228 ],
   alphaCSR[ 34 ][ 229 ],
   alphaCSR[ 34 ][ 230 ],
   alphaCSR[ 34 ][ 231 ],
   alphaCSR[ 34 ][ 232 ],
   alphaCSR[ 34 ][ 233 ],
   alphaCSR[ 34 ][ 234 ],
   alphaCSR[ 34 ][ 235 ],
   alphaCSR[ 34 ][ 236 ],
   alphaCSR[ 34 ][ 237 ],
   alphaCSR[ 34 ][ 238 ],
   alphaCSR[ 34 ][ 239 ],
   alphaCSR[ 34 ][ 240 ],
   alphaCSR[ 34 ][ 241 ],
   alphaCSR[ 34 ][ 242 ],
   alphaCSR[ 34 ][ 243 ],
   alphaCSR[ 34 ][ 244 ],
   alphaCSR[ 34 ][ 245 ],
   alphaCSR[ 34 ][ 246 ],
   alphaCSR[ 34 ][ 247 ],
   alphaCSR[ 34 ][ 248 ],
   alphaCSR[ 34 ][ 249 ],
   alphaCSR[ 34 ][ 250 ],
   alphaCSR[ 34 ][ 251 ],
   alphaCSR[ 34 ][ 252 ],
   alphaCSR[ 34 ][ 253 ],
   alphaCSR[ 34 ][ 254 ],
   alphaCSR[ 34 ][ 255 ],
   alphaCSR[ 34 ][ 256 ],
   alphaCSR[ 34 ][ 257 ],
   alphaCSR[ 34 ][ 258 ],
   alphaCSR[ 34 ][ 259 ],
   alphaCSR[ 34 ][ 260 ],
   alphaCSR[ 34 ][ 261 ],
   alphaCSR[ 34 ][ 262 ],
   alphaCSR[ 34 ][ 263 ],
   alphaCSR[ 34 ][ 264 ],
   alphaCSR[ 34 ][ 265 ],
   alphaCSR[ 34 ][ 266 ],
   alphaCSR[ 34 ][ 267 ],
   alphaCSR[ 34 ][ 268 ],
   alphaCSR[ 34 ][ 269 ],
   alphaCSR[ 34 ][ 270 ],
   alphaCSR[ 34 ][ 271 ],
   alphaCSR[ 34 ][ 272 ],
   alphaCSR[ 34 ][ 273 ],
   alphaCSR[ 34 ][ 274 ],
   alphaCSR[ 34 ][ 275 ],
   alphaCSR[ 34 ][ 276 ],
   alphaCSR[ 34 ][ 277 ],
   alphaCSR[ 34 ][ 278 ],
   alphaCSR[ 34 ][ 279 ],
   alphaCSR[ 34 ][ 280 ],
   alphaCSR[ 34 ][ 281 ],
   alphaCSR[ 34 ][ 282 ],
   alphaCSR[ 34 ][ 283 ],
   alphaCSR[ 34 ][ 284 ],
   alphaCSR[ 34 ][ 285 ],
   alphaCSR[ 34 ][ 286 ],
   alphaCSR[ 34 ][ 287 ],
   alphaCSR[ 34 ][ 288 ],
   alphaCSR[ 34 ][ 289 ],
   alphaCSR[ 34 ][ 290 ],
   alphaCSR[ 34 ][ 291 ],
   alphaCSR[ 34 ][ 292 ],
   alphaCSR[ 34 ][ 293 ],
   alphaCSR[ 34 ][ 294 ],
   alphaCSR[ 34 ][ 295 ],
   alphaCSR[ 34 ][ 296 ],
   alphaCSR[ 34 ][ 297 ],
   alphaCSR[ 34 ][ 298 ],
   alphaCSR[ 34 ][ 299 ],
   alphaCSR[ 34 ][ 300 ],
   alphaCSR[ 34 ][ 301 ],
   alphaCSR[ 34 ][ 302 ],
   alphaCSR[ 34 ][ 303 ],
   alphaCSR[ 34 ][ 304 ],
   alphaCSR[ 34 ][ 305 ],
   alphaCSR[ 34 ][ 306 ],
   alphaCSR[ 34 ][ 307 ],
   alphaCSR[ 34 ][ 308 ],
   alphaCSR[ 34 ][ 309 ],
   alphaCSR[ 34 ][ 310 ],
   alphaCSR[ 34 ][ 311 ],
   alphaCSR[ 34 ][ 312 ],
   alphaCSR[ 34 ][ 313 ],
   alphaCSR[ 34 ][ 314 ],
   alphaCSR[ 34 ][ 315 ],
   alphaCSR[ 34 ][ 316 ],
   alphaCSR[ 34 ][ 317 ],
   alphaCSR[ 34 ][ 318 ],
   alphaCSR[ 34 ][ 319 ],
   alphaCSR[ 34 ][ 320 ],
   alphaCSR[ 34 ][ 321 ],
   alphaCSR[ 34 ][ 322 ],
   alphaCSR[ 34 ][ 323 ],
   alphaCSR[ 34 ][ 324 ],
   alphaCSR[ 34 ][ 325 ],
   alphaCSR[ 34 ][ 326 ],
   alphaCSR[ 34 ][ 327 ],
   alphaCSR[ 34 ][ 328 ],
   alphaCSR[ 34 ][ 329 ],
   alphaCSR[ 34 ][ 330 ],
   alphaCSR[ 34 ][ 331 ],
   alphaCSR[ 34 ][ 332 ],
   alphaCSR[ 34 ][ 333 ],
   alphaCSR[ 34 ][ 334 ],
   alphaCSR[ 34 ][ 335 ],
   alphaCSR[ 34 ][ 336 ],
   alphaCSR[ 34 ][ 337 ],
   alphaCSR[ 34 ][ 338 ],
   alphaCSR[ 34 ][ 339 ],
   alphaCSR[ 34 ][ 340 ],
   alphaCSR[ 34 ][ 341 ],
   alphaCSR[ 34 ][ 342 ],
   alphaCSR[ 34 ][ 343 ],
   alphaCSR[ 34 ][ 344 ],
   alphaCSR[ 34 ][ 345 ],
   alphaCSR[ 34 ][ 346 ],
   alphaCSR[ 34 ][ 347 ],
   alphaCSR[ 34 ][ 348 ],
   alphaCSR[ 34 ][ 349 ],
   alphaCSR[ 34 ][ 350 ],
   alphaCSR[ 34 ][ 351 ],
   alphaCSR[ 34 ][ 352 ],
   alphaCSR[ 34 ][ 353 ],
   alphaCSR[ 34 ][ 354 ],
   alphaCSR[ 34 ][ 355 ],
   alphaCSR[ 34 ][ 356 ],
   alphaCSR[ 34 ][ 357 ],
   alphaCSR[ 34 ][ 358 ],
   alphaCSR[ 34 ][ 359 ],
   alphaCSR[ 34 ][ 360 ],
   alphaCSR[ 34 ][ 361 ],
   alphaCSR[ 34 ][ 362 ],
   alphaCSR[ 34 ][ 363 ],
   alphaCSR[ 34 ][ 364 ],
   alphaCSR[ 34 ][ 365 ],
   alphaCSR[ 34 ][ 366 ],
   alphaCSR[ 34 ][ 367 ],
   alphaCSR[ 34 ][ 368 ],
   alphaCSR[ 34 ][ 369 ],
   alphaCSR[ 34 ][ 370 ],
   alphaCSR[ 34 ][ 371 ],
   alphaCSR[ 34 ][ 372 ],
   alphaCSR[ 34 ][ 373 ],
   alphaCSR[ 34 ][ 374 ],
   alphaCSR[ 34 ][ 375 ],
   alphaCSR[ 34 ][ 376 ],
   alphaCSR[ 34 ][ 377 ],
   alphaCSR[ 34 ][ 378 ],
   alphaCSR[ 34 ][ 379 ],
   alphaCSR[ 34 ][ 380 ],
   alphaCSR[ 34 ][ 381 ],
   alphaCSR[ 34 ][ 382 ],
   alphaCSR[ 34 ][ 383 ],
   alphaCSR[ 35 ][ 0 ],
   alphaCSR[ 35 ][ 1 ],
   alphaCSR[ 35 ][ 2 ],
   alphaCSR[ 35 ][ 3 ],
   alphaCSR[ 35 ][ 4 ],
   alphaCSR[ 35 ][ 5 ],
   alphaCSR[ 35 ][ 6 ],
   alphaCSR[ 35 ][ 7 ],
   alphaCSR[ 35 ][ 8 ],
   alphaCSR[ 35 ][ 9 ],
   alphaCSR[ 35 ][ 10 ],
   alphaCSR[ 35 ][ 11 ],
   alphaCSR[ 35 ][ 12 ],
   alphaCSR[ 35 ][ 13 ],
   alphaCSR[ 35 ][ 14 ],
   alphaCSR[ 35 ][ 15 ],
   alphaCSR[ 35 ][ 16 ],
   alphaCSR[ 35 ][ 17 ],
   alphaCSR[ 35 ][ 18 ],
   alphaCSR[ 35 ][ 19 ],
   alphaCSR[ 35 ][ 20 ],
   alphaCSR[ 35 ][ 21 ],
   alphaCSR[ 35 ][ 22 ],
   alphaCSR[ 35 ][ 23 ],
   alphaCSR[ 35 ][ 24 ],
   alphaCSR[ 35 ][ 25 ],
   alphaCSR[ 35 ][ 26 ],
   alphaCSR[ 35 ][ 27 ],
   alphaCSR[ 35 ][ 28 ],
   alphaCSR[ 35 ][ 29 ],
   alphaCSR[ 35 ][ 30 ],
   alphaCSR[ 35 ][ 31 ],
   alphaCSR[ 35 ][ 32 ],
   alphaCSR[ 35 ][ 33 ],
   alphaCSR[ 35 ][ 34 ],
   alphaCSR[ 35 ][ 35 ],
   alphaCSR[ 35 ][ 36 ],
   alphaCSR[ 35 ][ 37 ],
   alphaCSR[ 35 ][ 38 ],
   alphaCSR[ 35 ][ 39 ],
   alphaCSR[ 35 ][ 40 ],
   alphaCSR[ 35 ][ 41 ],
   alphaCSR[ 35 ][ 42 ],
   alphaCSR[ 35 ][ 43 ],
   alphaCSR[ 35 ][ 44 ],
   alphaCSR[ 35 ][ 45 ],
   alphaCSR[ 35 ][ 46 ],
   alphaCSR[ 35 ][ 47 ],
   alphaCSR[ 35 ][ 48 ],
   alphaCSR[ 35 ][ 49 ],
   alphaCSR[ 35 ][ 50 ],
   alphaCSR[ 35 ][ 51 ],
   alphaCSR[ 35 ][ 52 ],
   alphaCSR[ 35 ][ 53 ],
   alphaCSR[ 35 ][ 54 ],
   alphaCSR[ 35 ][ 55 ],
   alphaCSR[ 35 ][ 56 ],
   alphaCSR[ 35 ][ 57 ],
   alphaCSR[ 35 ][ 58 ],
   alphaCSR[ 35 ][ 59 ],
   alphaCSR[ 35 ][ 60 ],
   alphaCSR[ 35 ][ 61 ],
   alphaCSR[ 35 ][ 62 ],
   alphaCSR[ 35 ][ 63 ],
   alphaCSR[ 35 ][ 64 ],
   alphaCSR[ 35 ][ 65 ],
   alphaCSR[ 35 ][ 66 ],
   alphaCSR[ 35 ][ 67 ],
   alphaCSR[ 35 ][ 68 ],
   alphaCSR[ 35 ][ 69 ],
   alphaCSR[ 35 ][ 70 ],
   alphaCSR[ 35 ][ 71 ],
   alphaCSR[ 35 ][ 72 ],
   alphaCSR[ 35 ][ 73 ],
   alphaCSR[ 35 ][ 74 ],
   alphaCSR[ 35 ][ 75 ],
   alphaCSR[ 35 ][ 76 ],
   alphaCSR[ 35 ][ 77 ],
   alphaCSR[ 35 ][ 78 ],
   alphaCSR[ 35 ][ 79 ],
   alphaCSR[ 35 ][ 80 ],
   alphaCSR[ 35 ][ 81 ],
   alphaCSR[ 35 ][ 82 ],
   alphaCSR[ 35 ][ 83 ],
   alphaCSR[ 35 ][ 84 ],
   alphaCSR[ 35 ][ 85 ],
   alphaCSR[ 35 ][ 86 ],
   alphaCSR[ 35 ][ 87 ],
   alphaCSR[ 35 ][ 88 ],
   alphaCSR[ 35 ][ 89 ],
   alphaCSR[ 35 ][ 90 ],
   alphaCSR[ 35 ][ 91 ],
   alphaCSR[ 35 ][ 92 ],
   alphaCSR[ 35 ][ 93 ],
   alphaCSR[ 35 ][ 94 ],
   alphaCSR[ 35 ][ 95 ],
   alphaCSR[ 35 ][ 96 ],
   alphaCSR[ 35 ][ 97 ],
   alphaCSR[ 35 ][ 98 ],
   alphaCSR[ 35 ][ 99 ],
   alphaCSR[ 35 ][ 100 ],
   alphaCSR[ 35 ][ 101 ],
   alphaCSR[ 35 ][ 102 ],
   alphaCSR[ 35 ][ 103 ],
   alphaCSR[ 35 ][ 104 ],
   alphaCSR[ 35 ][ 105 ],
   alphaCSR[ 35 ][ 106 ],
   alphaCSR[ 35 ][ 107 ],
   alphaCSR[ 35 ][ 108 ],
   alphaCSR[ 35 ][ 109 ],
   alphaCSR[ 35 ][ 110 ],
   alphaCSR[ 35 ][ 111 ],
   alphaCSR[ 35 ][ 112 ],
   alphaCSR[ 35 ][ 113 ],
   alphaCSR[ 35 ][ 114 ],
   alphaCSR[ 35 ][ 115 ],
   alphaCSR[ 35 ][ 116 ],
   alphaCSR[ 35 ][ 117 ],
   alphaCSR[ 35 ][ 118 ],
   alphaCSR[ 35 ][ 119 ],
   alphaCSR[ 35 ][ 120 ],
   alphaCSR[ 35 ][ 121 ],
   alphaCSR[ 35 ][ 122 ],
   alphaCSR[ 35 ][ 123 ],
   alphaCSR[ 35 ][ 124 ],
   alphaCSR[ 35 ][ 125 ],
   alphaCSR[ 35 ][ 126 ],
   alphaCSR[ 35 ][ 127 ],
   alphaCSR[ 35 ][ 128 ],
   alphaCSR[ 35 ][ 129 ],
   alphaCSR[ 35 ][ 130 ],
   alphaCSR[ 35 ][ 131 ],
   alphaCSR[ 35 ][ 132 ],
   alphaCSR[ 35 ][ 133 ],
   alphaCSR[ 35 ][ 134 ],
   alphaCSR[ 35 ][ 135 ],
   alphaCSR[ 35 ][ 136 ],
   alphaCSR[ 35 ][ 137 ],
   alphaCSR[ 35 ][ 138 ],
   alphaCSR[ 35 ][ 139 ],
   alphaCSR[ 35 ][ 140 ],
   alphaCSR[ 35 ][ 141 ],
   alphaCSR[ 35 ][ 142 ],
   alphaCSR[ 35 ][ 143 ],
   alphaCSR[ 35 ][ 144 ],
   alphaCSR[ 35 ][ 145 ],
   alphaCSR[ 35 ][ 146 ],
   alphaCSR[ 35 ][ 147 ],
   alphaCSR[ 35 ][ 148 ],
   alphaCSR[ 35 ][ 149 ],
   alphaCSR[ 35 ][ 150 ],
   alphaCSR[ 35 ][ 151 ],
   alphaCSR[ 35 ][ 152 ],
   alphaCSR[ 35 ][ 153 ],
   alphaCSR[ 35 ][ 154 ],
   alphaCSR[ 35 ][ 155 ],
   alphaCSR[ 35 ][ 156 ],
   alphaCSR[ 35 ][ 157 ],
   alphaCSR[ 35 ][ 158 ],
   alphaCSR[ 35 ][ 159 ],
   alphaCSR[ 35 ][ 160 ],
   alphaCSR[ 35 ][ 161 ],
   alphaCSR[ 35 ][ 162 ],
   alphaCSR[ 35 ][ 163 ],
   alphaCSR[ 35 ][ 164 ],
   alphaCSR[ 35 ][ 165 ],
   alphaCSR[ 35 ][ 166 ],
   alphaCSR[ 35 ][ 167 ],
   alphaCSR[ 35 ][ 168 ],
   alphaCSR[ 35 ][ 169 ],
   alphaCSR[ 35 ][ 170 ],
   alphaCSR[ 35 ][ 171 ],
   alphaCSR[ 35 ][ 172 ],
   alphaCSR[ 35 ][ 173 ],
   alphaCSR[ 35 ][ 174 ],
   alphaCSR[ 35 ][ 175 ],
   alphaCSR[ 35 ][ 176 ],
   alphaCSR[ 35 ][ 177 ],
   alphaCSR[ 35 ][ 178 ],
   alphaCSR[ 35 ][ 179 ],
   alphaCSR[ 35 ][ 180 ],
   alphaCSR[ 35 ][ 181 ],
   alphaCSR[ 35 ][ 182 ],
   alphaCSR[ 35 ][ 183 ],
   alphaCSR[ 35 ][ 184 ],
   alphaCSR[ 35 ][ 185 ],
   alphaCSR[ 35 ][ 186 ],
   alphaCSR[ 35 ][ 187 ],
   alphaCSR[ 35 ][ 188 ],
   alphaCSR[ 35 ][ 189 ],
   alphaCSR[ 35 ][ 190 ],
   alphaCSR[ 35 ][ 191 ],
   alphaCSR[ 35 ][ 192 ],
   alphaCSR[ 35 ][ 193 ],
   alphaCSR[ 35 ][ 194 ],
   alphaCSR[ 35 ][ 195 ],
   alphaCSR[ 35 ][ 196 ],
   alphaCSR[ 35 ][ 197 ],
   alphaCSR[ 35 ][ 198 ],
   alphaCSR[ 35 ][ 199 ],
   alphaCSR[ 35 ][ 200 ],
   alphaCSR[ 35 ][ 201 ],
   alphaCSR[ 35 ][ 202 ],
   alphaCSR[ 35 ][ 203 ],
   alphaCSR[ 35 ][ 204 ],
   alphaCSR[ 35 ][ 205 ],
   alphaCSR[ 35 ][ 206 ],
   alphaCSR[ 35 ][ 207 ],
   alphaCSR[ 35 ][ 208 ],
   alphaCSR[ 35 ][ 209 ],
   alphaCSR[ 35 ][ 210 ],
   alphaCSR[ 35 ][ 211 ],
   alphaCSR[ 35 ][ 212 ],
   alphaCSR[ 35 ][ 213 ],
   alphaCSR[ 35 ][ 214 ],
   alphaCSR[ 35 ][ 215 ],
   alphaCSR[ 35 ][ 216 ],
   alphaCSR[ 35 ][ 217 ],
   alphaCSR[ 35 ][ 218 ],
   alphaCSR[ 35 ][ 219 ],
   alphaCSR[ 35 ][ 220 ],
   alphaCSR[ 35 ][ 221 ],
   alphaCSR[ 35 ][ 222 ],
   alphaCSR[ 35 ][ 223 ],
   alphaCSR[ 35 ][ 224 ],
   alphaCSR[ 35 ][ 225 ],
   alphaCSR[ 35 ][ 226 ],
   alphaCSR[ 35 ][ 227 ],
   alphaCSR[ 35 ][ 228 ],
   alphaCSR[ 35 ][ 229 ],
   alphaCSR[ 35 ][ 230 ],
   alphaCSR[ 35 ][ 231 ],
   alphaCSR[ 35 ][ 232 ],
   alphaCSR[ 35 ][ 233 ],
   alphaCSR[ 35 ][ 234 ],
   alphaCSR[ 35 ][ 235 ],
   alphaCSR[ 35 ][ 236 ],
   alphaCSR[ 35 ][ 237 ],
   alphaCSR[ 35 ][ 238 ],
   alphaCSR[ 35 ][ 239 ],
   alphaCSR[ 35 ][ 240 ],
   alphaCSR[ 35 ][ 241 ],
   alphaCSR[ 35 ][ 242 ],
   alphaCSR[ 35 ][ 243 ],
   alphaCSR[ 35 ][ 244 ],
   alphaCSR[ 35 ][ 245 ],
   alphaCSR[ 35 ][ 246 ],
   alphaCSR[ 35 ][ 247 ],
   alphaCSR[ 35 ][ 248 ],
   alphaCSR[ 35 ][ 249 ],
   alphaCSR[ 35 ][ 250 ],
   alphaCSR[ 35 ][ 251 ],
   alphaCSR[ 35 ][ 252 ],
   alphaCSR[ 35 ][ 253 ],
   alphaCSR[ 35 ][ 254 ],
   alphaCSR[ 35 ][ 255 ],
   alphaCSR[ 35 ][ 256 ],
   alphaCSR[ 35 ][ 257 ],
   alphaCSR[ 35 ][ 258 ],
   alphaCSR[ 35 ][ 259 ],
   alphaCSR[ 35 ][ 260 ],
   alphaCSR[ 35 ][ 261 ],
   alphaCSR[ 35 ][ 262 ],
   alphaCSR[ 35 ][ 263 ],
   alphaCSR[ 35 ][ 264 ],
   alphaCSR[ 35 ][ 265 ],
   alphaCSR[ 35 ][ 266 ],
   alphaCSR[ 35 ][ 267 ],
   alphaCSR[ 35 ][ 268 ],
   alphaCSR[ 35 ][ 269 ],
   alphaCSR[ 35 ][ 270 ],
   alphaCSR[ 35 ][ 271 ],
   alphaCSR[ 35 ][ 272 ],
   alphaCSR[ 35 ][ 273 ],
   alphaCSR[ 35 ][ 274 ],
   alphaCSR[ 35 ][ 275 ],
   alphaCSR[ 35 ][ 276 ],
   alphaCSR[ 35 ][ 277 ],
   alphaCSR[ 35 ][ 278 ],
   alphaCSR[ 35 ][ 279 ],
   alphaCSR[ 35 ][ 280 ],
   alphaCSR[ 35 ][ 281 ],
   alphaCSR[ 35 ][ 282 ],
   alphaCSR[ 35 ][ 283 ],
   alphaCSR[ 35 ][ 284 ],
   alphaCSR[ 35 ][ 285 ],
   alphaCSR[ 35 ][ 286 ],
   alphaCSR[ 35 ][ 287 ],
   alphaCSR[ 35 ][ 288 ],
   alphaCSR[ 35 ][ 289 ],
   alphaCSR[ 35 ][ 290 ],
   alphaCSR[ 35 ][ 291 ],
   alphaCSR[ 35 ][ 292 ],
   alphaCSR[ 35 ][ 293 ],
   alphaCSR[ 35 ][ 294 ],
   alphaCSR[ 35 ][ 295 ],
   alphaCSR[ 35 ][ 296 ],
   alphaCSR[ 35 ][ 297 ],
   alphaCSR[ 35 ][ 298 ],
   alphaCSR[ 35 ][ 299 ],
   alphaCSR[ 35 ][ 300 ],
   alphaCSR[ 35 ][ 301 ],
   alphaCSR[ 35 ][ 302 ],
   alphaCSR[ 35 ][ 303 ],
   alphaCSR[ 35 ][ 304 ],
   alphaCSR[ 35 ][ 305 ],
   alphaCSR[ 35 ][ 306 ],
   alphaCSR[ 35 ][ 307 ],
   alphaCSR[ 35 ][ 308 ],
   alphaCSR[ 35 ][ 309 ],
   alphaCSR[ 35 ][ 310 ],
   alphaCSR[ 35 ][ 311 ],
   alphaCSR[ 35 ][ 312 ],
   alphaCSR[ 35 ][ 313 ],
   alphaCSR[ 35 ][ 314 ],
   alphaCSR[ 35 ][ 315 ],
   alphaCSR[ 35 ][ 316 ],
   alphaCSR[ 35 ][ 317 ],
   alphaCSR[ 35 ][ 318 ],
   alphaCSR[ 35 ][ 319 ],
   alphaCSR[ 35 ][ 320 ],
   alphaCSR[ 35 ][ 321 ],
   alphaCSR[ 35 ][ 322 ],
   alphaCSR[ 35 ][ 323 ],
   alphaCSR[ 35 ][ 324 ],
   alphaCSR[ 35 ][ 325 ],
   alphaCSR[ 35 ][ 326 ],
   alphaCSR[ 35 ][ 327 ],
   alphaCSR[ 35 ][ 328 ],
   alphaCSR[ 35 ][ 329 ],
   alphaCSR[ 35 ][ 330 ],
   alphaCSR[ 35 ][ 331 ],
   alphaCSR[ 35 ][ 332 ],
   alphaCSR[ 35 ][ 333 ],
   alphaCSR[ 35 ][ 334 ],
   alphaCSR[ 35 ][ 335 ],
   alphaCSR[ 35 ][ 336 ],
   alphaCSR[ 35 ][ 337 ],
   alphaCSR[ 35 ][ 338 ],
   alphaCSR[ 35 ][ 339 ],
   alphaCSR[ 35 ][ 340 ],
   alphaCSR[ 35 ][ 341 ],
   alphaCSR[ 35 ][ 342 ],
   alphaCSR[ 35 ][ 343 ],
   alphaCSR[ 35 ][ 344 ],
   alphaCSR[ 35 ][ 345 ],
   alphaCSR[ 35 ][ 346 ],
   alphaCSR[ 35 ][ 347 ],
   alphaCSR[ 35 ][ 348 ],
   alphaCSR[ 35 ][ 349 ],
   alphaCSR[ 35 ][ 350 ],
   alphaCSR[ 35 ][ 351 ],
   alphaCSR[ 35 ][ 352 ],
   alphaCSR[ 35 ][ 353 ],
   alphaCSR[ 35 ][ 354 ],
   alphaCSR[ 35 ][ 355 ],
   alphaCSR[ 35 ][ 356 ],
   alphaCSR[ 35 ][ 357 ],
   alphaCSR[ 35 ][ 358 ],
   alphaCSR[ 35 ][ 359 ],
   alphaCSR[ 35 ][ 360 ],
   alphaCSR[ 35 ][ 361 ],
   alphaCSR[ 35 ][ 362 ],
   alphaCSR[ 35 ][ 363 ],
   alphaCSR[ 35 ][ 364 ],
   alphaCSR[ 35 ][ 365 ],
   alphaCSR[ 35 ][ 366 ],
   alphaCSR[ 35 ][ 367 ],
   alphaCSR[ 35 ][ 368 ],
   alphaCSR[ 35 ][ 369 ],
   alphaCSR[ 35 ][ 370 ],
   alphaCSR[ 35 ][ 371 ],
   alphaCSR[ 35 ][ 372 ],
   alphaCSR[ 35 ][ 373 ],
   alphaCSR[ 35 ][ 374 ],
   alphaCSR[ 35 ][ 375 ],
   alphaCSR[ 35 ][ 376 ],
   alphaCSR[ 35 ][ 377 ],
   alphaCSR[ 35 ][ 378 ],
   alphaCSR[ 35 ][ 379 ],
   alphaCSR[ 35 ][ 380 ],
   alphaCSR[ 35 ][ 381 ],
   alphaCSR[ 35 ][ 382 ],
   alphaCSR[ 35 ][ 383 ],
   alphaCSR[ 36 ][ 0 ],
   alphaCSR[ 36 ][ 1 ],
   alphaCSR[ 36 ][ 2 ],
   alphaCSR[ 36 ][ 3 ],
   alphaCSR[ 36 ][ 4 ],
   alphaCSR[ 36 ][ 5 ],
   alphaCSR[ 36 ][ 6 ],
   alphaCSR[ 36 ][ 7 ],
   alphaCSR[ 36 ][ 8 ],
   alphaCSR[ 36 ][ 9 ],
   alphaCSR[ 36 ][ 10 ],
   alphaCSR[ 36 ][ 11 ],
   alphaCSR[ 36 ][ 12 ],
   alphaCSR[ 36 ][ 13 ],
   alphaCSR[ 36 ][ 14 ],
   alphaCSR[ 36 ][ 15 ],
   alphaCSR[ 36 ][ 16 ],
   alphaCSR[ 36 ][ 17 ],
   alphaCSR[ 36 ][ 18 ],
   alphaCSR[ 36 ][ 19 ],
   alphaCSR[ 36 ][ 20 ],
   alphaCSR[ 36 ][ 21 ],
   alphaCSR[ 36 ][ 22 ],
   alphaCSR[ 36 ][ 23 ],
   alphaCSR[ 36 ][ 24 ],
   alphaCSR[ 36 ][ 25 ],
   alphaCSR[ 36 ][ 26 ],
   alphaCSR[ 36 ][ 27 ],
   alphaCSR[ 36 ][ 28 ],
   alphaCSR[ 36 ][ 29 ],
   alphaCSR[ 36 ][ 30 ],
   alphaCSR[ 36 ][ 31 ],
   alphaCSR[ 36 ][ 32 ],
   alphaCSR[ 36 ][ 33 ],
   alphaCSR[ 36 ][ 34 ],
   alphaCSR[ 36 ][ 35 ],
   alphaCSR[ 36 ][ 36 ],
   alphaCSR[ 36 ][ 37 ],
   alphaCSR[ 36 ][ 38 ],
   alphaCSR[ 36 ][ 39 ],
   alphaCSR[ 36 ][ 40 ],
   alphaCSR[ 36 ][ 41 ],
   alphaCSR[ 36 ][ 42 ],
   alphaCSR[ 36 ][ 43 ],
   alphaCSR[ 36 ][ 44 ],
   alphaCSR[ 36 ][ 45 ],
   alphaCSR[ 36 ][ 46 ],
   alphaCSR[ 36 ][ 47 ],
   alphaCSR[ 36 ][ 48 ],
   alphaCSR[ 36 ][ 49 ],
   alphaCSR[ 36 ][ 50 ],
   alphaCSR[ 36 ][ 51 ],
   alphaCSR[ 36 ][ 52 ],
   alphaCSR[ 36 ][ 53 ],
   alphaCSR[ 36 ][ 54 ],
   alphaCSR[ 36 ][ 55 ],
   alphaCSR[ 36 ][ 56 ],
   alphaCSR[ 36 ][ 57 ],
   alphaCSR[ 36 ][ 58 ],
   alphaCSR[ 36 ][ 59 ],
   alphaCSR[ 36 ][ 60 ],
   alphaCSR[ 36 ][ 61 ],
   alphaCSR[ 36 ][ 62 ],
   alphaCSR[ 36 ][ 63 ],
   alphaCSR[ 36 ][ 64 ],
   alphaCSR[ 36 ][ 65 ],
   alphaCSR[ 36 ][ 66 ],
   alphaCSR[ 36 ][ 67 ],
   alphaCSR[ 36 ][ 68 ],
   alphaCSR[ 36 ][ 69 ],
   alphaCSR[ 36 ][ 70 ],
   alphaCSR[ 36 ][ 71 ],
   alphaCSR[ 36 ][ 72 ],
   alphaCSR[ 36 ][ 73 ],
   alphaCSR[ 36 ][ 74 ],
   alphaCSR[ 36 ][ 75 ],
   alphaCSR[ 36 ][ 76 ],
   alphaCSR[ 36 ][ 77 ],
   alphaCSR[ 36 ][ 78 ],
   alphaCSR[ 36 ][ 79 ],
   alphaCSR[ 36 ][ 80 ],
   alphaCSR[ 36 ][ 81 ],
   alphaCSR[ 36 ][ 82 ],
   alphaCSR[ 36 ][ 83 ],
   alphaCSR[ 36 ][ 84 ],
   alphaCSR[ 36 ][ 85 ],
   alphaCSR[ 36 ][ 86 ],
   alphaCSR[ 36 ][ 87 ],
   alphaCSR[ 36 ][ 88 ],
   alphaCSR[ 36 ][ 89 ],
   alphaCSR[ 36 ][ 90 ],
   alphaCSR[ 36 ][ 91 ],
   alphaCSR[ 36 ][ 92 ],
   alphaCSR[ 36 ][ 93 ],
   alphaCSR[ 36 ][ 94 ],
   alphaCSR[ 36 ][ 95 ],
   alphaCSR[ 36 ][ 96 ],
   alphaCSR[ 36 ][ 97 ],
   alphaCSR[ 36 ][ 98 ],
   alphaCSR[ 36 ][ 99 ],
   alphaCSR[ 36 ][ 100 ],
   alphaCSR[ 36 ][ 101 ],
   alphaCSR[ 36 ][ 102 ],
   alphaCSR[ 36 ][ 103 ],
   alphaCSR[ 36 ][ 104 ],
   alphaCSR[ 36 ][ 105 ],
   alphaCSR[ 36 ][ 106 ],
   alphaCSR[ 36 ][ 107 ],
   alphaCSR[ 36 ][ 108 ],
   alphaCSR[ 36 ][ 109 ],
   alphaCSR[ 36 ][ 110 ],
   alphaCSR[ 36 ][ 111 ],
   alphaCSR[ 36 ][ 112 ],
   alphaCSR[ 36 ][ 113 ],
   alphaCSR[ 36 ][ 114 ],
   alphaCSR[ 36 ][ 115 ],
   alphaCSR[ 36 ][ 116 ],
   alphaCSR[ 36 ][ 117 ],
   alphaCSR[ 36 ][ 118 ],
   alphaCSR[ 36 ][ 119 ],
   alphaCSR[ 36 ][ 120 ],
   alphaCSR[ 36 ][ 121 ],
   alphaCSR[ 36 ][ 122 ],
   alphaCSR[ 36 ][ 123 ],
   alphaCSR[ 36 ][ 124 ],
   alphaCSR[ 36 ][ 125 ],
   alphaCSR[ 36 ][ 126 ],
   alphaCSR[ 36 ][ 127 ],
   alphaCSR[ 36 ][ 128 ],
   alphaCSR[ 36 ][ 129 ],
   alphaCSR[ 36 ][ 130 ],
   alphaCSR[ 36 ][ 131 ],
   alphaCSR[ 36 ][ 132 ],
   alphaCSR[ 36 ][ 133 ],
   alphaCSR[ 36 ][ 134 ],
   alphaCSR[ 36 ][ 135 ],
   alphaCSR[ 36 ][ 136 ],
   alphaCSR[ 36 ][ 137 ],
   alphaCSR[ 36 ][ 138 ],
   alphaCSR[ 36 ][ 139 ],
   alphaCSR[ 36 ][ 140 ],
   alphaCSR[ 36 ][ 141 ],
   alphaCSR[ 36 ][ 142 ],
   alphaCSR[ 36 ][ 143 ],
   alphaCSR[ 36 ][ 144 ],
   alphaCSR[ 36 ][ 145 ],
   alphaCSR[ 36 ][ 146 ],
   alphaCSR[ 36 ][ 147 ],
   alphaCSR[ 36 ][ 148 ],
   alphaCSR[ 36 ][ 149 ],
   alphaCSR[ 36 ][ 150 ],
   alphaCSR[ 36 ][ 151 ],
   alphaCSR[ 36 ][ 152 ],
   alphaCSR[ 36 ][ 153 ],
   alphaCSR[ 36 ][ 154 ],
   alphaCSR[ 36 ][ 155 ],
   alphaCSR[ 36 ][ 156 ],
   alphaCSR[ 36 ][ 157 ],
   alphaCSR[ 36 ][ 158 ],
   alphaCSR[ 36 ][ 159 ],
   alphaCSR[ 36 ][ 160 ],
   alphaCSR[ 36 ][ 161 ],
   alphaCSR[ 36 ][ 162 ],
   alphaCSR[ 36 ][ 163 ],
   alphaCSR[ 36 ][ 164 ],
   alphaCSR[ 36 ][ 165 ],
   alphaCSR[ 36 ][ 166 ],
   alphaCSR[ 36 ][ 167 ],
   alphaCSR[ 36 ][ 168 ],
   alphaCSR[ 36 ][ 169 ],
   alphaCSR[ 36 ][ 170 ],
   alphaCSR[ 36 ][ 171 ],
   alphaCSR[ 36 ][ 172 ],
   alphaCSR[ 36 ][ 173 ],
   alphaCSR[ 36 ][ 174 ],
   alphaCSR[ 36 ][ 175 ],
   alphaCSR[ 36 ][ 176 ],
   alphaCSR[ 36 ][ 177 ],
   alphaCSR[ 36 ][ 178 ],
   alphaCSR[ 36 ][ 179 ],
   alphaCSR[ 36 ][ 180 ],
   alphaCSR[ 36 ][ 181 ],
   alphaCSR[ 36 ][ 182 ],
   alphaCSR[ 36 ][ 183 ],
   alphaCSR[ 36 ][ 184 ],
   alphaCSR[ 36 ][ 185 ],
   alphaCSR[ 36 ][ 186 ],
   alphaCSR[ 36 ][ 187 ],
   alphaCSR[ 36 ][ 188 ],
   alphaCSR[ 36 ][ 189 ],
   alphaCSR[ 36 ][ 190 ],
   alphaCSR[ 36 ][ 191 ],
   alphaCSR[ 36 ][ 192 ],
   alphaCSR[ 36 ][ 193 ],
   alphaCSR[ 36 ][ 194 ],
   alphaCSR[ 36 ][ 195 ],
   alphaCSR[ 36 ][ 196 ],
   alphaCSR[ 36 ][ 197 ],
   alphaCSR[ 36 ][ 198 ],
   alphaCSR[ 36 ][ 199 ],
   alphaCSR[ 36 ][ 200 ],
   alphaCSR[ 36 ][ 201 ],
   alphaCSR[ 36 ][ 202 ],
   alphaCSR[ 36 ][ 203 ],
   alphaCSR[ 36 ][ 204 ],
   alphaCSR[ 36 ][ 205 ],
   alphaCSR[ 36 ][ 206 ],
   alphaCSR[ 36 ][ 207 ],
   alphaCSR[ 36 ][ 208 ],
   alphaCSR[ 36 ][ 209 ],
   alphaCSR[ 36 ][ 210 ],
   alphaCSR[ 36 ][ 211 ],
   alphaCSR[ 36 ][ 212 ],
   alphaCSR[ 36 ][ 213 ],
   alphaCSR[ 36 ][ 214 ],
   alphaCSR[ 36 ][ 215 ],
   alphaCSR[ 36 ][ 216 ],
   alphaCSR[ 36 ][ 217 ],
   alphaCSR[ 36 ][ 218 ],
   alphaCSR[ 36 ][ 219 ],
   alphaCSR[ 36 ][ 220 ],
   alphaCSR[ 36 ][ 221 ],
   alphaCSR[ 36 ][ 222 ],
   alphaCSR[ 36 ][ 223 ],
   alphaCSR[ 36 ][ 224 ],
   alphaCSR[ 36 ][ 225 ],
   alphaCSR[ 36 ][ 226 ],
   alphaCSR[ 36 ][ 227 ],
   alphaCSR[ 36 ][ 228 ],
   alphaCSR[ 36 ][ 229 ],
   alphaCSR[ 36 ][ 230 ],
   alphaCSR[ 36 ][ 231 ],
   alphaCSR[ 36 ][ 232 ],
   alphaCSR[ 36 ][ 233 ],
   alphaCSR[ 36 ][ 234 ],
   alphaCSR[ 36 ][ 235 ],
   alphaCSR[ 36 ][ 236 ],
   alphaCSR[ 36 ][ 237 ],
   alphaCSR[ 36 ][ 238 ],
   alphaCSR[ 36 ][ 239 ],
   alphaCSR[ 36 ][ 240 ],
   alphaCSR[ 36 ][ 241 ],
   alphaCSR[ 36 ][ 242 ],
   alphaCSR[ 36 ][ 243 ],
   alphaCSR[ 36 ][ 244 ],
   alphaCSR[ 36 ][ 245 ],
   alphaCSR[ 36 ][ 246 ],
   alphaCSR[ 36 ][ 247 ],
   alphaCSR[ 36 ][ 248 ],
   alphaCSR[ 36 ][ 249 ],
   alphaCSR[ 36 ][ 250 ],
   alphaCSR[ 36 ][ 251 ],
   alphaCSR[ 36 ][ 252 ],
   alphaCSR[ 36 ][ 253 ],
   alphaCSR[ 36 ][ 254 ],
   alphaCSR[ 36 ][ 255 ],
   alphaCSR[ 36 ][ 256 ],
   alphaCSR[ 36 ][ 257 ],
   alphaCSR[ 36 ][ 258 ],
   alphaCSR[ 36 ][ 259 ],
   alphaCSR[ 36 ][ 260 ],
   alphaCSR[ 36 ][ 261 ],
   alphaCSR[ 36 ][ 262 ],
   alphaCSR[ 36 ][ 263 ],
   alphaCSR[ 36 ][ 264 ],
   alphaCSR[ 36 ][ 265 ],
   alphaCSR[ 36 ][ 266 ],
   alphaCSR[ 36 ][ 267 ],
   alphaCSR[ 36 ][ 268 ],
   alphaCSR[ 36 ][ 269 ],
   alphaCSR[ 36 ][ 270 ],
   alphaCSR[ 36 ][ 271 ],
   alphaCSR[ 36 ][ 272 ],
   alphaCSR[ 36 ][ 273 ],
   alphaCSR[ 36 ][ 274 ],
   alphaCSR[ 36 ][ 275 ],
   alphaCSR[ 36 ][ 276 ],
   alphaCSR[ 36 ][ 277 ],
   alphaCSR[ 36 ][ 278 ],
   alphaCSR[ 36 ][ 279 ],
   alphaCSR[ 36 ][ 280 ],
   alphaCSR[ 36 ][ 281 ],
   alphaCSR[ 36 ][ 282 ],
   alphaCSR[ 36 ][ 283 ],
   alphaCSR[ 36 ][ 284 ],
   alphaCSR[ 36 ][ 285 ],
   alphaCSR[ 36 ][ 286 ],
   alphaCSR[ 36 ][ 287 ],
   alphaCSR[ 36 ][ 288 ],
   alphaCSR[ 36 ][ 289 ],
   alphaCSR[ 36 ][ 290 ],
   alphaCSR[ 36 ][ 291 ],
   alphaCSR[ 36 ][ 292 ],
   alphaCSR[ 36 ][ 293 ],
   alphaCSR[ 36 ][ 294 ],
   alphaCSR[ 36 ][ 295 ],
   alphaCSR[ 36 ][ 296 ],
   alphaCSR[ 36 ][ 297 ],
   alphaCSR[ 36 ][ 298 ],
   alphaCSR[ 36 ][ 299 ],
   alphaCSR[ 36 ][ 300 ],
   alphaCSR[ 36 ][ 301 ],
   alphaCSR[ 36 ][ 302 ],
   alphaCSR[ 36 ][ 303 ],
   alphaCSR[ 36 ][ 304 ],
   alphaCSR[ 36 ][ 305 ],
   alphaCSR[ 36 ][ 306 ],
   alphaCSR[ 36 ][ 307 ],
   alphaCSR[ 36 ][ 308 ],
   alphaCSR[ 36 ][ 309 ],
   alphaCSR[ 36 ][ 310 ],
   alphaCSR[ 36 ][ 311 ],
   alphaCSR[ 36 ][ 312 ],
   alphaCSR[ 36 ][ 313 ],
   alphaCSR[ 36 ][ 314 ],
   alphaCSR[ 36 ][ 315 ],
   alphaCSR[ 36 ][ 316 ],
   alphaCSR[ 36 ][ 317 ],
   alphaCSR[ 36 ][ 318 ],
   alphaCSR[ 36 ][ 319 ],
   alphaCSR[ 36 ][ 320 ],
   alphaCSR[ 36 ][ 321 ],
   alphaCSR[ 36 ][ 322 ],
   alphaCSR[ 36 ][ 323 ],
   alphaCSR[ 36 ][ 324 ],
   alphaCSR[ 36 ][ 325 ],
   alphaCSR[ 36 ][ 326 ],
   alphaCSR[ 36 ][ 327 ],
   alphaCSR[ 36 ][ 328 ],
   alphaCSR[ 36 ][ 329 ],
   alphaCSR[ 36 ][ 330 ],
   alphaCSR[ 36 ][ 331 ],
   alphaCSR[ 36 ][ 332 ],
   alphaCSR[ 36 ][ 333 ],
   alphaCSR[ 36 ][ 334 ],
   alphaCSR[ 36 ][ 335 ],
   alphaCSR[ 36 ][ 336 ],
   alphaCSR[ 36 ][ 337 ],
   alphaCSR[ 36 ][ 338 ],
   alphaCSR[ 36 ][ 339 ],
   alphaCSR[ 36 ][ 340 ],
   alphaCSR[ 36 ][ 341 ],
   alphaCSR[ 36 ][ 342 ],
   alphaCSR[ 36 ][ 343 ],
   alphaCSR[ 36 ][ 344 ],
   alphaCSR[ 36 ][ 345 ],
   alphaCSR[ 36 ][ 346 ],
   alphaCSR[ 36 ][ 347 ],
   alphaCSR[ 36 ][ 348 ],
   alphaCSR[ 36 ][ 349 ],
   alphaCSR[ 36 ][ 350 ],
   alphaCSR[ 36 ][ 351 ],
   alphaCSR[ 36 ][ 352 ],
   alphaCSR[ 36 ][ 353 ],
   alphaCSR[ 36 ][ 354 ],
   alphaCSR[ 36 ][ 355 ],
   alphaCSR[ 36 ][ 356 ],
   alphaCSR[ 36 ][ 357 ],
   alphaCSR[ 36 ][ 358 ],
   alphaCSR[ 36 ][ 359 ],
   alphaCSR[ 36 ][ 360 ],
   alphaCSR[ 36 ][ 361 ],
   alphaCSR[ 36 ][ 362 ],
   alphaCSR[ 36 ][ 363 ],
   alphaCSR[ 36 ][ 364 ],
   alphaCSR[ 36 ][ 365 ],
   alphaCSR[ 36 ][ 366 ],
   alphaCSR[ 36 ][ 367 ],
   alphaCSR[ 36 ][ 368 ],
   alphaCSR[ 36 ][ 369 ],
   alphaCSR[ 36 ][ 370 ],
   alphaCSR[ 36 ][ 371 ],
   alphaCSR[ 36 ][ 372 ],
   alphaCSR[ 36 ][ 373 ],
   alphaCSR[ 36 ][ 374 ],
   alphaCSR[ 36 ][ 375 ],
   alphaCSR[ 36 ][ 376 ],
   alphaCSR[ 36 ][ 377 ],
   alphaCSR[ 36 ][ 378 ],
   alphaCSR[ 36 ][ 379 ],
   alphaCSR[ 36 ][ 380 ],
   alphaCSR[ 36 ][ 381 ],
   alphaCSR[ 36 ][ 382 ],
   alphaCSR[ 36 ][ 383 ],
   alphaCSR[ 37 ][ 0 ],
   alphaCSR[ 37 ][ 1 ],
   alphaCSR[ 37 ][ 2 ],
   alphaCSR[ 37 ][ 3 ],
   alphaCSR[ 37 ][ 4 ],
   alphaCSR[ 37 ][ 5 ],
   alphaCSR[ 37 ][ 6 ],
   alphaCSR[ 37 ][ 7 ],
   alphaCSR[ 37 ][ 8 ],
   alphaCSR[ 37 ][ 9 ],
   alphaCSR[ 37 ][ 10 ],
   alphaCSR[ 37 ][ 11 ],
   alphaCSR[ 37 ][ 12 ],
   alphaCSR[ 37 ][ 13 ],
   alphaCSR[ 37 ][ 14 ],
   alphaCSR[ 37 ][ 15 ],
   alphaCSR[ 37 ][ 16 ],
   alphaCSR[ 37 ][ 17 ],
   alphaCSR[ 37 ][ 18 ],
   alphaCSR[ 37 ][ 19 ],
   alphaCSR[ 37 ][ 20 ],
   alphaCSR[ 37 ][ 21 ],
   alphaCSR[ 37 ][ 22 ],
   alphaCSR[ 37 ][ 23 ],
   alphaCSR[ 37 ][ 24 ],
   alphaCSR[ 37 ][ 25 ],
   alphaCSR[ 37 ][ 26 ],
   alphaCSR[ 37 ][ 27 ],
   alphaCSR[ 37 ][ 28 ],
   alphaCSR[ 37 ][ 29 ],
   alphaCSR[ 37 ][ 30 ],
   alphaCSR[ 37 ][ 31 ],
   alphaCSR[ 37 ][ 32 ],
   alphaCSR[ 37 ][ 33 ],
   alphaCSR[ 37 ][ 34 ],
   alphaCSR[ 37 ][ 35 ],
   alphaCSR[ 37 ][ 36 ],
   alphaCSR[ 37 ][ 37 ],
   alphaCSR[ 37 ][ 38 ],
   alphaCSR[ 37 ][ 39 ],
   alphaCSR[ 37 ][ 40 ],
   alphaCSR[ 37 ][ 41 ],
   alphaCSR[ 37 ][ 42 ],
   alphaCSR[ 37 ][ 43 ],
   alphaCSR[ 37 ][ 44 ],
   alphaCSR[ 37 ][ 45 ],
   alphaCSR[ 37 ][ 46 ],
   alphaCSR[ 37 ][ 47 ],
   alphaCSR[ 37 ][ 48 ],
   alphaCSR[ 37 ][ 49 ],
   alphaCSR[ 37 ][ 50 ],
   alphaCSR[ 37 ][ 51 ],
   alphaCSR[ 37 ][ 52 ],
   alphaCSR[ 37 ][ 53 ],
   alphaCSR[ 37 ][ 54 ],
   alphaCSR[ 37 ][ 55 ],
   alphaCSR[ 37 ][ 56 ],
   alphaCSR[ 37 ][ 57 ],
   alphaCSR[ 37 ][ 58 ],
   alphaCSR[ 37 ][ 59 ],
   alphaCSR[ 37 ][ 60 ],
   alphaCSR[ 37 ][ 61 ],
   alphaCSR[ 37 ][ 62 ],
   alphaCSR[ 37 ][ 63 ],
   alphaCSR[ 37 ][ 64 ],
   alphaCSR[ 37 ][ 65 ],
   alphaCSR[ 37 ][ 66 ],
   alphaCSR[ 37 ][ 67 ],
   alphaCSR[ 37 ][ 68 ],
   alphaCSR[ 37 ][ 69 ],
   alphaCSR[ 37 ][ 70 ],
   alphaCSR[ 37 ][ 71 ],
   alphaCSR[ 37 ][ 72 ],
   alphaCSR[ 37 ][ 73 ],
   alphaCSR[ 37 ][ 74 ],
   alphaCSR[ 37 ][ 75 ],
   alphaCSR[ 37 ][ 76 ],
   alphaCSR[ 37 ][ 77 ],
   alphaCSR[ 37 ][ 78 ],
   alphaCSR[ 37 ][ 79 ],
   alphaCSR[ 37 ][ 80 ],
   alphaCSR[ 37 ][ 81 ],
   alphaCSR[ 37 ][ 82 ],
   alphaCSR[ 37 ][ 83 ],
   alphaCSR[ 37 ][ 84 ],
   alphaCSR[ 37 ][ 85 ],
   alphaCSR[ 37 ][ 86 ],
   alphaCSR[ 37 ][ 87 ],
   alphaCSR[ 37 ][ 88 ],
   alphaCSR[ 37 ][ 89 ],
   alphaCSR[ 37 ][ 90 ],
   alphaCSR[ 37 ][ 91 ],
   alphaCSR[ 37 ][ 92 ],
   alphaCSR[ 37 ][ 93 ],
   alphaCSR[ 37 ][ 94 ],
   alphaCSR[ 37 ][ 95 ],
   alphaCSR[ 37 ][ 96 ],
   alphaCSR[ 37 ][ 97 ],
   alphaCSR[ 37 ][ 98 ],
   alphaCSR[ 37 ][ 99 ],
   alphaCSR[ 37 ][ 100 ],
   alphaCSR[ 37 ][ 101 ],
   alphaCSR[ 37 ][ 102 ],
   alphaCSR[ 37 ][ 103 ],
   alphaCSR[ 37 ][ 104 ],
   alphaCSR[ 37 ][ 105 ],
   alphaCSR[ 37 ][ 106 ],
   alphaCSR[ 37 ][ 107 ],
   alphaCSR[ 37 ][ 108 ],
   alphaCSR[ 37 ][ 109 ],
   alphaCSR[ 37 ][ 110 ],
   alphaCSR[ 37 ][ 111 ],
   alphaCSR[ 37 ][ 112 ],
   alphaCSR[ 37 ][ 113 ],
   alphaCSR[ 37 ][ 114 ],
   alphaCSR[ 37 ][ 115 ],
   alphaCSR[ 37 ][ 116 ],
   alphaCSR[ 37 ][ 117 ],
   alphaCSR[ 37 ][ 118 ],
   alphaCSR[ 37 ][ 119 ],
   alphaCSR[ 37 ][ 120 ],
   alphaCSR[ 37 ][ 121 ],
   alphaCSR[ 37 ][ 122 ],
   alphaCSR[ 37 ][ 123 ],
   alphaCSR[ 37 ][ 124 ],
   alphaCSR[ 37 ][ 125 ],
   alphaCSR[ 37 ][ 126 ],
   alphaCSR[ 37 ][ 127 ],
   alphaCSR[ 37 ][ 128 ],
   alphaCSR[ 37 ][ 129 ],
   alphaCSR[ 37 ][ 130 ],
   alphaCSR[ 37 ][ 131 ],
   alphaCSR[ 37 ][ 132 ],
   alphaCSR[ 37 ][ 133 ],
   alphaCSR[ 37 ][ 134 ],
   alphaCSR[ 37 ][ 135 ],
   alphaCSR[ 37 ][ 136 ],
   alphaCSR[ 37 ][ 137 ],
   alphaCSR[ 37 ][ 138 ],
   alphaCSR[ 37 ][ 139 ],
   alphaCSR[ 37 ][ 140 ],
   alphaCSR[ 37 ][ 141 ],
   alphaCSR[ 37 ][ 142 ],
   alphaCSR[ 37 ][ 143 ],
   alphaCSR[ 37 ][ 144 ],
   alphaCSR[ 37 ][ 145 ],
   alphaCSR[ 37 ][ 146 ],
   alphaCSR[ 37 ][ 147 ],
   alphaCSR[ 37 ][ 148 ],
   alphaCSR[ 37 ][ 149 ],
   alphaCSR[ 37 ][ 150 ],
   alphaCSR[ 37 ][ 151 ],
   alphaCSR[ 37 ][ 152 ],
   alphaCSR[ 37 ][ 153 ],
   alphaCSR[ 37 ][ 154 ],
   alphaCSR[ 37 ][ 155 ],
   alphaCSR[ 37 ][ 156 ],
   alphaCSR[ 37 ][ 157 ],
   alphaCSR[ 37 ][ 158 ],
   alphaCSR[ 37 ][ 159 ],
   alphaCSR[ 37 ][ 160 ],
   alphaCSR[ 37 ][ 161 ],
   alphaCSR[ 37 ][ 162 ],
   alphaCSR[ 37 ][ 163 ],
   alphaCSR[ 37 ][ 164 ],
   alphaCSR[ 37 ][ 165 ],
   alphaCSR[ 37 ][ 166 ],
   alphaCSR[ 37 ][ 167 ],
   alphaCSR[ 37 ][ 168 ],
   alphaCSR[ 37 ][ 169 ],
   alphaCSR[ 37 ][ 170 ],
   alphaCSR[ 37 ][ 171 ],
   alphaCSR[ 37 ][ 172 ],
   alphaCSR[ 37 ][ 173 ],
   alphaCSR[ 37 ][ 174 ],
   alphaCSR[ 37 ][ 175 ],
   alphaCSR[ 37 ][ 176 ],
   alphaCSR[ 37 ][ 177 ],
   alphaCSR[ 37 ][ 178 ],
   alphaCSR[ 37 ][ 179 ],
   alphaCSR[ 37 ][ 180 ],
   alphaCSR[ 37 ][ 181 ],
   alphaCSR[ 37 ][ 182 ],
   alphaCSR[ 37 ][ 183 ],
   alphaCSR[ 37 ][ 184 ],
   alphaCSR[ 37 ][ 185 ],
   alphaCSR[ 37 ][ 186 ],
   alphaCSR[ 37 ][ 187 ],
   alphaCSR[ 37 ][ 188 ],
   alphaCSR[ 37 ][ 189 ],
   alphaCSR[ 37 ][ 190 ],
   alphaCSR[ 37 ][ 191 ],
   alphaCSR[ 37 ][ 192 ],
   alphaCSR[ 37 ][ 193 ],
   alphaCSR[ 37 ][ 194 ],
   alphaCSR[ 37 ][ 195 ],
   alphaCSR[ 37 ][ 196 ],
   alphaCSR[ 37 ][ 197 ],
   alphaCSR[ 37 ][ 198 ],
   alphaCSR[ 37 ][ 199 ],
   alphaCSR[ 37 ][ 200 ],
   alphaCSR[ 37 ][ 201 ],
   alphaCSR[ 37 ][ 202 ],
   alphaCSR[ 37 ][ 203 ],
   alphaCSR[ 37 ][ 204 ],
   alphaCSR[ 37 ][ 205 ],
   alphaCSR[ 37 ][ 206 ],
   alphaCSR[ 37 ][ 207 ],
   alphaCSR[ 37 ][ 208 ],
   alphaCSR[ 37 ][ 209 ],
   alphaCSR[ 37 ][ 210 ],
   alphaCSR[ 37 ][ 211 ],
   alphaCSR[ 37 ][ 212 ],
   alphaCSR[ 37 ][ 213 ],
   alphaCSR[ 37 ][ 214 ],
   alphaCSR[ 37 ][ 215 ],
   alphaCSR[ 37 ][ 216 ],
   alphaCSR[ 37 ][ 217 ],
   alphaCSR[ 37 ][ 218 ],
   alphaCSR[ 37 ][ 219 ],
   alphaCSR[ 37 ][ 220 ],
   alphaCSR[ 37 ][ 221 ],
   alphaCSR[ 37 ][ 222 ],
   alphaCSR[ 37 ][ 223 ],
   alphaCSR[ 37 ][ 224 ],
   alphaCSR[ 37 ][ 225 ],
   alphaCSR[ 37 ][ 226 ],
   alphaCSR[ 37 ][ 227 ],
   alphaCSR[ 37 ][ 228 ],
   alphaCSR[ 37 ][ 229 ],
   alphaCSR[ 37 ][ 230 ],
   alphaCSR[ 37 ][ 231 ],
   alphaCSR[ 37 ][ 232 ],
   alphaCSR[ 37 ][ 233 ],
   alphaCSR[ 37 ][ 234 ],
   alphaCSR[ 37 ][ 235 ],
   alphaCSR[ 37 ][ 236 ],
   alphaCSR[ 37 ][ 237 ],
   alphaCSR[ 37 ][ 238 ],
   alphaCSR[ 37 ][ 239 ],
   alphaCSR[ 37 ][ 240 ],
   alphaCSR[ 37 ][ 241 ],
   alphaCSR[ 37 ][ 242 ],
   alphaCSR[ 37 ][ 243 ],
   alphaCSR[ 37 ][ 244 ],
   alphaCSR[ 37 ][ 245 ],
   alphaCSR[ 37 ][ 246 ],
   alphaCSR[ 37 ][ 247 ],
   alphaCSR[ 37 ][ 248 ],
   alphaCSR[ 37 ][ 249 ],
   alphaCSR[ 37 ][ 250 ],
   alphaCSR[ 37 ][ 251 ],
   alphaCSR[ 37 ][ 252 ],
   alphaCSR[ 37 ][ 253 ],
   alphaCSR[ 37 ][ 254 ],
   alphaCSR[ 37 ][ 255 ],
   alphaCSR[ 37 ][ 256 ],
   alphaCSR[ 37 ][ 257 ],
   alphaCSR[ 37 ][ 258 ],
   alphaCSR[ 37 ][ 259 ],
   alphaCSR[ 37 ][ 260 ],
   alphaCSR[ 37 ][ 261 ],
   alphaCSR[ 37 ][ 262 ],
   alphaCSR[ 37 ][ 263 ],
   alphaCSR[ 37 ][ 264 ],
   alphaCSR[ 37 ][ 265 ],
   alphaCSR[ 37 ][ 266 ],
   alphaCSR[ 37 ][ 267 ],
   alphaCSR[ 37 ][ 268 ],
   alphaCSR[ 37 ][ 269 ],
   alphaCSR[ 37 ][ 270 ],
   alphaCSR[ 37 ][ 271 ],
   alphaCSR[ 37 ][ 272 ],
   alphaCSR[ 37 ][ 273 ],
   alphaCSR[ 37 ][ 274 ],
   alphaCSR[ 37 ][ 275 ],
   alphaCSR[ 37 ][ 276 ],
   alphaCSR[ 37 ][ 277 ],
   alphaCSR[ 37 ][ 278 ],
   alphaCSR[ 37 ][ 279 ],
   alphaCSR[ 37 ][ 280 ],
   alphaCSR[ 37 ][ 281 ],
   alphaCSR[ 37 ][ 282 ],
   alphaCSR[ 37 ][ 283 ],
   alphaCSR[ 37 ][ 284 ],
   alphaCSR[ 37 ][ 285 ],
   alphaCSR[ 37 ][ 286 ],
   alphaCSR[ 37 ][ 287 ],
   alphaCSR[ 37 ][ 288 ],
   alphaCSR[ 37 ][ 289 ],
   alphaCSR[ 37 ][ 290 ],
   alphaCSR[ 37 ][ 291 ],
   alphaCSR[ 37 ][ 292 ],
   alphaCSR[ 37 ][ 293 ],
   alphaCSR[ 37 ][ 294 ],
   alphaCSR[ 37 ][ 295 ],
   alphaCSR[ 37 ][ 296 ],
   alphaCSR[ 37 ][ 297 ],
   alphaCSR[ 37 ][ 298 ],
   alphaCSR[ 37 ][ 299 ],
   alphaCSR[ 37 ][ 300 ],
   alphaCSR[ 37 ][ 301 ],
   alphaCSR[ 37 ][ 302 ],
   alphaCSR[ 37 ][ 303 ],
   alphaCSR[ 37 ][ 304 ],
   alphaCSR[ 37 ][ 305 ],
   alphaCSR[ 37 ][ 306 ],
   alphaCSR[ 37 ][ 307 ],
   alphaCSR[ 37 ][ 308 ],
   alphaCSR[ 37 ][ 309 ],
   alphaCSR[ 37 ][ 310 ],
   alphaCSR[ 37 ][ 311 ],
   alphaCSR[ 37 ][ 312 ],
   alphaCSR[ 37 ][ 313 ],
   alphaCSR[ 37 ][ 314 ],
   alphaCSR[ 37 ][ 315 ],
   alphaCSR[ 37 ][ 316 ],
   alphaCSR[ 37 ][ 317 ],
   alphaCSR[ 37 ][ 318 ],
   alphaCSR[ 37 ][ 319 ],
   alphaCSR[ 37 ][ 320 ],
   alphaCSR[ 37 ][ 321 ],
   alphaCSR[ 37 ][ 322 ],
   alphaCSR[ 37 ][ 323 ],
   alphaCSR[ 37 ][ 324 ],
   alphaCSR[ 37 ][ 325 ],
   alphaCSR[ 37 ][ 326 ],
   alphaCSR[ 37 ][ 327 ],
   alphaCSR[ 37 ][ 328 ],
   alphaCSR[ 37 ][ 329 ],
   alphaCSR[ 37 ][ 330 ],
   alphaCSR[ 37 ][ 331 ],
   alphaCSR[ 37 ][ 332 ],
   alphaCSR[ 37 ][ 333 ],
   alphaCSR[ 37 ][ 334 ],
   alphaCSR[ 37 ][ 335 ],
   alphaCSR[ 37 ][ 336 ],
   alphaCSR[ 37 ][ 337 ],
   alphaCSR[ 37 ][ 338 ],
   alphaCSR[ 37 ][ 339 ],
   alphaCSR[ 37 ][ 340 ],
   alphaCSR[ 37 ][ 341 ],
   alphaCSR[ 37 ][ 342 ],
   alphaCSR[ 37 ][ 343 ],
   alphaCSR[ 37 ][ 344 ],
   alphaCSR[ 37 ][ 345 ],
   alphaCSR[ 37 ][ 346 ],
   alphaCSR[ 37 ][ 347 ],
   alphaCSR[ 37 ][ 348 ],
   alphaCSR[ 37 ][ 349 ],
   alphaCSR[ 37 ][ 350 ],
   alphaCSR[ 37 ][ 351 ],
   alphaCSR[ 37 ][ 352 ],
   alphaCSR[ 37 ][ 353 ],
   alphaCSR[ 37 ][ 354 ],
   alphaCSR[ 37 ][ 355 ],
   alphaCSR[ 37 ][ 356 ],
   alphaCSR[ 37 ][ 357 ],
   alphaCSR[ 37 ][ 358 ],
   alphaCSR[ 37 ][ 359 ],
   alphaCSR[ 37 ][ 360 ],
   alphaCSR[ 37 ][ 361 ],
   alphaCSR[ 37 ][ 362 ],
   alphaCSR[ 37 ][ 363 ],
   alphaCSR[ 37 ][ 364 ],
   alphaCSR[ 37 ][ 365 ],
   alphaCSR[ 37 ][ 366 ],
   alphaCSR[ 37 ][ 367 ],
   alphaCSR[ 37 ][ 368 ],
   alphaCSR[ 37 ][ 369 ],
   alphaCSR[ 37 ][ 370 ],
   alphaCSR[ 37 ][ 371 ],
   alphaCSR[ 37 ][ 372 ],
   alphaCSR[ 37 ][ 373 ],
   alphaCSR[ 37 ][ 374 ],
   alphaCSR[ 37 ][ 375 ],
   alphaCSR[ 37 ][ 376 ],
   alphaCSR[ 37 ][ 377 ],
   alphaCSR[ 37 ][ 378 ],
   alphaCSR[ 37 ][ 379 ],
   alphaCSR[ 37 ][ 380 ],
   alphaCSR[ 37 ][ 381 ],
   alphaCSR[ 37 ][ 382 ],
   alphaCSR[ 37 ][ 383 ],
   alphaCSR[ 38 ][ 0 ],
   alphaCSR[ 38 ][ 1 ],
   alphaCSR[ 38 ][ 2 ],
   alphaCSR[ 38 ][ 3 ],
   alphaCSR[ 38 ][ 4 ],
   alphaCSR[ 38 ][ 5 ],
   alphaCSR[ 38 ][ 6 ],
   alphaCSR[ 38 ][ 7 ],
   alphaCSR[ 38 ][ 8 ],
   alphaCSR[ 38 ][ 9 ],
   alphaCSR[ 38 ][ 10 ],
   alphaCSR[ 38 ][ 11 ],
   alphaCSR[ 38 ][ 12 ],
   alphaCSR[ 38 ][ 13 ],
   alphaCSR[ 38 ][ 14 ],
   alphaCSR[ 38 ][ 15 ],
   alphaCSR[ 38 ][ 16 ],
   alphaCSR[ 38 ][ 17 ],
   alphaCSR[ 38 ][ 18 ],
   alphaCSR[ 38 ][ 19 ],
   alphaCSR[ 38 ][ 20 ],
   alphaCSR[ 38 ][ 21 ],
   alphaCSR[ 38 ][ 22 ],
   alphaCSR[ 38 ][ 23 ],
   alphaCSR[ 38 ][ 24 ],
   alphaCSR[ 38 ][ 25 ],
   alphaCSR[ 38 ][ 26 ],
   alphaCSR[ 38 ][ 27 ],
   alphaCSR[ 38 ][ 28 ],
   alphaCSR[ 38 ][ 29 ],
   alphaCSR[ 38 ][ 30 ],
   alphaCSR[ 38 ][ 31 ],
   alphaCSR[ 38 ][ 32 ],
   alphaCSR[ 38 ][ 33 ],
   alphaCSR[ 38 ][ 34 ],
   alphaCSR[ 38 ][ 35 ],
   alphaCSR[ 38 ][ 36 ],
   alphaCSR[ 38 ][ 37 ],
   alphaCSR[ 38 ][ 38 ],
   alphaCSR[ 38 ][ 39 ],
   alphaCSR[ 38 ][ 40 ],
   alphaCSR[ 38 ][ 41 ],
   alphaCSR[ 38 ][ 42 ],
   alphaCSR[ 38 ][ 43 ],
   alphaCSR[ 38 ][ 44 ],
   alphaCSR[ 38 ][ 45 ],
   alphaCSR[ 38 ][ 46 ],
   alphaCSR[ 38 ][ 47 ],
   alphaCSR[ 38 ][ 48 ],
   alphaCSR[ 38 ][ 49 ],
   alphaCSR[ 38 ][ 50 ],
   alphaCSR[ 38 ][ 51 ],
   alphaCSR[ 38 ][ 52 ],
   alphaCSR[ 38 ][ 53 ],
   alphaCSR[ 38 ][ 54 ],
   alphaCSR[ 38 ][ 55 ],
   alphaCSR[ 38 ][ 56 ],
   alphaCSR[ 38 ][ 57 ],
   alphaCSR[ 38 ][ 58 ],
   alphaCSR[ 38 ][ 59 ],
   alphaCSR[ 38 ][ 60 ],
   alphaCSR[ 38 ][ 61 ],
   alphaCSR[ 38 ][ 62 ],
   alphaCSR[ 38 ][ 63 ],
   alphaCSR[ 38 ][ 64 ],
   alphaCSR[ 38 ][ 65 ],
   alphaCSR[ 38 ][ 66 ],
   alphaCSR[ 38 ][ 67 ],
   alphaCSR[ 38 ][ 68 ],
   alphaCSR[ 38 ][ 69 ],
   alphaCSR[ 38 ][ 70 ],
   alphaCSR[ 38 ][ 71 ],
   alphaCSR[ 38 ][ 72 ],
   alphaCSR[ 38 ][ 73 ],
   alphaCSR[ 38 ][ 74 ],
   alphaCSR[ 38 ][ 75 ],
   alphaCSR[ 38 ][ 76 ],
   alphaCSR[ 38 ][ 77 ],
   alphaCSR[ 38 ][ 78 ],
   alphaCSR[ 38 ][ 79 ],
   alphaCSR[ 38 ][ 80 ],
   alphaCSR[ 38 ][ 81 ],
   alphaCSR[ 38 ][ 82 ],
   alphaCSR[ 38 ][ 83 ],
   alphaCSR[ 38 ][ 84 ],
   alphaCSR[ 38 ][ 85 ],
   alphaCSR[ 38 ][ 86 ],
   alphaCSR[ 38 ][ 87 ],
   alphaCSR[ 38 ][ 88 ],
   alphaCSR[ 38 ][ 89 ],
   alphaCSR[ 38 ][ 90 ],
   alphaCSR[ 38 ][ 91 ],
   alphaCSR[ 38 ][ 92 ],
   alphaCSR[ 38 ][ 93 ],
   alphaCSR[ 38 ][ 94 ],
   alphaCSR[ 38 ][ 95 ],
   alphaCSR[ 38 ][ 96 ],
   alphaCSR[ 38 ][ 97 ],
   alphaCSR[ 38 ][ 98 ],
   alphaCSR[ 38 ][ 99 ],
   alphaCSR[ 38 ][ 100 ],
   alphaCSR[ 38 ][ 101 ],
   alphaCSR[ 38 ][ 102 ],
   alphaCSR[ 38 ][ 103 ],
   alphaCSR[ 38 ][ 104 ],
   alphaCSR[ 38 ][ 105 ],
   alphaCSR[ 38 ][ 106 ],
   alphaCSR[ 38 ][ 107 ],
   alphaCSR[ 38 ][ 108 ],
   alphaCSR[ 38 ][ 109 ],
   alphaCSR[ 38 ][ 110 ],
   alphaCSR[ 38 ][ 111 ],
   alphaCSR[ 38 ][ 112 ],
   alphaCSR[ 38 ][ 113 ],
   alphaCSR[ 38 ][ 114 ],
   alphaCSR[ 38 ][ 115 ],
   alphaCSR[ 38 ][ 116 ],
   alphaCSR[ 38 ][ 117 ],
   alphaCSR[ 38 ][ 118 ],
   alphaCSR[ 38 ][ 119 ],
   alphaCSR[ 38 ][ 120 ],
   alphaCSR[ 38 ][ 121 ],
   alphaCSR[ 38 ][ 122 ],
   alphaCSR[ 38 ][ 123 ],
   alphaCSR[ 38 ][ 124 ],
   alphaCSR[ 38 ][ 125 ],
   alphaCSR[ 38 ][ 126 ],
   alphaCSR[ 38 ][ 127 ],
   alphaCSR[ 38 ][ 128 ],
   alphaCSR[ 38 ][ 129 ],
   alphaCSR[ 38 ][ 130 ],
   alphaCSR[ 38 ][ 131 ],
   alphaCSR[ 38 ][ 132 ],
   alphaCSR[ 38 ][ 133 ],
   alphaCSR[ 38 ][ 134 ],
   alphaCSR[ 38 ][ 135 ],
   alphaCSR[ 38 ][ 136 ],
   alphaCSR[ 38 ][ 137 ],
   alphaCSR[ 38 ][ 138 ],
   alphaCSR[ 38 ][ 139 ],
   alphaCSR[ 38 ][ 140 ],
   alphaCSR[ 38 ][ 141 ],
   alphaCSR[ 38 ][ 142 ],
   alphaCSR[ 38 ][ 143 ],
   alphaCSR[ 38 ][ 144 ],
   alphaCSR[ 38 ][ 145 ],
   alphaCSR[ 38 ][ 146 ],
   alphaCSR[ 38 ][ 147 ],
   alphaCSR[ 38 ][ 148 ],
   alphaCSR[ 38 ][ 149 ],
   alphaCSR[ 38 ][ 150 ],
   alphaCSR[ 38 ][ 151 ],
   alphaCSR[ 38 ][ 152 ],
   alphaCSR[ 38 ][ 153 ],
   alphaCSR[ 38 ][ 154 ],
   alphaCSR[ 38 ][ 155 ],
   alphaCSR[ 38 ][ 156 ],
   alphaCSR[ 38 ][ 157 ],
   alphaCSR[ 38 ][ 158 ],
   alphaCSR[ 38 ][ 159 ],
   alphaCSR[ 38 ][ 160 ],
   alphaCSR[ 38 ][ 161 ],
   alphaCSR[ 38 ][ 162 ],
   alphaCSR[ 38 ][ 163 ],
   alphaCSR[ 38 ][ 164 ],
   alphaCSR[ 38 ][ 165 ],
   alphaCSR[ 38 ][ 166 ],
   alphaCSR[ 38 ][ 167 ],
   alphaCSR[ 38 ][ 168 ],
   alphaCSR[ 38 ][ 169 ],
   alphaCSR[ 38 ][ 170 ],
   alphaCSR[ 38 ][ 171 ],
   alphaCSR[ 38 ][ 172 ],
   alphaCSR[ 38 ][ 173 ],
   alphaCSR[ 38 ][ 174 ],
   alphaCSR[ 38 ][ 175 ],
   alphaCSR[ 38 ][ 176 ],
   alphaCSR[ 38 ][ 177 ],
   alphaCSR[ 38 ][ 178 ],
   alphaCSR[ 38 ][ 179 ],
   alphaCSR[ 38 ][ 180 ],
   alphaCSR[ 38 ][ 181 ],
   alphaCSR[ 38 ][ 182 ],
   alphaCSR[ 38 ][ 183 ],
   alphaCSR[ 38 ][ 184 ],
   alphaCSR[ 38 ][ 185 ],
   alphaCSR[ 38 ][ 186 ],
   alphaCSR[ 38 ][ 187 ],
   alphaCSR[ 38 ][ 188 ],
   alphaCSR[ 38 ][ 189 ],
   alphaCSR[ 38 ][ 190 ],
   alphaCSR[ 38 ][ 191 ],
   alphaCSR[ 38 ][ 192 ],
   alphaCSR[ 38 ][ 193 ],
   alphaCSR[ 38 ][ 194 ],
   alphaCSR[ 38 ][ 195 ],
   alphaCSR[ 38 ][ 196 ],
   alphaCSR[ 38 ][ 197 ],
   alphaCSR[ 38 ][ 198 ],
   alphaCSR[ 38 ][ 199 ],
   alphaCSR[ 38 ][ 200 ],
   alphaCSR[ 38 ][ 201 ],
   alphaCSR[ 38 ][ 202 ],
   alphaCSR[ 38 ][ 203 ],
   alphaCSR[ 38 ][ 204 ],
   alphaCSR[ 38 ][ 205 ],
   alphaCSR[ 38 ][ 206 ],
   alphaCSR[ 38 ][ 207 ],
   alphaCSR[ 38 ][ 208 ],
   alphaCSR[ 38 ][ 209 ],
   alphaCSR[ 38 ][ 210 ],
   alphaCSR[ 38 ][ 211 ],
   alphaCSR[ 38 ][ 212 ],
   alphaCSR[ 38 ][ 213 ],
   alphaCSR[ 38 ][ 214 ],
   alphaCSR[ 38 ][ 215 ],
   alphaCSR[ 38 ][ 216 ],
   alphaCSR[ 38 ][ 217 ],
   alphaCSR[ 38 ][ 218 ],
   alphaCSR[ 38 ][ 219 ],
   alphaCSR[ 38 ][ 220 ],
   alphaCSR[ 38 ][ 221 ],
   alphaCSR[ 38 ][ 222 ],
   alphaCSR[ 38 ][ 223 ],
   alphaCSR[ 38 ][ 224 ],
   alphaCSR[ 38 ][ 225 ],
   alphaCSR[ 38 ][ 226 ],
   alphaCSR[ 38 ][ 227 ],
   alphaCSR[ 38 ][ 228 ],
   alphaCSR[ 38 ][ 229 ],
   alphaCSR[ 38 ][ 230 ],
   alphaCSR[ 38 ][ 231 ],
   alphaCSR[ 38 ][ 232 ],
   alphaCSR[ 38 ][ 233 ],
   alphaCSR[ 38 ][ 234 ],
   alphaCSR[ 38 ][ 235 ],
   alphaCSR[ 38 ][ 236 ],
   alphaCSR[ 38 ][ 237 ],
   alphaCSR[ 38 ][ 238 ],
   alphaCSR[ 38 ][ 239 ],
   alphaCSR[ 38 ][ 240 ],
   alphaCSR[ 38 ][ 241 ],
   alphaCSR[ 38 ][ 242 ],
   alphaCSR[ 38 ][ 243 ],
   alphaCSR[ 38 ][ 244 ],
   alphaCSR[ 38 ][ 245 ],
   alphaCSR[ 38 ][ 246 ],
   alphaCSR[ 38 ][ 247 ],
   alphaCSR[ 38 ][ 248 ],
   alphaCSR[ 38 ][ 249 ],
   alphaCSR[ 38 ][ 250 ],
   alphaCSR[ 38 ][ 251 ],
   alphaCSR[ 38 ][ 252 ],
   alphaCSR[ 38 ][ 253 ],
   alphaCSR[ 38 ][ 254 ],
   alphaCSR[ 38 ][ 255 ],
   alphaCSR[ 38 ][ 256 ],
   alphaCSR[ 38 ][ 257 ],
   alphaCSR[ 38 ][ 258 ],
   alphaCSR[ 38 ][ 259 ],
   alphaCSR[ 38 ][ 260 ],
   alphaCSR[ 38 ][ 261 ],
   alphaCSR[ 38 ][ 262 ],
   alphaCSR[ 38 ][ 263 ],
   alphaCSR[ 38 ][ 264 ],
   alphaCSR[ 38 ][ 265 ],
   alphaCSR[ 38 ][ 266 ],
   alphaCSR[ 38 ][ 267 ],
   alphaCSR[ 38 ][ 268 ],
   alphaCSR[ 38 ][ 269 ],
   alphaCSR[ 38 ][ 270 ],
   alphaCSR[ 38 ][ 271 ],
   alphaCSR[ 38 ][ 272 ],
   alphaCSR[ 38 ][ 273 ],
   alphaCSR[ 38 ][ 274 ],
   alphaCSR[ 38 ][ 275 ],
   alphaCSR[ 38 ][ 276 ],
   alphaCSR[ 38 ][ 277 ],
   alphaCSR[ 38 ][ 278 ],
   alphaCSR[ 38 ][ 279 ],
   alphaCSR[ 38 ][ 280 ],
   alphaCSR[ 38 ][ 281 ],
   alphaCSR[ 38 ][ 282 ],
   alphaCSR[ 38 ][ 283 ],
   alphaCSR[ 38 ][ 284 ],
   alphaCSR[ 38 ][ 285 ],
   alphaCSR[ 38 ][ 286 ],
   alphaCSR[ 38 ][ 287 ],
   alphaCSR[ 38 ][ 288 ],
   alphaCSR[ 38 ][ 289 ],
   alphaCSR[ 38 ][ 290 ],
   alphaCSR[ 38 ][ 291 ],
   alphaCSR[ 38 ][ 292 ],
   alphaCSR[ 38 ][ 293 ],
   alphaCSR[ 38 ][ 294 ],
   alphaCSR[ 38 ][ 295 ],
   alphaCSR[ 38 ][ 296 ],
   alphaCSR[ 38 ][ 297 ],
   alphaCSR[ 38 ][ 298 ],
   alphaCSR[ 38 ][ 299 ],
   alphaCSR[ 38 ][ 300 ],
   alphaCSR[ 38 ][ 301 ],
   alphaCSR[ 38 ][ 302 ],
   alphaCSR[ 38 ][ 303 ],
   alphaCSR[ 38 ][ 304 ],
   alphaCSR[ 38 ][ 305 ],
   alphaCSR[ 38 ][ 306 ],
   alphaCSR[ 38 ][ 307 ],
   alphaCSR[ 38 ][ 308 ],
   alphaCSR[ 38 ][ 309 ],
   alphaCSR[ 38 ][ 310 ],
   alphaCSR[ 38 ][ 311 ],
   alphaCSR[ 38 ][ 312 ],
   alphaCSR[ 38 ][ 313 ],
   alphaCSR[ 38 ][ 314 ],
   alphaCSR[ 38 ][ 315 ],
   alphaCSR[ 38 ][ 316 ],
   alphaCSR[ 38 ][ 317 ],
   alphaCSR[ 38 ][ 318 ],
   alphaCSR[ 38 ][ 319 ],
   alphaCSR[ 38 ][ 320 ],
   alphaCSR[ 38 ][ 321 ],
   alphaCSR[ 38 ][ 322 ],
   alphaCSR[ 38 ][ 323 ],
   alphaCSR[ 38 ][ 324 ],
   alphaCSR[ 38 ][ 325 ],
   alphaCSR[ 38 ][ 326 ],
   alphaCSR[ 38 ][ 327 ],
   alphaCSR[ 38 ][ 328 ],
   alphaCSR[ 38 ][ 329 ],
   alphaCSR[ 38 ][ 330 ],
   alphaCSR[ 38 ][ 331 ],
   alphaCSR[ 38 ][ 332 ],
   alphaCSR[ 38 ][ 333 ],
   alphaCSR[ 38 ][ 334 ],
   alphaCSR[ 38 ][ 335 ],
   alphaCSR[ 38 ][ 336 ],
   alphaCSR[ 38 ][ 337 ],
   alphaCSR[ 38 ][ 338 ],
   alphaCSR[ 38 ][ 339 ],
   alphaCSR[ 38 ][ 340 ],
   alphaCSR[ 38 ][ 341 ],
   alphaCSR[ 38 ][ 342 ],
   alphaCSR[ 38 ][ 343 ],
   alphaCSR[ 38 ][ 344 ],
   alphaCSR[ 38 ][ 345 ],
   alphaCSR[ 38 ][ 346 ],
   alphaCSR[ 38 ][ 347 ],
   alphaCSR[ 38 ][ 348 ],
   alphaCSR[ 38 ][ 349 ],
   alphaCSR[ 38 ][ 350 ],
   alphaCSR[ 38 ][ 351 ],
   alphaCSR[ 38 ][ 352 ],
   alphaCSR[ 38 ][ 353 ],
   alphaCSR[ 38 ][ 354 ],
   alphaCSR[ 38 ][ 355 ],
   alphaCSR[ 38 ][ 356 ],
   alphaCSR[ 38 ][ 357 ],
   alphaCSR[ 38 ][ 358 ],
   alphaCSR[ 38 ][ 359 ],
   alphaCSR[ 38 ][ 360 ],
   alphaCSR[ 38 ][ 361 ],
   alphaCSR[ 38 ][ 362 ],
   alphaCSR[ 38 ][ 363 ],
   alphaCSR[ 38 ][ 364 ],
   alphaCSR[ 38 ][ 365 ],
   alphaCSR[ 38 ][ 366 ],
   alphaCSR[ 38 ][ 367 ],
   alphaCSR[ 38 ][ 368 ],
   alphaCSR[ 38 ][ 369 ],
   alphaCSR[ 38 ][ 370 ],
   alphaCSR[ 38 ][ 371 ],
   alphaCSR[ 38 ][ 372 ],
   alphaCSR[ 38 ][ 373 ],
   alphaCSR[ 38 ][ 374 ],
   alphaCSR[ 38 ][ 375 ],
   alphaCSR[ 38 ][ 376 ],
   alphaCSR[ 38 ][ 377 ],
   alphaCSR[ 38 ][ 378 ],
   alphaCSR[ 38 ][ 379 ],
   alphaCSR[ 38 ][ 380 ],
   alphaCSR[ 38 ][ 381 ],
   alphaCSR[ 38 ][ 382 ],
   alphaCSR[ 38 ][ 383 ],
   alphaCSR[ 39 ][ 0 ],
   alphaCSR[ 39 ][ 1 ],
   alphaCSR[ 39 ][ 2 ],
   alphaCSR[ 39 ][ 3 ],
   alphaCSR[ 39 ][ 4 ],
   alphaCSR[ 39 ][ 5 ],
   alphaCSR[ 39 ][ 6 ],
   alphaCSR[ 39 ][ 7 ],
   alphaCSR[ 39 ][ 8 ],
   alphaCSR[ 39 ][ 9 ],
   alphaCSR[ 39 ][ 10 ],
   alphaCSR[ 39 ][ 11 ],
   alphaCSR[ 39 ][ 12 ],
   alphaCSR[ 39 ][ 13 ],
   alphaCSR[ 39 ][ 14 ],
   alphaCSR[ 39 ][ 15 ],
   alphaCSR[ 39 ][ 16 ],
   alphaCSR[ 39 ][ 17 ],
   alphaCSR[ 39 ][ 18 ],
   alphaCSR[ 39 ][ 19 ],
   alphaCSR[ 39 ][ 20 ],
   alphaCSR[ 39 ][ 21 ],
   alphaCSR[ 39 ][ 22 ],
   alphaCSR[ 39 ][ 23 ],
   alphaCSR[ 39 ][ 24 ],
   alphaCSR[ 39 ][ 25 ],
   alphaCSR[ 39 ][ 26 ],
   alphaCSR[ 39 ][ 27 ],
   alphaCSR[ 39 ][ 28 ],
   alphaCSR[ 39 ][ 29 ],
   alphaCSR[ 39 ][ 30 ],
   alphaCSR[ 39 ][ 31 ],
   alphaCSR[ 39 ][ 32 ],
   alphaCSR[ 39 ][ 33 ],
   alphaCSR[ 39 ][ 34 ],
   alphaCSR[ 39 ][ 35 ],
   alphaCSR[ 39 ][ 36 ],
   alphaCSR[ 39 ][ 37 ],
   alphaCSR[ 39 ][ 38 ],
   alphaCSR[ 39 ][ 39 ],
   alphaCSR[ 39 ][ 40 ],
   alphaCSR[ 39 ][ 41 ],
   alphaCSR[ 39 ][ 42 ],
   alphaCSR[ 39 ][ 43 ],
   alphaCSR[ 39 ][ 44 ],
   alphaCSR[ 39 ][ 45 ],
   alphaCSR[ 39 ][ 46 ],
   alphaCSR[ 39 ][ 47 ],
   alphaCSR[ 39 ][ 48 ],
   alphaCSR[ 39 ][ 49 ],
   alphaCSR[ 39 ][ 50 ],
   alphaCSR[ 39 ][ 51 ],
   alphaCSR[ 39 ][ 52 ],
   alphaCSR[ 39 ][ 53 ],
   alphaCSR[ 39 ][ 54 ],
   alphaCSR[ 39 ][ 55 ],
   alphaCSR[ 39 ][ 56 ],
   alphaCSR[ 39 ][ 57 ],
   alphaCSR[ 39 ][ 58 ],
   alphaCSR[ 39 ][ 59 ],
   alphaCSR[ 39 ][ 60 ],
   alphaCSR[ 39 ][ 61 ],
   alphaCSR[ 39 ][ 62 ],
   alphaCSR[ 39 ][ 63 ],
   alphaCSR[ 39 ][ 64 ],
   alphaCSR[ 39 ][ 65 ],
   alphaCSR[ 39 ][ 66 ],
   alphaCSR[ 39 ][ 67 ],
   alphaCSR[ 39 ][ 68 ],
   alphaCSR[ 39 ][ 69 ],
   alphaCSR[ 39 ][ 70 ],
   alphaCSR[ 39 ][ 71 ],
   alphaCSR[ 39 ][ 72 ],
   alphaCSR[ 39 ][ 73 ],
   alphaCSR[ 39 ][ 74 ],
   alphaCSR[ 39 ][ 75 ],
   alphaCSR[ 39 ][ 76 ],
   alphaCSR[ 39 ][ 77 ],
   alphaCSR[ 39 ][ 78 ],
   alphaCSR[ 39 ][ 79 ],
   alphaCSR[ 39 ][ 80 ],
   alphaCSR[ 39 ][ 81 ],
   alphaCSR[ 39 ][ 82 ],
   alphaCSR[ 39 ][ 83 ],
   alphaCSR[ 39 ][ 84 ],
   alphaCSR[ 39 ][ 85 ],
   alphaCSR[ 39 ][ 86 ],
   alphaCSR[ 39 ][ 87 ],
   alphaCSR[ 39 ][ 88 ],
   alphaCSR[ 39 ][ 89 ],
   alphaCSR[ 39 ][ 90 ],
   alphaCSR[ 39 ][ 91 ],
   alphaCSR[ 39 ][ 92 ],
   alphaCSR[ 39 ][ 93 ],
   alphaCSR[ 39 ][ 94 ],
   alphaCSR[ 39 ][ 95 ],
   alphaCSR[ 39 ][ 96 ],
   alphaCSR[ 39 ][ 97 ],
   alphaCSR[ 39 ][ 98 ],
   alphaCSR[ 39 ][ 99 ],
   alphaCSR[ 39 ][ 100 ],
   alphaCSR[ 39 ][ 101 ],
   alphaCSR[ 39 ][ 102 ],
   alphaCSR[ 39 ][ 103 ],
   alphaCSR[ 39 ][ 104 ],
   alphaCSR[ 39 ][ 105 ],
   alphaCSR[ 39 ][ 106 ],
   alphaCSR[ 39 ][ 107 ],
   alphaCSR[ 39 ][ 108 ],
   alphaCSR[ 39 ][ 109 ],
   alphaCSR[ 39 ][ 110 ],
   alphaCSR[ 39 ][ 111 ],
   alphaCSR[ 39 ][ 112 ],
   alphaCSR[ 39 ][ 113 ],
   alphaCSR[ 39 ][ 114 ],
   alphaCSR[ 39 ][ 115 ],
   alphaCSR[ 39 ][ 116 ],
   alphaCSR[ 39 ][ 117 ],
   alphaCSR[ 39 ][ 118 ],
   alphaCSR[ 39 ][ 119 ],
   alphaCSR[ 39 ][ 120 ],
   alphaCSR[ 39 ][ 121 ],
   alphaCSR[ 39 ][ 122 ],
   alphaCSR[ 39 ][ 123 ],
   alphaCSR[ 39 ][ 124 ],
   alphaCSR[ 39 ][ 125 ],
   alphaCSR[ 39 ][ 126 ],
   alphaCSR[ 39 ][ 127 ],
   alphaCSR[ 39 ][ 128 ],
   alphaCSR[ 39 ][ 129 ],
   alphaCSR[ 39 ][ 130 ],
   alphaCSR[ 39 ][ 131 ],
   alphaCSR[ 39 ][ 132 ],
   alphaCSR[ 39 ][ 133 ],
   alphaCSR[ 39 ][ 134 ],
   alphaCSR[ 39 ][ 135 ],
   alphaCSR[ 39 ][ 136 ],
   alphaCSR[ 39 ][ 137 ],
   alphaCSR[ 39 ][ 138 ],
   alphaCSR[ 39 ][ 139 ],
   alphaCSR[ 39 ][ 140 ],
   alphaCSR[ 39 ][ 141 ],
   alphaCSR[ 39 ][ 142 ],
   alphaCSR[ 39 ][ 143 ],
   alphaCSR[ 39 ][ 144 ],
   alphaCSR[ 39 ][ 145 ],
   alphaCSR[ 39 ][ 146 ],
   alphaCSR[ 39 ][ 147 ],
   alphaCSR[ 39 ][ 148 ],
   alphaCSR[ 39 ][ 149 ],
   alphaCSR[ 39 ][ 150 ],
   alphaCSR[ 39 ][ 151 ],
   alphaCSR[ 39 ][ 152 ],
   alphaCSR[ 39 ][ 153 ],
   alphaCSR[ 39 ][ 154 ],
   alphaCSR[ 39 ][ 155 ],
   alphaCSR[ 39 ][ 156 ],
   alphaCSR[ 39 ][ 157 ],
   alphaCSR[ 39 ][ 158 ],
   alphaCSR[ 39 ][ 159 ],
   alphaCSR[ 39 ][ 160 ],
   alphaCSR[ 39 ][ 161 ],
   alphaCSR[ 39 ][ 162 ],
   alphaCSR[ 39 ][ 163 ],
   alphaCSR[ 39 ][ 164 ],
   alphaCSR[ 39 ][ 165 ],
   alphaCSR[ 39 ][ 166 ],
   alphaCSR[ 39 ][ 167 ],
   alphaCSR[ 39 ][ 168 ],
   alphaCSR[ 39 ][ 169 ],
   alphaCSR[ 39 ][ 170 ],
   alphaCSR[ 39 ][ 171 ],
   alphaCSR[ 39 ][ 172 ],
   alphaCSR[ 39 ][ 173 ],
   alphaCSR[ 39 ][ 174 ],
   alphaCSR[ 39 ][ 175 ],
   alphaCSR[ 39 ][ 176 ],
   alphaCSR[ 39 ][ 177 ],
   alphaCSR[ 39 ][ 178 ],
   alphaCSR[ 39 ][ 179 ],
   alphaCSR[ 39 ][ 180 ],
   alphaCSR[ 39 ][ 181 ],
   alphaCSR[ 39 ][ 182 ],
   alphaCSR[ 39 ][ 183 ],
   alphaCSR[ 39 ][ 184 ],
   alphaCSR[ 39 ][ 185 ],
   alphaCSR[ 39 ][ 186 ],
   alphaCSR[ 39 ][ 187 ],
   alphaCSR[ 39 ][ 188 ],
   alphaCSR[ 39 ][ 189 ],
   alphaCSR[ 39 ][ 190 ],
   alphaCSR[ 39 ][ 191 ],
   alphaCSR[ 39 ][ 192 ],
   alphaCSR[ 39 ][ 193 ],
   alphaCSR[ 39 ][ 194 ],
   alphaCSR[ 39 ][ 195 ],
   alphaCSR[ 39 ][ 196 ],
   alphaCSR[ 39 ][ 197 ],
   alphaCSR[ 39 ][ 198 ],
   alphaCSR[ 39 ][ 199 ],
   alphaCSR[ 39 ][ 200 ],
   alphaCSR[ 39 ][ 201 ],
   alphaCSR[ 39 ][ 202 ],
   alphaCSR[ 39 ][ 203 ],
   alphaCSR[ 39 ][ 204 ],
   alphaCSR[ 39 ][ 205 ],
   alphaCSR[ 39 ][ 206 ],
   alphaCSR[ 39 ][ 207 ],
   alphaCSR[ 39 ][ 208 ],
   alphaCSR[ 39 ][ 209 ],
   alphaCSR[ 39 ][ 210 ],
   alphaCSR[ 39 ][ 211 ],
   alphaCSR[ 39 ][ 212 ],
   alphaCSR[ 39 ][ 213 ],
   alphaCSR[ 39 ][ 214 ],
   alphaCSR[ 39 ][ 215 ],
   alphaCSR[ 39 ][ 216 ],
   alphaCSR[ 39 ][ 217 ],
   alphaCSR[ 39 ][ 218 ],
   alphaCSR[ 39 ][ 219 ],
   alphaCSR[ 39 ][ 220 ],
   alphaCSR[ 39 ][ 221 ],
   alphaCSR[ 39 ][ 222 ],
   alphaCSR[ 39 ][ 223 ],
   alphaCSR[ 39 ][ 224 ],
   alphaCSR[ 39 ][ 225 ],
   alphaCSR[ 39 ][ 226 ],
   alphaCSR[ 39 ][ 227 ],
   alphaCSR[ 39 ][ 228 ],
   alphaCSR[ 39 ][ 229 ],
   alphaCSR[ 39 ][ 230 ],
   alphaCSR[ 39 ][ 231 ],
   alphaCSR[ 39 ][ 232 ],
   alphaCSR[ 39 ][ 233 ],
   alphaCSR[ 39 ][ 234 ],
   alphaCSR[ 39 ][ 235 ],
   alphaCSR[ 39 ][ 236 ],
   alphaCSR[ 39 ][ 237 ],
   alphaCSR[ 39 ][ 238 ],
   alphaCSR[ 39 ][ 239 ],
   alphaCSR[ 39 ][ 240 ],
   alphaCSR[ 39 ][ 241 ],
   alphaCSR[ 39 ][ 242 ],
   alphaCSR[ 39 ][ 243 ],
   alphaCSR[ 39 ][ 244 ],
   alphaCSR[ 39 ][ 245 ],
   alphaCSR[ 39 ][ 246 ],
   alphaCSR[ 39 ][ 247 ],
   alphaCSR[ 39 ][ 248 ],
   alphaCSR[ 39 ][ 249 ],
   alphaCSR[ 39 ][ 250 ],
   alphaCSR[ 39 ][ 251 ],
   alphaCSR[ 39 ][ 252 ],
   alphaCSR[ 39 ][ 253 ],
   alphaCSR[ 39 ][ 254 ],
   alphaCSR[ 39 ][ 255 ],
   alphaCSR[ 39 ][ 256 ],
   alphaCSR[ 39 ][ 257 ],
   alphaCSR[ 39 ][ 258 ],
   alphaCSR[ 39 ][ 259 ],
   alphaCSR[ 39 ][ 260 ],
   alphaCSR[ 39 ][ 261 ],
   alphaCSR[ 39 ][ 262 ],
   alphaCSR[ 39 ][ 263 ],
   alphaCSR[ 39 ][ 264 ],
   alphaCSR[ 39 ][ 265 ],
   alphaCSR[ 39 ][ 266 ],
   alphaCSR[ 39 ][ 267 ],
   alphaCSR[ 39 ][ 268 ],
   alphaCSR[ 39 ][ 269 ],
   alphaCSR[ 39 ][ 270 ],
   alphaCSR[ 39 ][ 271 ],
   alphaCSR[ 39 ][ 272 ],
   alphaCSR[ 39 ][ 273 ],
   alphaCSR[ 39 ][ 274 ],
   alphaCSR[ 39 ][ 275 ],
   alphaCSR[ 39 ][ 276 ],
   alphaCSR[ 39 ][ 277 ],
   alphaCSR[ 39 ][ 278 ],
   alphaCSR[ 39 ][ 279 ],
   alphaCSR[ 39 ][ 280 ],
   alphaCSR[ 39 ][ 281 ],
   alphaCSR[ 39 ][ 282 ],
   alphaCSR[ 39 ][ 283 ],
   alphaCSR[ 39 ][ 284 ],
   alphaCSR[ 39 ][ 285 ],
   alphaCSR[ 39 ][ 286 ],
   alphaCSR[ 39 ][ 287 ],
   alphaCSR[ 39 ][ 288 ],
   alphaCSR[ 39 ][ 289 ],
   alphaCSR[ 39 ][ 290 ],
   alphaCSR[ 39 ][ 291 ],
   alphaCSR[ 39 ][ 292 ],
   alphaCSR[ 39 ][ 293 ],
   alphaCSR[ 39 ][ 294 ],
   alphaCSR[ 39 ][ 295 ],
   alphaCSR[ 39 ][ 296 ],
   alphaCSR[ 39 ][ 297 ],
   alphaCSR[ 39 ][ 298 ],
   alphaCSR[ 39 ][ 299 ],
   alphaCSR[ 39 ][ 300 ],
   alphaCSR[ 39 ][ 301 ],
   alphaCSR[ 39 ][ 302 ],
   alphaCSR[ 39 ][ 303 ],
   alphaCSR[ 39 ][ 304 ],
   alphaCSR[ 39 ][ 305 ],
   alphaCSR[ 39 ][ 306 ],
   alphaCSR[ 39 ][ 307 ],
   alphaCSR[ 39 ][ 308 ],
   alphaCSR[ 39 ][ 309 ],
   alphaCSR[ 39 ][ 310 ],
   alphaCSR[ 39 ][ 311 ],
   alphaCSR[ 39 ][ 312 ],
   alphaCSR[ 39 ][ 313 ],
   alphaCSR[ 39 ][ 314 ],
   alphaCSR[ 39 ][ 315 ],
   alphaCSR[ 39 ][ 316 ],
   alphaCSR[ 39 ][ 317 ],
   alphaCSR[ 39 ][ 318 ],
   alphaCSR[ 39 ][ 319 ],
   alphaCSR[ 39 ][ 320 ],
   alphaCSR[ 39 ][ 321 ],
   alphaCSR[ 39 ][ 322 ],
   alphaCSR[ 39 ][ 323 ],
   alphaCSR[ 39 ][ 324 ],
   alphaCSR[ 39 ][ 325 ],
   alphaCSR[ 39 ][ 326 ],
   alphaCSR[ 39 ][ 327 ],
   alphaCSR[ 39 ][ 328 ],
   alphaCSR[ 39 ][ 329 ],
   alphaCSR[ 39 ][ 330 ],
   alphaCSR[ 39 ][ 331 ],
   alphaCSR[ 39 ][ 332 ],
   alphaCSR[ 39 ][ 333 ],
   alphaCSR[ 39 ][ 334 ],
   alphaCSR[ 39 ][ 335 ],
   alphaCSR[ 39 ][ 336 ],
   alphaCSR[ 39 ][ 337 ],
   alphaCSR[ 39 ][ 338 ],
   alphaCSR[ 39 ][ 339 ],
   alphaCSR[ 39 ][ 340 ],
   alphaCSR[ 39 ][ 341 ],
   alphaCSR[ 39 ][ 342 ],
   alphaCSR[ 39 ][ 343 ],
   alphaCSR[ 39 ][ 344 ],
   alphaCSR[ 39 ][ 345 ],
   alphaCSR[ 39 ][ 346 ],
   alphaCSR[ 39 ][ 347 ],
   alphaCSR[ 39 ][ 348 ],
   alphaCSR[ 39 ][ 349 ],
   alphaCSR[ 39 ][ 350 ],
   alphaCSR[ 39 ][ 351 ],
   alphaCSR[ 39 ][ 352 ],
   alphaCSR[ 39 ][ 353 ],
   alphaCSR[ 39 ][ 354 ],
   alphaCSR[ 39 ][ 355 ],
   alphaCSR[ 39 ][ 356 ],
   alphaCSR[ 39 ][ 357 ],
   alphaCSR[ 39 ][ 358 ],
   alphaCSR[ 39 ][ 359 ],
   alphaCSR[ 39 ][ 360 ],
   alphaCSR[ 39 ][ 361 ],
   alphaCSR[ 39 ][ 362 ],
   alphaCSR[ 39 ][ 363 ],
   alphaCSR[ 39 ][ 364 ],
   alphaCSR[ 39 ][ 365 ],
   alphaCSR[ 39 ][ 366 ],
   alphaCSR[ 39 ][ 367 ],
   alphaCSR[ 39 ][ 368 ],
   alphaCSR[ 39 ][ 369 ],
   alphaCSR[ 39 ][ 370 ],
   alphaCSR[ 39 ][ 371 ],
   alphaCSR[ 39 ][ 372 ],
   alphaCSR[ 39 ][ 373 ],
   alphaCSR[ 39 ][ 374 ],
   alphaCSR[ 39 ][ 375 ],
   alphaCSR[ 39 ][ 376 ],
   alphaCSR[ 39 ][ 377 ],
   alphaCSR[ 39 ][ 378 ],
   alphaCSR[ 39 ][ 379 ],
   alphaCSR[ 39 ][ 380 ],
   alphaCSR[ 39 ][ 381 ],
   alphaCSR[ 39 ][ 382 ],
   alphaCSR[ 39 ][ 383 ],
   alphaCSR[ 40 ][ 0 ],
   alphaCSR[ 40 ][ 1 ],
   alphaCSR[ 40 ][ 2 ],
   alphaCSR[ 40 ][ 3 ],
   alphaCSR[ 40 ][ 4 ],
   alphaCSR[ 40 ][ 5 ],
   alphaCSR[ 40 ][ 6 ],
   alphaCSR[ 40 ][ 7 ],
   alphaCSR[ 40 ][ 8 ],
   alphaCSR[ 40 ][ 9 ],
   alphaCSR[ 40 ][ 10 ],
   alphaCSR[ 40 ][ 11 ],
   alphaCSR[ 40 ][ 12 ],
   alphaCSR[ 40 ][ 13 ],
   alphaCSR[ 40 ][ 14 ],
   alphaCSR[ 40 ][ 15 ],
   alphaCSR[ 40 ][ 16 ],
   alphaCSR[ 40 ][ 17 ],
   alphaCSR[ 40 ][ 18 ],
   alphaCSR[ 40 ][ 19 ],
   alphaCSR[ 40 ][ 20 ],
   alphaCSR[ 40 ][ 21 ],
   alphaCSR[ 40 ][ 22 ],
   alphaCSR[ 40 ][ 23 ],
   alphaCSR[ 40 ][ 24 ],
   alphaCSR[ 40 ][ 25 ],
   alphaCSR[ 40 ][ 26 ],
   alphaCSR[ 40 ][ 27 ],
   alphaCSR[ 40 ][ 28 ],
   alphaCSR[ 40 ][ 29 ],
   alphaCSR[ 40 ][ 30 ],
   alphaCSR[ 40 ][ 31 ],
   alphaCSR[ 40 ][ 32 ],
   alphaCSR[ 40 ][ 33 ],
   alphaCSR[ 40 ][ 34 ],
   alphaCSR[ 40 ][ 35 ],
   alphaCSR[ 40 ][ 36 ],
   alphaCSR[ 40 ][ 37 ],
   alphaCSR[ 40 ][ 38 ],
   alphaCSR[ 40 ][ 39 ],
   alphaCSR[ 40 ][ 40 ],
   alphaCSR[ 40 ][ 41 ],
   alphaCSR[ 40 ][ 42 ],
   alphaCSR[ 40 ][ 43 ],
   alphaCSR[ 40 ][ 44 ],
   alphaCSR[ 40 ][ 45 ],
   alphaCSR[ 40 ][ 46 ],
   alphaCSR[ 40 ][ 47 ],
   alphaCSR[ 40 ][ 48 ],
   alphaCSR[ 40 ][ 49 ],
   alphaCSR[ 40 ][ 50 ],
   alphaCSR[ 40 ][ 51 ],
   alphaCSR[ 40 ][ 52 ],
   alphaCSR[ 40 ][ 53 ],
   alphaCSR[ 40 ][ 54 ],
   alphaCSR[ 40 ][ 55 ],
   alphaCSR[ 40 ][ 56 ],
   alphaCSR[ 40 ][ 57 ],
   alphaCSR[ 40 ][ 58 ],
   alphaCSR[ 40 ][ 59 ],
   alphaCSR[ 40 ][ 60 ],
   alphaCSR[ 40 ][ 61 ],
   alphaCSR[ 40 ][ 62 ],
   alphaCSR[ 40 ][ 63 ],
   alphaCSR[ 40 ][ 64 ],
   alphaCSR[ 40 ][ 65 ],
   alphaCSR[ 40 ][ 66 ],
   alphaCSR[ 40 ][ 67 ],
   alphaCSR[ 40 ][ 68 ],
   alphaCSR[ 40 ][ 69 ],
   alphaCSR[ 40 ][ 70 ],
   alphaCSR[ 40 ][ 71 ],
   alphaCSR[ 40 ][ 72 ],
   alphaCSR[ 40 ][ 73 ],
   alphaCSR[ 40 ][ 74 ],
   alphaCSR[ 40 ][ 75 ],
   alphaCSR[ 40 ][ 76 ],
   alphaCSR[ 40 ][ 77 ],
   alphaCSR[ 40 ][ 78 ],
   alphaCSR[ 40 ][ 79 ],
   alphaCSR[ 40 ][ 80 ],
   alphaCSR[ 40 ][ 81 ],
   alphaCSR[ 40 ][ 82 ],
   alphaCSR[ 40 ][ 83 ],
   alphaCSR[ 40 ][ 84 ],
   alphaCSR[ 40 ][ 85 ],
   alphaCSR[ 40 ][ 86 ],
   alphaCSR[ 40 ][ 87 ],
   alphaCSR[ 40 ][ 88 ],
   alphaCSR[ 40 ][ 89 ],
   alphaCSR[ 40 ][ 90 ],
   alphaCSR[ 40 ][ 91 ],
   alphaCSR[ 40 ][ 92 ],
   alphaCSR[ 40 ][ 93 ],
   alphaCSR[ 40 ][ 94 ],
   alphaCSR[ 40 ][ 95 ],
   alphaCSR[ 40 ][ 96 ],
   alphaCSR[ 40 ][ 97 ],
   alphaCSR[ 40 ][ 98 ],
   alphaCSR[ 40 ][ 99 ],
   alphaCSR[ 40 ][ 100 ],
   alphaCSR[ 40 ][ 101 ],
   alphaCSR[ 40 ][ 102 ],
   alphaCSR[ 40 ][ 103 ],
   alphaCSR[ 40 ][ 104 ],
   alphaCSR[ 40 ][ 105 ],
   alphaCSR[ 40 ][ 106 ],
   alphaCSR[ 40 ][ 107 ],
   alphaCSR[ 40 ][ 108 ],
   alphaCSR[ 40 ][ 109 ],
   alphaCSR[ 40 ][ 110 ],
   alphaCSR[ 40 ][ 111 ],
   alphaCSR[ 40 ][ 112 ],
   alphaCSR[ 40 ][ 113 ],
   alphaCSR[ 40 ][ 114 ],
   alphaCSR[ 40 ][ 115 ],
   alphaCSR[ 40 ][ 116 ],
   alphaCSR[ 40 ][ 117 ],
   alphaCSR[ 40 ][ 118 ],
   alphaCSR[ 40 ][ 119 ],
   alphaCSR[ 40 ][ 120 ],
   alphaCSR[ 40 ][ 121 ],
   alphaCSR[ 40 ][ 122 ],
   alphaCSR[ 40 ][ 123 ],
   alphaCSR[ 40 ][ 124 ],
   alphaCSR[ 40 ][ 125 ],
   alphaCSR[ 40 ][ 126 ],
   alphaCSR[ 40 ][ 127 ],
   alphaCSR[ 40 ][ 128 ],
   alphaCSR[ 40 ][ 129 ],
   alphaCSR[ 40 ][ 130 ],
   alphaCSR[ 40 ][ 131 ],
   alphaCSR[ 40 ][ 132 ],
   alphaCSR[ 40 ][ 133 ],
   alphaCSR[ 40 ][ 134 ],
   alphaCSR[ 40 ][ 135 ],
   alphaCSR[ 40 ][ 136 ],
   alphaCSR[ 40 ][ 137 ],
   alphaCSR[ 40 ][ 138 ],
   alphaCSR[ 40 ][ 139 ],
   alphaCSR[ 40 ][ 140 ],
   alphaCSR[ 40 ][ 141 ],
   alphaCSR[ 40 ][ 142 ],
   alphaCSR[ 40 ][ 143 ],
   alphaCSR[ 40 ][ 144 ],
   alphaCSR[ 40 ][ 145 ],
   alphaCSR[ 40 ][ 146 ],
   alphaCSR[ 40 ][ 147 ],
   alphaCSR[ 40 ][ 148 ],
   alphaCSR[ 40 ][ 149 ],
   alphaCSR[ 40 ][ 150 ],
   alphaCSR[ 40 ][ 151 ],
   alphaCSR[ 40 ][ 152 ],
   alphaCSR[ 40 ][ 153 ],
   alphaCSR[ 40 ][ 154 ],
   alphaCSR[ 40 ][ 155 ],
   alphaCSR[ 40 ][ 156 ],
   alphaCSR[ 40 ][ 157 ],
   alphaCSR[ 40 ][ 158 ],
   alphaCSR[ 40 ][ 159 ],
   alphaCSR[ 40 ][ 160 ],
   alphaCSR[ 40 ][ 161 ],
   alphaCSR[ 40 ][ 162 ],
   alphaCSR[ 40 ][ 163 ],
   alphaCSR[ 40 ][ 164 ],
   alphaCSR[ 40 ][ 165 ],
   alphaCSR[ 40 ][ 166 ],
   alphaCSR[ 40 ][ 167 ],
   alphaCSR[ 40 ][ 168 ],
   alphaCSR[ 40 ][ 169 ],
   alphaCSR[ 40 ][ 170 ],
   alphaCSR[ 40 ][ 171 ],
   alphaCSR[ 40 ][ 172 ],
   alphaCSR[ 40 ][ 173 ],
   alphaCSR[ 40 ][ 174 ],
   alphaCSR[ 40 ][ 175 ],
   alphaCSR[ 40 ][ 176 ],
   alphaCSR[ 40 ][ 177 ],
   alphaCSR[ 40 ][ 178 ],
   alphaCSR[ 40 ][ 179 ],
   alphaCSR[ 40 ][ 180 ],
   alphaCSR[ 40 ][ 181 ],
   alphaCSR[ 40 ][ 182 ],
   alphaCSR[ 40 ][ 183 ],
   alphaCSR[ 40 ][ 184 ],
   alphaCSR[ 40 ][ 185 ],
   alphaCSR[ 40 ][ 186 ],
   alphaCSR[ 40 ][ 187 ],
   alphaCSR[ 40 ][ 188 ],
   alphaCSR[ 40 ][ 189 ],
   alphaCSR[ 40 ][ 190 ],
   alphaCSR[ 40 ][ 191 ],
   alphaCSR[ 40 ][ 192 ],
   alphaCSR[ 40 ][ 193 ],
   alphaCSR[ 40 ][ 194 ],
   alphaCSR[ 40 ][ 195 ],
   alphaCSR[ 40 ][ 196 ],
   alphaCSR[ 40 ][ 197 ],
   alphaCSR[ 40 ][ 198 ],
   alphaCSR[ 40 ][ 199 ],
   alphaCSR[ 40 ][ 200 ],
   alphaCSR[ 40 ][ 201 ],
   alphaCSR[ 40 ][ 202 ],
   alphaCSR[ 40 ][ 203 ],
   alphaCSR[ 40 ][ 204 ],
   alphaCSR[ 40 ][ 205 ],
   alphaCSR[ 40 ][ 206 ],
   alphaCSR[ 40 ][ 207 ],
   alphaCSR[ 40 ][ 208 ],
   alphaCSR[ 40 ][ 209 ],
   alphaCSR[ 40 ][ 210 ],
   alphaCSR[ 40 ][ 211 ],
   alphaCSR[ 40 ][ 212 ],
   alphaCSR[ 40 ][ 213 ],
   alphaCSR[ 40 ][ 214 ],
   alphaCSR[ 40 ][ 215 ],
   alphaCSR[ 40 ][ 216 ],
   alphaCSR[ 40 ][ 217 ],
   alphaCSR[ 40 ][ 218 ],
   alphaCSR[ 40 ][ 219 ],
   alphaCSR[ 40 ][ 220 ],
   alphaCSR[ 40 ][ 221 ],
   alphaCSR[ 40 ][ 222 ],
   alphaCSR[ 40 ][ 223 ],
   alphaCSR[ 40 ][ 224 ],
   alphaCSR[ 40 ][ 225 ],
   alphaCSR[ 40 ][ 226 ],
   alphaCSR[ 40 ][ 227 ],
   alphaCSR[ 40 ][ 228 ],
   alphaCSR[ 40 ][ 229 ],
   alphaCSR[ 40 ][ 230 ],
   alphaCSR[ 40 ][ 231 ],
   alphaCSR[ 40 ][ 232 ],
   alphaCSR[ 40 ][ 233 ],
   alphaCSR[ 40 ][ 234 ],
   alphaCSR[ 40 ][ 235 ],
   alphaCSR[ 40 ][ 236 ],
   alphaCSR[ 40 ][ 237 ],
   alphaCSR[ 40 ][ 238 ],
   alphaCSR[ 40 ][ 239 ],
   alphaCSR[ 40 ][ 240 ],
   alphaCSR[ 40 ][ 241 ],
   alphaCSR[ 40 ][ 242 ],
   alphaCSR[ 40 ][ 243 ],
   alphaCSR[ 40 ][ 244 ],
   alphaCSR[ 40 ][ 245 ],
   alphaCSR[ 40 ][ 246 ],
   alphaCSR[ 40 ][ 247 ],
   alphaCSR[ 40 ][ 248 ],
   alphaCSR[ 40 ][ 249 ],
   alphaCSR[ 40 ][ 250 ],
   alphaCSR[ 40 ][ 251 ],
   alphaCSR[ 40 ][ 252 ],
   alphaCSR[ 40 ][ 253 ],
   alphaCSR[ 40 ][ 254 ],
   alphaCSR[ 40 ][ 255 ],
   alphaCSR[ 40 ][ 256 ],
   alphaCSR[ 40 ][ 257 ],
   alphaCSR[ 40 ][ 258 ],
   alphaCSR[ 40 ][ 259 ],
   alphaCSR[ 40 ][ 260 ],
   alphaCSR[ 40 ][ 261 ],
   alphaCSR[ 40 ][ 262 ],
   alphaCSR[ 40 ][ 263 ],
   alphaCSR[ 40 ][ 264 ],
   alphaCSR[ 40 ][ 265 ],
   alphaCSR[ 40 ][ 266 ],
   alphaCSR[ 40 ][ 267 ],
   alphaCSR[ 40 ][ 268 ],
   alphaCSR[ 40 ][ 269 ],
   alphaCSR[ 40 ][ 270 ],
   alphaCSR[ 40 ][ 271 ],
   alphaCSR[ 40 ][ 272 ],
   alphaCSR[ 40 ][ 273 ],
   alphaCSR[ 40 ][ 274 ],
   alphaCSR[ 40 ][ 275 ],
   alphaCSR[ 40 ][ 276 ],
   alphaCSR[ 40 ][ 277 ],
   alphaCSR[ 40 ][ 278 ],
   alphaCSR[ 40 ][ 279 ],
   alphaCSR[ 40 ][ 280 ],
   alphaCSR[ 40 ][ 281 ],
   alphaCSR[ 40 ][ 282 ],
   alphaCSR[ 40 ][ 283 ],
   alphaCSR[ 40 ][ 284 ],
   alphaCSR[ 40 ][ 285 ],
   alphaCSR[ 40 ][ 286 ],
   alphaCSR[ 40 ][ 287 ],
   alphaCSR[ 40 ][ 288 ],
   alphaCSR[ 40 ][ 289 ],
   alphaCSR[ 40 ][ 290 ],
   alphaCSR[ 40 ][ 291 ],
   alphaCSR[ 40 ][ 292 ],
   alphaCSR[ 40 ][ 293 ],
   alphaCSR[ 40 ][ 294 ],
   alphaCSR[ 40 ][ 295 ],
   alphaCSR[ 40 ][ 296 ],
   alphaCSR[ 40 ][ 297 ],
   alphaCSR[ 40 ][ 298 ],
   alphaCSR[ 40 ][ 299 ],
   alphaCSR[ 40 ][ 300 ],
   alphaCSR[ 40 ][ 301 ],
   alphaCSR[ 40 ][ 302 ],
   alphaCSR[ 40 ][ 303 ],
   alphaCSR[ 40 ][ 304 ],
   alphaCSR[ 40 ][ 305 ],
   alphaCSR[ 40 ][ 306 ],
   alphaCSR[ 40 ][ 307 ],
   alphaCSR[ 40 ][ 308 ],
   alphaCSR[ 40 ][ 309 ],
   alphaCSR[ 40 ][ 310 ],
   alphaCSR[ 40 ][ 311 ],
   alphaCSR[ 40 ][ 312 ],
   alphaCSR[ 40 ][ 313 ],
   alphaCSR[ 40 ][ 314 ],
   alphaCSR[ 40 ][ 315 ],
   alphaCSR[ 40 ][ 316 ],
   alphaCSR[ 40 ][ 317 ],
   alphaCSR[ 40 ][ 318 ],
   alphaCSR[ 40 ][ 319 ],
   alphaCSR[ 40 ][ 320 ],
   alphaCSR[ 40 ][ 321 ],
   alphaCSR[ 40 ][ 322 ],
   alphaCSR[ 40 ][ 323 ],
   alphaCSR[ 40 ][ 324 ],
   alphaCSR[ 40 ][ 325 ],
   alphaCSR[ 40 ][ 326 ],
   alphaCSR[ 40 ][ 327 ],
   alphaCSR[ 40 ][ 328 ],
   alphaCSR[ 40 ][ 329 ],
   alphaCSR[ 40 ][ 330 ],
   alphaCSR[ 40 ][ 331 ],
   alphaCSR[ 40 ][ 332 ],
   alphaCSR[ 40 ][ 333 ],
   alphaCSR[ 40 ][ 334 ],
   alphaCSR[ 40 ][ 335 ],
   alphaCSR[ 40 ][ 336 ],
   alphaCSR[ 40 ][ 337 ],
   alphaCSR[ 40 ][ 338 ],
   alphaCSR[ 40 ][ 339 ],
   alphaCSR[ 40 ][ 340 ],
   alphaCSR[ 40 ][ 341 ],
   alphaCSR[ 40 ][ 342 ],
   alphaCSR[ 40 ][ 343 ],
   alphaCSR[ 40 ][ 344 ],
   alphaCSR[ 40 ][ 345 ],
   alphaCSR[ 40 ][ 346 ],
   alphaCSR[ 40 ][ 347 ],
   alphaCSR[ 40 ][ 348 ],
   alphaCSR[ 40 ][ 349 ],
   alphaCSR[ 40 ][ 350 ],
   alphaCSR[ 40 ][ 351 ],
   alphaCSR[ 40 ][ 352 ],
   alphaCSR[ 40 ][ 353 ],
   alphaCSR[ 40 ][ 354 ],
   alphaCSR[ 40 ][ 355 ],
   alphaCSR[ 40 ][ 356 ],
   alphaCSR[ 40 ][ 357 ],
   alphaCSR[ 40 ][ 358 ],
   alphaCSR[ 40 ][ 359 ],
   alphaCSR[ 40 ][ 360 ],
   alphaCSR[ 40 ][ 361 ],
   alphaCSR[ 40 ][ 362 ],
   alphaCSR[ 40 ][ 363 ],
   alphaCSR[ 40 ][ 364 ],
   alphaCSR[ 40 ][ 365 ],
   alphaCSR[ 40 ][ 366 ],
   alphaCSR[ 40 ][ 367 ],
   alphaCSR[ 40 ][ 368 ],
   alphaCSR[ 40 ][ 369 ],
   alphaCSR[ 40 ][ 370 ],
   alphaCSR[ 40 ][ 371 ],
   alphaCSR[ 40 ][ 372 ],
   alphaCSR[ 40 ][ 373 ],
   alphaCSR[ 40 ][ 374 ],
   alphaCSR[ 40 ][ 375 ],
   alphaCSR[ 40 ][ 376 ],
   alphaCSR[ 40 ][ 377 ],
   alphaCSR[ 40 ][ 378 ],
   alphaCSR[ 40 ][ 379 ],
   alphaCSR[ 40 ][ 380 ],
   alphaCSR[ 40 ][ 381 ],
   alphaCSR[ 40 ][ 382 ],
   alphaCSR[ 40 ][ 383 ],
   alphaCSR[ 41 ][ 0 ],
   alphaCSR[ 41 ][ 1 ],
   alphaCSR[ 41 ][ 2 ],
   alphaCSR[ 41 ][ 3 ],
   alphaCSR[ 41 ][ 4 ],
   alphaCSR[ 41 ][ 5 ],
   alphaCSR[ 41 ][ 6 ],
   alphaCSR[ 41 ][ 7 ],
   alphaCSR[ 41 ][ 8 ],
   alphaCSR[ 41 ][ 9 ],
   alphaCSR[ 41 ][ 10 ],
   alphaCSR[ 41 ][ 11 ],
   alphaCSR[ 41 ][ 12 ],
   alphaCSR[ 41 ][ 13 ],
   alphaCSR[ 41 ][ 14 ],
   alphaCSR[ 41 ][ 15 ],
   alphaCSR[ 41 ][ 16 ],
   alphaCSR[ 41 ][ 17 ],
   alphaCSR[ 41 ][ 18 ],
   alphaCSR[ 41 ][ 19 ],
   alphaCSR[ 41 ][ 20 ],
   alphaCSR[ 41 ][ 21 ],
   alphaCSR[ 41 ][ 22 ],
   alphaCSR[ 41 ][ 23 ],
   alphaCSR[ 41 ][ 24 ],
   alphaCSR[ 41 ][ 25 ],
   alphaCSR[ 41 ][ 26 ],
   alphaCSR[ 41 ][ 27 ],
   alphaCSR[ 41 ][ 28 ],
   alphaCSR[ 41 ][ 29 ],
   alphaCSR[ 41 ][ 30 ],
   alphaCSR[ 41 ][ 31 ],
   alphaCSR[ 41 ][ 32 ],
   alphaCSR[ 41 ][ 33 ],
   alphaCSR[ 41 ][ 34 ],
   alphaCSR[ 41 ][ 35 ],
   alphaCSR[ 41 ][ 36 ],
   alphaCSR[ 41 ][ 37 ],
   alphaCSR[ 41 ][ 38 ],
   alphaCSR[ 41 ][ 39 ],
   alphaCSR[ 41 ][ 40 ],
   alphaCSR[ 41 ][ 41 ],
   alphaCSR[ 41 ][ 42 ],
   alphaCSR[ 41 ][ 43 ],
   alphaCSR[ 41 ][ 44 ],
   alphaCSR[ 41 ][ 45 ],
   alphaCSR[ 41 ][ 46 ],
   alphaCSR[ 41 ][ 47 ],
   alphaCSR[ 41 ][ 48 ],
   alphaCSR[ 41 ][ 49 ],
   alphaCSR[ 41 ][ 50 ],
   alphaCSR[ 41 ][ 51 ],
   alphaCSR[ 41 ][ 52 ],
   alphaCSR[ 41 ][ 53 ],
   alphaCSR[ 41 ][ 54 ],
   alphaCSR[ 41 ][ 55 ],
   alphaCSR[ 41 ][ 56 ],
   alphaCSR[ 41 ][ 57 ],
   alphaCSR[ 41 ][ 58 ],
   alphaCSR[ 41 ][ 59 ],
   alphaCSR[ 41 ][ 60 ],
   alphaCSR[ 41 ][ 61 ],
   alphaCSR[ 41 ][ 62 ],
   alphaCSR[ 41 ][ 63 ],
   alphaCSR[ 41 ][ 64 ],
   alphaCSR[ 41 ][ 65 ],
   alphaCSR[ 41 ][ 66 ],
   alphaCSR[ 41 ][ 67 ],
   alphaCSR[ 41 ][ 68 ],
   alphaCSR[ 41 ][ 69 ],
   alphaCSR[ 41 ][ 70 ],
   alphaCSR[ 41 ][ 71 ],
   alphaCSR[ 41 ][ 72 ],
   alphaCSR[ 41 ][ 73 ],
   alphaCSR[ 41 ][ 74 ],
   alphaCSR[ 41 ][ 75 ],
   alphaCSR[ 41 ][ 76 ],
   alphaCSR[ 41 ][ 77 ],
   alphaCSR[ 41 ][ 78 ],
   alphaCSR[ 41 ][ 79 ],
   alphaCSR[ 41 ][ 80 ],
   alphaCSR[ 41 ][ 81 ],
   alphaCSR[ 41 ][ 82 ],
   alphaCSR[ 41 ][ 83 ],
   alphaCSR[ 41 ][ 84 ],
   alphaCSR[ 41 ][ 85 ],
   alphaCSR[ 41 ][ 86 ],
   alphaCSR[ 41 ][ 87 ],
   alphaCSR[ 41 ][ 88 ],
   alphaCSR[ 41 ][ 89 ],
   alphaCSR[ 41 ][ 90 ],
   alphaCSR[ 41 ][ 91 ],
   alphaCSR[ 41 ][ 92 ],
   alphaCSR[ 41 ][ 93 ],
   alphaCSR[ 41 ][ 94 ],
   alphaCSR[ 41 ][ 95 ],
   alphaCSR[ 41 ][ 96 ],
   alphaCSR[ 41 ][ 97 ],
   alphaCSR[ 41 ][ 98 ],
   alphaCSR[ 41 ][ 99 ],
   alphaCSR[ 41 ][ 100 ],
   alphaCSR[ 41 ][ 101 ],
   alphaCSR[ 41 ][ 102 ],
   alphaCSR[ 41 ][ 103 ],
   alphaCSR[ 41 ][ 104 ],
   alphaCSR[ 41 ][ 105 ],
   alphaCSR[ 41 ][ 106 ],
   alphaCSR[ 41 ][ 107 ],
   alphaCSR[ 41 ][ 108 ],
   alphaCSR[ 41 ][ 109 ],
   alphaCSR[ 41 ][ 110 ],
   alphaCSR[ 41 ][ 111 ],
   alphaCSR[ 41 ][ 112 ],
   alphaCSR[ 41 ][ 113 ],
   alphaCSR[ 41 ][ 114 ],
   alphaCSR[ 41 ][ 115 ],
   alphaCSR[ 41 ][ 116 ],
   alphaCSR[ 41 ][ 117 ],
   alphaCSR[ 41 ][ 118 ],
   alphaCSR[ 41 ][ 119 ],
   alphaCSR[ 41 ][ 120 ],
   alphaCSR[ 41 ][ 121 ],
   alphaCSR[ 41 ][ 122 ],
   alphaCSR[ 41 ][ 123 ],
   alphaCSR[ 41 ][ 124 ],
   alphaCSR[ 41 ][ 125 ],
   alphaCSR[ 41 ][ 126 ],
   alphaCSR[ 41 ][ 127 ],
   alphaCSR[ 41 ][ 128 ],
   alphaCSR[ 41 ][ 129 ],
   alphaCSR[ 41 ][ 130 ],
   alphaCSR[ 41 ][ 131 ],
   alphaCSR[ 41 ][ 132 ],
   alphaCSR[ 41 ][ 133 ],
   alphaCSR[ 41 ][ 134 ],
   alphaCSR[ 41 ][ 135 ],
   alphaCSR[ 41 ][ 136 ],
   alphaCSR[ 41 ][ 137 ],
   alphaCSR[ 41 ][ 138 ],
   alphaCSR[ 41 ][ 139 ],
   alphaCSR[ 41 ][ 140 ],
   alphaCSR[ 41 ][ 141 ],
   alphaCSR[ 41 ][ 142 ],
   alphaCSR[ 41 ][ 143 ],
   alphaCSR[ 41 ][ 144 ],
   alphaCSR[ 41 ][ 145 ],
   alphaCSR[ 41 ][ 146 ],
   alphaCSR[ 41 ][ 147 ],
   alphaCSR[ 41 ][ 148 ],
   alphaCSR[ 41 ][ 149 ],
   alphaCSR[ 41 ][ 150 ],
   alphaCSR[ 41 ][ 151 ],
   alphaCSR[ 41 ][ 152 ],
   alphaCSR[ 41 ][ 153 ],
   alphaCSR[ 41 ][ 154 ],
   alphaCSR[ 41 ][ 155 ],
   alphaCSR[ 41 ][ 156 ],
   alphaCSR[ 41 ][ 157 ],
   alphaCSR[ 41 ][ 158 ],
   alphaCSR[ 41 ][ 159 ],
   alphaCSR[ 41 ][ 160 ],
   alphaCSR[ 41 ][ 161 ],
   alphaCSR[ 41 ][ 162 ],
   alphaCSR[ 41 ][ 163 ],
   alphaCSR[ 41 ][ 164 ],
   alphaCSR[ 41 ][ 165 ],
   alphaCSR[ 41 ][ 166 ],
   alphaCSR[ 41 ][ 167 ],
   alphaCSR[ 41 ][ 168 ],
   alphaCSR[ 41 ][ 169 ],
   alphaCSR[ 41 ][ 170 ],
   alphaCSR[ 41 ][ 171 ],
   alphaCSR[ 41 ][ 172 ],
   alphaCSR[ 41 ][ 173 ],
   alphaCSR[ 41 ][ 174 ],
   alphaCSR[ 41 ][ 175 ],
   alphaCSR[ 41 ][ 176 ],
   alphaCSR[ 41 ][ 177 ],
   alphaCSR[ 41 ][ 178 ],
   alphaCSR[ 41 ][ 179 ],
   alphaCSR[ 41 ][ 180 ],
   alphaCSR[ 41 ][ 181 ],
   alphaCSR[ 41 ][ 182 ],
   alphaCSR[ 41 ][ 183 ],
   alphaCSR[ 41 ][ 184 ],
   alphaCSR[ 41 ][ 185 ],
   alphaCSR[ 41 ][ 186 ],
   alphaCSR[ 41 ][ 187 ],
   alphaCSR[ 41 ][ 188 ],
   alphaCSR[ 41 ][ 189 ],
   alphaCSR[ 41 ][ 190 ],
   alphaCSR[ 41 ][ 191 ],
   alphaCSR[ 41 ][ 192 ],
   alphaCSR[ 41 ][ 193 ],
   alphaCSR[ 41 ][ 194 ],
   alphaCSR[ 41 ][ 195 ],
   alphaCSR[ 41 ][ 196 ],
   alphaCSR[ 41 ][ 197 ],
   alphaCSR[ 41 ][ 198 ],
   alphaCSR[ 41 ][ 199 ],
   alphaCSR[ 41 ][ 200 ],
   alphaCSR[ 41 ][ 201 ],
   alphaCSR[ 41 ][ 202 ],
   alphaCSR[ 41 ][ 203 ],
   alphaCSR[ 41 ][ 204 ],
   alphaCSR[ 41 ][ 205 ],
   alphaCSR[ 41 ][ 206 ],
   alphaCSR[ 41 ][ 207 ],
   alphaCSR[ 41 ][ 208 ],
   alphaCSR[ 41 ][ 209 ],
   alphaCSR[ 41 ][ 210 ],
   alphaCSR[ 41 ][ 211 ],
   alphaCSR[ 41 ][ 212 ],
   alphaCSR[ 41 ][ 213 ],
   alphaCSR[ 41 ][ 214 ],
   alphaCSR[ 41 ][ 215 ],
   alphaCSR[ 41 ][ 216 ],
   alphaCSR[ 41 ][ 217 ],
   alphaCSR[ 41 ][ 218 ],
   alphaCSR[ 41 ][ 219 ],
   alphaCSR[ 41 ][ 220 ],
   alphaCSR[ 41 ][ 221 ],
   alphaCSR[ 41 ][ 222 ],
   alphaCSR[ 41 ][ 223 ],
   alphaCSR[ 41 ][ 224 ],
   alphaCSR[ 41 ][ 225 ],
   alphaCSR[ 41 ][ 226 ],
   alphaCSR[ 41 ][ 227 ],
   alphaCSR[ 41 ][ 228 ],
   alphaCSR[ 41 ][ 229 ],
   alphaCSR[ 41 ][ 230 ],
   alphaCSR[ 41 ][ 231 ],
   alphaCSR[ 41 ][ 232 ],
   alphaCSR[ 41 ][ 233 ],
   alphaCSR[ 41 ][ 234 ],
   alphaCSR[ 41 ][ 235 ],
   alphaCSR[ 41 ][ 236 ],
   alphaCSR[ 41 ][ 237 ],
   alphaCSR[ 41 ][ 238 ],
   alphaCSR[ 41 ][ 239 ],
   alphaCSR[ 41 ][ 240 ],
   alphaCSR[ 41 ][ 241 ],
   alphaCSR[ 41 ][ 242 ],
   alphaCSR[ 41 ][ 243 ],
   alphaCSR[ 41 ][ 244 ],
   alphaCSR[ 41 ][ 245 ],
   alphaCSR[ 41 ][ 246 ],
   alphaCSR[ 41 ][ 247 ],
   alphaCSR[ 41 ][ 248 ],
   alphaCSR[ 41 ][ 249 ],
   alphaCSR[ 41 ][ 250 ],
   alphaCSR[ 41 ][ 251 ],
   alphaCSR[ 41 ][ 252 ],
   alphaCSR[ 41 ][ 253 ],
   alphaCSR[ 41 ][ 254 ],
   alphaCSR[ 41 ][ 255 ],
   alphaCSR[ 41 ][ 256 ],
   alphaCSR[ 41 ][ 257 ],
   alphaCSR[ 41 ][ 258 ],
   alphaCSR[ 41 ][ 259 ],
   alphaCSR[ 41 ][ 260 ],
   alphaCSR[ 41 ][ 261 ],
   alphaCSR[ 41 ][ 262 ],
   alphaCSR[ 41 ][ 263 ],
   alphaCSR[ 41 ][ 264 ],
   alphaCSR[ 41 ][ 265 ],
   alphaCSR[ 41 ][ 266 ],
   alphaCSR[ 41 ][ 267 ],
   alphaCSR[ 41 ][ 268 ],
   alphaCSR[ 41 ][ 269 ],
   alphaCSR[ 41 ][ 270 ],
   alphaCSR[ 41 ][ 271 ],
   alphaCSR[ 41 ][ 272 ],
   alphaCSR[ 41 ][ 273 ],
   alphaCSR[ 41 ][ 274 ],
   alphaCSR[ 41 ][ 275 ],
   alphaCSR[ 41 ][ 276 ],
   alphaCSR[ 41 ][ 277 ],
   alphaCSR[ 41 ][ 278 ],
   alphaCSR[ 41 ][ 279 ],
   alphaCSR[ 41 ][ 280 ],
   alphaCSR[ 41 ][ 281 ],
   alphaCSR[ 41 ][ 282 ],
   alphaCSR[ 41 ][ 283 ],
   alphaCSR[ 41 ][ 284 ],
   alphaCSR[ 41 ][ 285 ],
   alphaCSR[ 41 ][ 286 ],
   alphaCSR[ 41 ][ 287 ],
   alphaCSR[ 41 ][ 288 ],
   alphaCSR[ 41 ][ 289 ],
   alphaCSR[ 41 ][ 290 ],
   alphaCSR[ 41 ][ 291 ],
   alphaCSR[ 41 ][ 292 ],
   alphaCSR[ 41 ][ 293 ],
   alphaCSR[ 41 ][ 294 ],
   alphaCSR[ 41 ][ 295 ],
   alphaCSR[ 41 ][ 296 ],
   alphaCSR[ 41 ][ 297 ],
   alphaCSR[ 41 ][ 298 ],
   alphaCSR[ 41 ][ 299 ],
   alphaCSR[ 41 ][ 300 ],
   alphaCSR[ 41 ][ 301 ],
   alphaCSR[ 41 ][ 302 ],
   alphaCSR[ 41 ][ 303 ],
   alphaCSR[ 41 ][ 304 ],
   alphaCSR[ 41 ][ 305 ],
   alphaCSR[ 41 ][ 306 ],
   alphaCSR[ 41 ][ 307 ],
   alphaCSR[ 41 ][ 308 ],
   alphaCSR[ 41 ][ 309 ],
   alphaCSR[ 41 ][ 310 ],
   alphaCSR[ 41 ][ 311 ],
   alphaCSR[ 41 ][ 312 ],
   alphaCSR[ 41 ][ 313 ],
   alphaCSR[ 41 ][ 314 ],
   alphaCSR[ 41 ][ 315 ],
   alphaCSR[ 41 ][ 316 ],
   alphaCSR[ 41 ][ 317 ],
   alphaCSR[ 41 ][ 318 ],
   alphaCSR[ 41 ][ 319 ],
   alphaCSR[ 41 ][ 320 ],
   alphaCSR[ 41 ][ 321 ],
   alphaCSR[ 41 ][ 322 ],
   alphaCSR[ 41 ][ 323 ],
   alphaCSR[ 41 ][ 324 ],
   alphaCSR[ 41 ][ 325 ],
   alphaCSR[ 41 ][ 326 ],
   alphaCSR[ 41 ][ 327 ],
   alphaCSR[ 41 ][ 328 ],
   alphaCSR[ 41 ][ 329 ],
   alphaCSR[ 41 ][ 330 ],
   alphaCSR[ 41 ][ 331 ],
   alphaCSR[ 41 ][ 332 ],
   alphaCSR[ 41 ][ 333 ],
   alphaCSR[ 41 ][ 334 ],
   alphaCSR[ 41 ][ 335 ],
   alphaCSR[ 41 ][ 336 ],
   alphaCSR[ 41 ][ 337 ],
   alphaCSR[ 41 ][ 338 ],
   alphaCSR[ 41 ][ 339 ],
   alphaCSR[ 41 ][ 340 ],
   alphaCSR[ 41 ][ 341 ],
   alphaCSR[ 41 ][ 342 ],
   alphaCSR[ 41 ][ 343 ],
   alphaCSR[ 41 ][ 344 ],
   alphaCSR[ 41 ][ 345 ],
   alphaCSR[ 41 ][ 346 ],
   alphaCSR[ 41 ][ 347 ],
   alphaCSR[ 41 ][ 348 ],
   alphaCSR[ 41 ][ 349 ],
   alphaCSR[ 41 ][ 350 ],
   alphaCSR[ 41 ][ 351 ],
   alphaCSR[ 41 ][ 352 ],
   alphaCSR[ 41 ][ 353 ],
   alphaCSR[ 41 ][ 354 ],
   alphaCSR[ 41 ][ 355 ],
   alphaCSR[ 41 ][ 356 ],
   alphaCSR[ 41 ][ 357 ],
   alphaCSR[ 41 ][ 358 ],
   alphaCSR[ 41 ][ 359 ],
   alphaCSR[ 41 ][ 360 ],
   alphaCSR[ 41 ][ 361 ],
   alphaCSR[ 41 ][ 362 ],
   alphaCSR[ 41 ][ 363 ],
   alphaCSR[ 41 ][ 364 ],
   alphaCSR[ 41 ][ 365 ],
   alphaCSR[ 41 ][ 366 ],
   alphaCSR[ 41 ][ 367 ],
   alphaCSR[ 41 ][ 368 ],
   alphaCSR[ 41 ][ 369 ],
   alphaCSR[ 41 ][ 370 ],
   alphaCSR[ 41 ][ 371 ],
   alphaCSR[ 41 ][ 372 ],
   alphaCSR[ 41 ][ 373 ],
   alphaCSR[ 41 ][ 374 ],
   alphaCSR[ 41 ][ 375 ],
   alphaCSR[ 41 ][ 376 ],
   alphaCSR[ 41 ][ 377 ],
   alphaCSR[ 41 ][ 378 ],
   alphaCSR[ 41 ][ 379 ],
   alphaCSR[ 41 ][ 380 ],
   alphaCSR[ 41 ][ 381 ],
   alphaCSR[ 41 ][ 382 ],
   alphaCSR[ 41 ][ 383 ],
   alphaCSR[ 42 ][ 0 ],
   alphaCSR[ 42 ][ 1 ],
   alphaCSR[ 42 ][ 2 ],
   alphaCSR[ 42 ][ 3 ],
   alphaCSR[ 42 ][ 4 ],
   alphaCSR[ 42 ][ 5 ],
   alphaCSR[ 42 ][ 6 ],
   alphaCSR[ 42 ][ 7 ],
   alphaCSR[ 42 ][ 8 ],
   alphaCSR[ 42 ][ 9 ],
   alphaCSR[ 42 ][ 10 ],
   alphaCSR[ 42 ][ 11 ],
   alphaCSR[ 42 ][ 12 ],
   alphaCSR[ 42 ][ 13 ],
   alphaCSR[ 42 ][ 14 ],
   alphaCSR[ 42 ][ 15 ],
   alphaCSR[ 42 ][ 16 ],
   alphaCSR[ 42 ][ 17 ],
   alphaCSR[ 42 ][ 18 ],
   alphaCSR[ 42 ][ 19 ],
   alphaCSR[ 42 ][ 20 ],
   alphaCSR[ 42 ][ 21 ],
   alphaCSR[ 42 ][ 22 ],
   alphaCSR[ 42 ][ 23 ],
   alphaCSR[ 42 ][ 24 ],
   alphaCSR[ 42 ][ 25 ],
   alphaCSR[ 42 ][ 26 ],
   alphaCSR[ 42 ][ 27 ],
   alphaCSR[ 42 ][ 28 ],
   alphaCSR[ 42 ][ 29 ],
   alphaCSR[ 42 ][ 30 ],
   alphaCSR[ 42 ][ 31 ],
   alphaCSR[ 42 ][ 32 ],
   alphaCSR[ 42 ][ 33 ],
   alphaCSR[ 42 ][ 34 ],
   alphaCSR[ 42 ][ 35 ],
   alphaCSR[ 42 ][ 36 ],
   alphaCSR[ 42 ][ 37 ],
   alphaCSR[ 42 ][ 38 ],
   alphaCSR[ 42 ][ 39 ],
   alphaCSR[ 42 ][ 40 ],
   alphaCSR[ 42 ][ 41 ],
   alphaCSR[ 42 ][ 42 ],
   alphaCSR[ 42 ][ 43 ],
   alphaCSR[ 42 ][ 44 ],
   alphaCSR[ 42 ][ 45 ],
   alphaCSR[ 42 ][ 46 ],
   alphaCSR[ 42 ][ 47 ],
   alphaCSR[ 42 ][ 48 ],
   alphaCSR[ 42 ][ 49 ],
   alphaCSR[ 42 ][ 50 ],
   alphaCSR[ 42 ][ 51 ],
   alphaCSR[ 42 ][ 52 ],
   alphaCSR[ 42 ][ 53 ],
   alphaCSR[ 42 ][ 54 ],
   alphaCSR[ 42 ][ 55 ],
   alphaCSR[ 42 ][ 56 ],
   alphaCSR[ 42 ][ 57 ],
   alphaCSR[ 42 ][ 58 ],
   alphaCSR[ 42 ][ 59 ],
   alphaCSR[ 42 ][ 60 ],
   alphaCSR[ 42 ][ 61 ],
   alphaCSR[ 42 ][ 62 ],
   alphaCSR[ 42 ][ 63 ],
   alphaCSR[ 42 ][ 64 ],
   alphaCSR[ 42 ][ 65 ],
   alphaCSR[ 42 ][ 66 ],
   alphaCSR[ 42 ][ 67 ],
   alphaCSR[ 42 ][ 68 ],
   alphaCSR[ 42 ][ 69 ],
   alphaCSR[ 42 ][ 70 ],
   alphaCSR[ 42 ][ 71 ],
   alphaCSR[ 42 ][ 72 ],
   alphaCSR[ 42 ][ 73 ],
   alphaCSR[ 42 ][ 74 ],
   alphaCSR[ 42 ][ 75 ],
   alphaCSR[ 42 ][ 76 ],
   alphaCSR[ 42 ][ 77 ],
   alphaCSR[ 42 ][ 78 ],
   alphaCSR[ 42 ][ 79 ],
   alphaCSR[ 42 ][ 80 ],
   alphaCSR[ 42 ][ 81 ],
   alphaCSR[ 42 ][ 82 ],
   alphaCSR[ 42 ][ 83 ],
   alphaCSR[ 42 ][ 84 ],
   alphaCSR[ 42 ][ 85 ],
   alphaCSR[ 42 ][ 86 ],
   alphaCSR[ 42 ][ 87 ],
   alphaCSR[ 42 ][ 88 ],
   alphaCSR[ 42 ][ 89 ],
   alphaCSR[ 42 ][ 90 ],
   alphaCSR[ 42 ][ 91 ],
   alphaCSR[ 42 ][ 92 ],
   alphaCSR[ 42 ][ 93 ],
   alphaCSR[ 42 ][ 94 ],
   alphaCSR[ 42 ][ 95 ],
   alphaCSR[ 42 ][ 96 ],
   alphaCSR[ 42 ][ 97 ],
   alphaCSR[ 42 ][ 98 ],
   alphaCSR[ 42 ][ 99 ],
   alphaCSR[ 42 ][ 100 ],
   alphaCSR[ 42 ][ 101 ],
   alphaCSR[ 42 ][ 102 ],
   alphaCSR[ 42 ][ 103 ],
   alphaCSR[ 42 ][ 104 ],
   alphaCSR[ 42 ][ 105 ],
   alphaCSR[ 42 ][ 106 ],
   alphaCSR[ 42 ][ 107 ],
   alphaCSR[ 42 ][ 108 ],
   alphaCSR[ 42 ][ 109 ],
   alphaCSR[ 42 ][ 110 ],
   alphaCSR[ 42 ][ 111 ],
   alphaCSR[ 42 ][ 112 ],
   alphaCSR[ 42 ][ 113 ],
   alphaCSR[ 42 ][ 114 ],
   alphaCSR[ 42 ][ 115 ],
   alphaCSR[ 42 ][ 116 ],
   alphaCSR[ 42 ][ 117 ],
   alphaCSR[ 42 ][ 118 ],
   alphaCSR[ 42 ][ 119 ],
   alphaCSR[ 42 ][ 120 ],
   alphaCSR[ 42 ][ 121 ],
   alphaCSR[ 42 ][ 122 ],
   alphaCSR[ 42 ][ 123 ],
   alphaCSR[ 42 ][ 124 ],
   alphaCSR[ 42 ][ 125 ],
   alphaCSR[ 42 ][ 126 ],
   alphaCSR[ 42 ][ 127 ],
   alphaCSR[ 42 ][ 128 ],
   alphaCSR[ 42 ][ 129 ],
   alphaCSR[ 42 ][ 130 ],
   alphaCSR[ 42 ][ 131 ],
   alphaCSR[ 42 ][ 132 ],
   alphaCSR[ 42 ][ 133 ],
   alphaCSR[ 42 ][ 134 ],
   alphaCSR[ 42 ][ 135 ],
   alphaCSR[ 42 ][ 136 ],
   alphaCSR[ 42 ][ 137 ],
   alphaCSR[ 42 ][ 138 ],
   alphaCSR[ 42 ][ 139 ],
   alphaCSR[ 42 ][ 140 ],
   alphaCSR[ 42 ][ 141 ],
   alphaCSR[ 42 ][ 142 ],
   alphaCSR[ 42 ][ 143 ],
   alphaCSR[ 42 ][ 144 ],
   alphaCSR[ 42 ][ 145 ],
   alphaCSR[ 42 ][ 146 ],
   alphaCSR[ 42 ][ 147 ],
   alphaCSR[ 42 ][ 148 ],
   alphaCSR[ 42 ][ 149 ],
   alphaCSR[ 42 ][ 150 ],
   alphaCSR[ 42 ][ 151 ],
   alphaCSR[ 42 ][ 152 ],
   alphaCSR[ 42 ][ 153 ],
   alphaCSR[ 42 ][ 154 ],
   alphaCSR[ 42 ][ 155 ],
   alphaCSR[ 42 ][ 156 ],
   alphaCSR[ 42 ][ 157 ],
   alphaCSR[ 42 ][ 158 ],
   alphaCSR[ 42 ][ 159 ],
   alphaCSR[ 42 ][ 160 ],
   alphaCSR[ 42 ][ 161 ],
   alphaCSR[ 42 ][ 162 ],
   alphaCSR[ 42 ][ 163 ],
   alphaCSR[ 42 ][ 164 ],
   alphaCSR[ 42 ][ 165 ],
   alphaCSR[ 42 ][ 166 ],
   alphaCSR[ 42 ][ 167 ],
   alphaCSR[ 42 ][ 168 ],
   alphaCSR[ 42 ][ 169 ],
   alphaCSR[ 42 ][ 170 ],
   alphaCSR[ 42 ][ 171 ],
   alphaCSR[ 42 ][ 172 ],
   alphaCSR[ 42 ][ 173 ],
   alphaCSR[ 42 ][ 174 ],
   alphaCSR[ 42 ][ 175 ],
   alphaCSR[ 42 ][ 176 ],
   alphaCSR[ 42 ][ 177 ],
   alphaCSR[ 42 ][ 178 ],
   alphaCSR[ 42 ][ 179 ],
   alphaCSR[ 42 ][ 180 ],
   alphaCSR[ 42 ][ 181 ],
   alphaCSR[ 42 ][ 182 ],
   alphaCSR[ 42 ][ 183 ],
   alphaCSR[ 42 ][ 184 ],
   alphaCSR[ 42 ][ 185 ],
   alphaCSR[ 42 ][ 186 ],
   alphaCSR[ 42 ][ 187 ],
   alphaCSR[ 42 ][ 188 ],
   alphaCSR[ 42 ][ 189 ],
   alphaCSR[ 42 ][ 190 ],
   alphaCSR[ 42 ][ 191 ],
   alphaCSR[ 42 ][ 192 ],
   alphaCSR[ 42 ][ 193 ],
   alphaCSR[ 42 ][ 194 ],
   alphaCSR[ 42 ][ 195 ],
   alphaCSR[ 42 ][ 196 ],
   alphaCSR[ 42 ][ 197 ],
   alphaCSR[ 42 ][ 198 ],
   alphaCSR[ 42 ][ 199 ],
   alphaCSR[ 42 ][ 200 ],
   alphaCSR[ 42 ][ 201 ],
   alphaCSR[ 42 ][ 202 ],
   alphaCSR[ 42 ][ 203 ],
   alphaCSR[ 42 ][ 204 ],
   alphaCSR[ 42 ][ 205 ],
   alphaCSR[ 42 ][ 206 ],
   alphaCSR[ 42 ][ 207 ],
   alphaCSR[ 42 ][ 208 ],
   alphaCSR[ 42 ][ 209 ],
   alphaCSR[ 42 ][ 210 ],
   alphaCSR[ 42 ][ 211 ],
   alphaCSR[ 42 ][ 212 ],
   alphaCSR[ 42 ][ 213 ],
   alphaCSR[ 42 ][ 214 ],
   alphaCSR[ 42 ][ 215 ],
   alphaCSR[ 42 ][ 216 ],
   alphaCSR[ 42 ][ 217 ],
   alphaCSR[ 42 ][ 218 ],
   alphaCSR[ 42 ][ 219 ],
   alphaCSR[ 42 ][ 220 ],
   alphaCSR[ 42 ][ 221 ],
   alphaCSR[ 42 ][ 222 ],
   alphaCSR[ 42 ][ 223 ],
   alphaCSR[ 42 ][ 224 ],
   alphaCSR[ 42 ][ 225 ],
   alphaCSR[ 42 ][ 226 ],
   alphaCSR[ 42 ][ 227 ],
   alphaCSR[ 42 ][ 228 ],
   alphaCSR[ 42 ][ 229 ],
   alphaCSR[ 42 ][ 230 ],
   alphaCSR[ 42 ][ 231 ],
   alphaCSR[ 42 ][ 232 ],
   alphaCSR[ 42 ][ 233 ],
   alphaCSR[ 42 ][ 234 ],
   alphaCSR[ 42 ][ 235 ],
   alphaCSR[ 42 ][ 236 ],
   alphaCSR[ 42 ][ 237 ],
   alphaCSR[ 42 ][ 238 ],
   alphaCSR[ 42 ][ 239 ],
   alphaCSR[ 42 ][ 240 ],
   alphaCSR[ 42 ][ 241 ],
   alphaCSR[ 42 ][ 242 ],
   alphaCSR[ 42 ][ 243 ],
   alphaCSR[ 42 ][ 244 ],
   alphaCSR[ 42 ][ 245 ],
   alphaCSR[ 42 ][ 246 ],
   alphaCSR[ 42 ][ 247 ],
   alphaCSR[ 42 ][ 248 ],
   alphaCSR[ 42 ][ 249 ],
   alphaCSR[ 42 ][ 250 ],
   alphaCSR[ 42 ][ 251 ],
   alphaCSR[ 42 ][ 252 ],
   alphaCSR[ 42 ][ 253 ],
   alphaCSR[ 42 ][ 254 ],
   alphaCSR[ 42 ][ 255 ],
   alphaCSR[ 42 ][ 256 ],
   alphaCSR[ 42 ][ 257 ],
   alphaCSR[ 42 ][ 258 ],
   alphaCSR[ 42 ][ 259 ],
   alphaCSR[ 42 ][ 260 ],
   alphaCSR[ 42 ][ 261 ],
   alphaCSR[ 42 ][ 262 ],
   alphaCSR[ 42 ][ 263 ],
   alphaCSR[ 42 ][ 264 ],
   alphaCSR[ 42 ][ 265 ],
   alphaCSR[ 42 ][ 266 ],
   alphaCSR[ 42 ][ 267 ],
   alphaCSR[ 42 ][ 268 ],
   alphaCSR[ 42 ][ 269 ],
   alphaCSR[ 42 ][ 270 ],
   alphaCSR[ 42 ][ 271 ],
   alphaCSR[ 42 ][ 272 ],
   alphaCSR[ 42 ][ 273 ],
   alphaCSR[ 42 ][ 274 ],
   alphaCSR[ 42 ][ 275 ],
   alphaCSR[ 42 ][ 276 ],
   alphaCSR[ 42 ][ 277 ],
   alphaCSR[ 42 ][ 278 ],
   alphaCSR[ 42 ][ 279 ],
   alphaCSR[ 42 ][ 280 ],
   alphaCSR[ 42 ][ 281 ],
   alphaCSR[ 42 ][ 282 ],
   alphaCSR[ 42 ][ 283 ],
   alphaCSR[ 42 ][ 284 ],
   alphaCSR[ 42 ][ 285 ],
   alphaCSR[ 42 ][ 286 ],
   alphaCSR[ 42 ][ 287 ],
   alphaCSR[ 42 ][ 288 ],
   alphaCSR[ 42 ][ 289 ],
   alphaCSR[ 42 ][ 290 ],
   alphaCSR[ 42 ][ 291 ],
   alphaCSR[ 42 ][ 292 ],
   alphaCSR[ 42 ][ 293 ],
   alphaCSR[ 42 ][ 294 ],
   alphaCSR[ 42 ][ 295 ],
   alphaCSR[ 42 ][ 296 ],
   alphaCSR[ 42 ][ 297 ],
   alphaCSR[ 42 ][ 298 ],
   alphaCSR[ 42 ][ 299 ],
   alphaCSR[ 42 ][ 300 ],
   alphaCSR[ 42 ][ 301 ],
   alphaCSR[ 42 ][ 302 ],
   alphaCSR[ 42 ][ 303 ],
   alphaCSR[ 42 ][ 304 ],
   alphaCSR[ 42 ][ 305 ],
   alphaCSR[ 42 ][ 306 ],
   alphaCSR[ 42 ][ 307 ],
   alphaCSR[ 42 ][ 308 ],
   alphaCSR[ 42 ][ 309 ],
   alphaCSR[ 42 ][ 310 ],
   alphaCSR[ 42 ][ 311 ],
   alphaCSR[ 42 ][ 312 ],
   alphaCSR[ 42 ][ 313 ],
   alphaCSR[ 42 ][ 314 ],
   alphaCSR[ 42 ][ 315 ],
   alphaCSR[ 42 ][ 316 ],
   alphaCSR[ 42 ][ 317 ],
   alphaCSR[ 42 ][ 318 ],
   alphaCSR[ 42 ][ 319 ],
   alphaCSR[ 42 ][ 320 ],
   alphaCSR[ 42 ][ 321 ],
   alphaCSR[ 42 ][ 322 ],
   alphaCSR[ 42 ][ 323 ],
   alphaCSR[ 42 ][ 324 ],
   alphaCSR[ 42 ][ 325 ],
   alphaCSR[ 42 ][ 326 ],
   alphaCSR[ 42 ][ 327 ],
   alphaCSR[ 42 ][ 328 ],
   alphaCSR[ 42 ][ 329 ],
   alphaCSR[ 42 ][ 330 ],
   alphaCSR[ 42 ][ 331 ],
   alphaCSR[ 42 ][ 332 ],
   alphaCSR[ 42 ][ 333 ],
   alphaCSR[ 42 ][ 334 ],
   alphaCSR[ 42 ][ 335 ],
   alphaCSR[ 42 ][ 336 ],
   alphaCSR[ 42 ][ 337 ],
   alphaCSR[ 42 ][ 338 ],
   alphaCSR[ 42 ][ 339 ],
   alphaCSR[ 42 ][ 340 ],
   alphaCSR[ 42 ][ 341 ],
   alphaCSR[ 42 ][ 342 ],
   alphaCSR[ 42 ][ 343 ],
   alphaCSR[ 42 ][ 344 ],
   alphaCSR[ 42 ][ 345 ],
   alphaCSR[ 42 ][ 346 ],
   alphaCSR[ 42 ][ 347 ],
   alphaCSR[ 42 ][ 348 ],
   alphaCSR[ 42 ][ 349 ],
   alphaCSR[ 42 ][ 350 ],
   alphaCSR[ 42 ][ 351 ],
   alphaCSR[ 42 ][ 352 ],
   alphaCSR[ 42 ][ 353 ],
   alphaCSR[ 42 ][ 354 ],
   alphaCSR[ 42 ][ 355 ],
   alphaCSR[ 42 ][ 356 ],
   alphaCSR[ 42 ][ 357 ],
   alphaCSR[ 42 ][ 358 ],
   alphaCSR[ 42 ][ 359 ],
   alphaCSR[ 42 ][ 360 ],
   alphaCSR[ 42 ][ 361 ],
   alphaCSR[ 42 ][ 362 ],
   alphaCSR[ 42 ][ 363 ],
   alphaCSR[ 42 ][ 364 ],
   alphaCSR[ 42 ][ 365 ],
   alphaCSR[ 42 ][ 366 ],
   alphaCSR[ 42 ][ 367 ],
   alphaCSR[ 42 ][ 368 ],
   alphaCSR[ 42 ][ 369 ],
   alphaCSR[ 42 ][ 370 ],
   alphaCSR[ 42 ][ 371 ],
   alphaCSR[ 42 ][ 372 ],
   alphaCSR[ 42 ][ 373 ],
   alphaCSR[ 42 ][ 374 ],
   alphaCSR[ 42 ][ 375 ],
   alphaCSR[ 42 ][ 376 ],
   alphaCSR[ 42 ][ 377 ],
   alphaCSR[ 42 ][ 378 ],
   alphaCSR[ 42 ][ 379 ],
   alphaCSR[ 42 ][ 380 ],
   alphaCSR[ 42 ][ 381 ],
   alphaCSR[ 42 ][ 382 ],
   alphaCSR[ 42 ][ 383 ],
   alphaCSR[ 43 ][ 0 ],
   alphaCSR[ 43 ][ 1 ],
   alphaCSR[ 43 ][ 2 ],
   alphaCSR[ 43 ][ 3 ],
   alphaCSR[ 43 ][ 4 ],
   alphaCSR[ 43 ][ 5 ],
   alphaCSR[ 43 ][ 6 ],
   alphaCSR[ 43 ][ 7 ],
   alphaCSR[ 43 ][ 8 ],
   alphaCSR[ 43 ][ 9 ],
   alphaCSR[ 43 ][ 10 ],
   alphaCSR[ 43 ][ 11 ],
   alphaCSR[ 43 ][ 12 ],
   alphaCSR[ 43 ][ 13 ],
   alphaCSR[ 43 ][ 14 ],
   alphaCSR[ 43 ][ 15 ],
   alphaCSR[ 43 ][ 16 ],
   alphaCSR[ 43 ][ 17 ],
   alphaCSR[ 43 ][ 18 ],
   alphaCSR[ 43 ][ 19 ],
   alphaCSR[ 43 ][ 20 ],
   alphaCSR[ 43 ][ 21 ],
   alphaCSR[ 43 ][ 22 ],
   alphaCSR[ 43 ][ 23 ],
   alphaCSR[ 43 ][ 24 ],
   alphaCSR[ 43 ][ 25 ],
   alphaCSR[ 43 ][ 26 ],
   alphaCSR[ 43 ][ 27 ],
   alphaCSR[ 43 ][ 28 ],
   alphaCSR[ 43 ][ 29 ],
   alphaCSR[ 43 ][ 30 ],
   alphaCSR[ 43 ][ 31 ],
   alphaCSR[ 43 ][ 32 ],
   alphaCSR[ 43 ][ 33 ],
   alphaCSR[ 43 ][ 34 ],
   alphaCSR[ 43 ][ 35 ],
   alphaCSR[ 43 ][ 36 ],
   alphaCSR[ 43 ][ 37 ],
   alphaCSR[ 43 ][ 38 ],
   alphaCSR[ 43 ][ 39 ],
   alphaCSR[ 43 ][ 40 ],
   alphaCSR[ 43 ][ 41 ],
   alphaCSR[ 43 ][ 42 ],
   alphaCSR[ 43 ][ 43 ],
   alphaCSR[ 43 ][ 44 ],
   alphaCSR[ 43 ][ 45 ],
   alphaCSR[ 43 ][ 46 ],
   alphaCSR[ 43 ][ 47 ],
   alphaCSR[ 43 ][ 48 ],
   alphaCSR[ 43 ][ 49 ],
   alphaCSR[ 43 ][ 50 ],
   alphaCSR[ 43 ][ 51 ],
   alphaCSR[ 43 ][ 52 ],
   alphaCSR[ 43 ][ 53 ],
   alphaCSR[ 43 ][ 54 ],
   alphaCSR[ 43 ][ 55 ],
   alphaCSR[ 43 ][ 56 ],
   alphaCSR[ 43 ][ 57 ],
   alphaCSR[ 43 ][ 58 ],
   alphaCSR[ 43 ][ 59 ],
   alphaCSR[ 43 ][ 60 ],
   alphaCSR[ 43 ][ 61 ],
   alphaCSR[ 43 ][ 62 ],
   alphaCSR[ 43 ][ 63 ],
   alphaCSR[ 43 ][ 64 ],
   alphaCSR[ 43 ][ 65 ],
   alphaCSR[ 43 ][ 66 ],
   alphaCSR[ 43 ][ 67 ],
   alphaCSR[ 43 ][ 68 ],
   alphaCSR[ 43 ][ 69 ],
   alphaCSR[ 43 ][ 70 ],
   alphaCSR[ 43 ][ 71 ],
   alphaCSR[ 43 ][ 72 ],
   alphaCSR[ 43 ][ 73 ],
   alphaCSR[ 43 ][ 74 ],
   alphaCSR[ 43 ][ 75 ],
   alphaCSR[ 43 ][ 76 ],
   alphaCSR[ 43 ][ 77 ],
   alphaCSR[ 43 ][ 78 ],
   alphaCSR[ 43 ][ 79 ],
   alphaCSR[ 43 ][ 80 ],
   alphaCSR[ 43 ][ 81 ],
   alphaCSR[ 43 ][ 82 ],
   alphaCSR[ 43 ][ 83 ],
   alphaCSR[ 43 ][ 84 ],
   alphaCSR[ 43 ][ 85 ],
   alphaCSR[ 43 ][ 86 ],
   alphaCSR[ 43 ][ 87 ],
   alphaCSR[ 43 ][ 88 ],
   alphaCSR[ 43 ][ 89 ],
   alphaCSR[ 43 ][ 90 ],
   alphaCSR[ 43 ][ 91 ],
   alphaCSR[ 43 ][ 92 ],
   alphaCSR[ 43 ][ 93 ],
   alphaCSR[ 43 ][ 94 ],
   alphaCSR[ 43 ][ 95 ],
   alphaCSR[ 43 ][ 96 ],
   alphaCSR[ 43 ][ 97 ],
   alphaCSR[ 43 ][ 98 ],
   alphaCSR[ 43 ][ 99 ],
   alphaCSR[ 43 ][ 100 ],
   alphaCSR[ 43 ][ 101 ],
   alphaCSR[ 43 ][ 102 ],
   alphaCSR[ 43 ][ 103 ],
   alphaCSR[ 43 ][ 104 ],
   alphaCSR[ 43 ][ 105 ],
   alphaCSR[ 43 ][ 106 ],
   alphaCSR[ 43 ][ 107 ],
   alphaCSR[ 43 ][ 108 ],
   alphaCSR[ 43 ][ 109 ],
   alphaCSR[ 43 ][ 110 ],
   alphaCSR[ 43 ][ 111 ],
   alphaCSR[ 43 ][ 112 ],
   alphaCSR[ 43 ][ 113 ],
   alphaCSR[ 43 ][ 114 ],
   alphaCSR[ 43 ][ 115 ],
   alphaCSR[ 43 ][ 116 ],
   alphaCSR[ 43 ][ 117 ],
   alphaCSR[ 43 ][ 118 ],
   alphaCSR[ 43 ][ 119 ],
   alphaCSR[ 43 ][ 120 ],
   alphaCSR[ 43 ][ 121 ],
   alphaCSR[ 43 ][ 122 ],
   alphaCSR[ 43 ][ 123 ],
   alphaCSR[ 43 ][ 124 ],
   alphaCSR[ 43 ][ 125 ],
   alphaCSR[ 43 ][ 126 ],
   alphaCSR[ 43 ][ 127 ],
   alphaCSR[ 43 ][ 128 ],
   alphaCSR[ 43 ][ 129 ],
   alphaCSR[ 43 ][ 130 ],
   alphaCSR[ 43 ][ 131 ],
   alphaCSR[ 43 ][ 132 ],
   alphaCSR[ 43 ][ 133 ],
   alphaCSR[ 43 ][ 134 ],
   alphaCSR[ 43 ][ 135 ],
   alphaCSR[ 43 ][ 136 ],
   alphaCSR[ 43 ][ 137 ],
   alphaCSR[ 43 ][ 138 ],
   alphaCSR[ 43 ][ 139 ],
   alphaCSR[ 43 ][ 140 ],
   alphaCSR[ 43 ][ 141 ],
   alphaCSR[ 43 ][ 142 ],
   alphaCSR[ 43 ][ 143 ],
   alphaCSR[ 43 ][ 144 ],
   alphaCSR[ 43 ][ 145 ],
   alphaCSR[ 43 ][ 146 ],
   alphaCSR[ 43 ][ 147 ],
   alphaCSR[ 43 ][ 148 ],
   alphaCSR[ 43 ][ 149 ],
   alphaCSR[ 43 ][ 150 ],
   alphaCSR[ 43 ][ 151 ],
   alphaCSR[ 43 ][ 152 ],
   alphaCSR[ 43 ][ 153 ],
   alphaCSR[ 43 ][ 154 ],
   alphaCSR[ 43 ][ 155 ],
   alphaCSR[ 43 ][ 156 ],
   alphaCSR[ 43 ][ 157 ],
   alphaCSR[ 43 ][ 158 ],
   alphaCSR[ 43 ][ 159 ],
   alphaCSR[ 43 ][ 160 ],
   alphaCSR[ 43 ][ 161 ],
   alphaCSR[ 43 ][ 162 ],
   alphaCSR[ 43 ][ 163 ],
   alphaCSR[ 43 ][ 164 ],
   alphaCSR[ 43 ][ 165 ],
   alphaCSR[ 43 ][ 166 ],
   alphaCSR[ 43 ][ 167 ],
   alphaCSR[ 43 ][ 168 ],
   alphaCSR[ 43 ][ 169 ],
   alphaCSR[ 43 ][ 170 ],
   alphaCSR[ 43 ][ 171 ],
   alphaCSR[ 43 ][ 172 ],
   alphaCSR[ 43 ][ 173 ],
   alphaCSR[ 43 ][ 174 ],
   alphaCSR[ 43 ][ 175 ],
   alphaCSR[ 43 ][ 176 ],
   alphaCSR[ 43 ][ 177 ],
   alphaCSR[ 43 ][ 178 ],
   alphaCSR[ 43 ][ 179 ],
   alphaCSR[ 43 ][ 180 ],
   alphaCSR[ 43 ][ 181 ],
   alphaCSR[ 43 ][ 182 ],
   alphaCSR[ 43 ][ 183 ],
   alphaCSR[ 43 ][ 184 ],
   alphaCSR[ 43 ][ 185 ],
   alphaCSR[ 43 ][ 186 ],
   alphaCSR[ 43 ][ 187 ],
   alphaCSR[ 43 ][ 188 ],
   alphaCSR[ 43 ][ 189 ],
   alphaCSR[ 43 ][ 190 ],
   alphaCSR[ 43 ][ 191 ],
   alphaCSR[ 43 ][ 192 ],
   alphaCSR[ 43 ][ 193 ],
   alphaCSR[ 43 ][ 194 ],
   alphaCSR[ 43 ][ 195 ],
   alphaCSR[ 43 ][ 196 ],
   alphaCSR[ 43 ][ 197 ],
   alphaCSR[ 43 ][ 198 ],
   alphaCSR[ 43 ][ 199 ],
   alphaCSR[ 43 ][ 200 ],
   alphaCSR[ 43 ][ 201 ],
   alphaCSR[ 43 ][ 202 ],
   alphaCSR[ 43 ][ 203 ],
   alphaCSR[ 43 ][ 204 ],
   alphaCSR[ 43 ][ 205 ],
   alphaCSR[ 43 ][ 206 ],
   alphaCSR[ 43 ][ 207 ],
   alphaCSR[ 43 ][ 208 ],
   alphaCSR[ 43 ][ 209 ],
   alphaCSR[ 43 ][ 210 ],
   alphaCSR[ 43 ][ 211 ],
   alphaCSR[ 43 ][ 212 ],
   alphaCSR[ 43 ][ 213 ],
   alphaCSR[ 43 ][ 214 ],
   alphaCSR[ 43 ][ 215 ],
   alphaCSR[ 43 ][ 216 ],
   alphaCSR[ 43 ][ 217 ],
   alphaCSR[ 43 ][ 218 ],
   alphaCSR[ 43 ][ 219 ],
   alphaCSR[ 43 ][ 220 ],
   alphaCSR[ 43 ][ 221 ],
   alphaCSR[ 43 ][ 222 ],
   alphaCSR[ 43 ][ 223 ],
   alphaCSR[ 43 ][ 224 ],
   alphaCSR[ 43 ][ 225 ],
   alphaCSR[ 43 ][ 226 ],
   alphaCSR[ 43 ][ 227 ],
   alphaCSR[ 43 ][ 228 ],
   alphaCSR[ 43 ][ 229 ],
   alphaCSR[ 43 ][ 230 ],
   alphaCSR[ 43 ][ 231 ],
   alphaCSR[ 43 ][ 232 ],
   alphaCSR[ 43 ][ 233 ],
   alphaCSR[ 43 ][ 234 ],
   alphaCSR[ 43 ][ 235 ],
   alphaCSR[ 43 ][ 236 ],
   alphaCSR[ 43 ][ 237 ],
   alphaCSR[ 43 ][ 238 ],
   alphaCSR[ 43 ][ 239 ],
   alphaCSR[ 43 ][ 240 ],
   alphaCSR[ 43 ][ 241 ],
   alphaCSR[ 43 ][ 242 ],
   alphaCSR[ 43 ][ 243 ],
   alphaCSR[ 43 ][ 244 ],
   alphaCSR[ 43 ][ 245 ],
   alphaCSR[ 43 ][ 246 ],
   alphaCSR[ 43 ][ 247 ],
   alphaCSR[ 43 ][ 248 ],
   alphaCSR[ 43 ][ 249 ],
   alphaCSR[ 43 ][ 250 ],
   alphaCSR[ 43 ][ 251 ],
   alphaCSR[ 43 ][ 252 ],
   alphaCSR[ 43 ][ 253 ],
   alphaCSR[ 43 ][ 254 ],
   alphaCSR[ 43 ][ 255 ],
   alphaCSR[ 43 ][ 256 ],
   alphaCSR[ 43 ][ 257 ],
   alphaCSR[ 43 ][ 258 ],
   alphaCSR[ 43 ][ 259 ],
   alphaCSR[ 43 ][ 260 ],
   alphaCSR[ 43 ][ 261 ],
   alphaCSR[ 43 ][ 262 ],
   alphaCSR[ 43 ][ 263 ],
   alphaCSR[ 43 ][ 264 ],
   alphaCSR[ 43 ][ 265 ],
   alphaCSR[ 43 ][ 266 ],
   alphaCSR[ 43 ][ 267 ],
   alphaCSR[ 43 ][ 268 ],
   alphaCSR[ 43 ][ 269 ],
   alphaCSR[ 43 ][ 270 ],
   alphaCSR[ 43 ][ 271 ],
   alphaCSR[ 43 ][ 272 ],
   alphaCSR[ 43 ][ 273 ],
   alphaCSR[ 43 ][ 274 ],
   alphaCSR[ 43 ][ 275 ],
   alphaCSR[ 43 ][ 276 ],
   alphaCSR[ 43 ][ 277 ],
   alphaCSR[ 43 ][ 278 ],
   alphaCSR[ 43 ][ 279 ],
   alphaCSR[ 43 ][ 280 ],
   alphaCSR[ 43 ][ 281 ],
   alphaCSR[ 43 ][ 282 ],
   alphaCSR[ 43 ][ 283 ],
   alphaCSR[ 43 ][ 284 ],
   alphaCSR[ 43 ][ 285 ],
   alphaCSR[ 43 ][ 286 ],
   alphaCSR[ 43 ][ 287 ],
   alphaCSR[ 43 ][ 288 ],
   alphaCSR[ 43 ][ 289 ],
   alphaCSR[ 43 ][ 290 ],
   alphaCSR[ 43 ][ 291 ],
   alphaCSR[ 43 ][ 292 ],
   alphaCSR[ 43 ][ 293 ],
   alphaCSR[ 43 ][ 294 ],
   alphaCSR[ 43 ][ 295 ],
   alphaCSR[ 43 ][ 296 ],
   alphaCSR[ 43 ][ 297 ],
   alphaCSR[ 43 ][ 298 ],
   alphaCSR[ 43 ][ 299 ],
   alphaCSR[ 43 ][ 300 ],
   alphaCSR[ 43 ][ 301 ],
   alphaCSR[ 43 ][ 302 ],
   alphaCSR[ 43 ][ 303 ],
   alphaCSR[ 43 ][ 304 ],
   alphaCSR[ 43 ][ 305 ],
   alphaCSR[ 43 ][ 306 ],
   alphaCSR[ 43 ][ 307 ],
   alphaCSR[ 43 ][ 308 ],
   alphaCSR[ 43 ][ 309 ],
   alphaCSR[ 43 ][ 310 ],
   alphaCSR[ 43 ][ 311 ],
   alphaCSR[ 43 ][ 312 ],
   alphaCSR[ 43 ][ 313 ],
   alphaCSR[ 43 ][ 314 ],
   alphaCSR[ 43 ][ 315 ],
   alphaCSR[ 43 ][ 316 ],
   alphaCSR[ 43 ][ 317 ],
   alphaCSR[ 43 ][ 318 ],
   alphaCSR[ 43 ][ 319 ],
   alphaCSR[ 43 ][ 320 ],
   alphaCSR[ 43 ][ 321 ],
   alphaCSR[ 43 ][ 322 ],
   alphaCSR[ 43 ][ 323 ],
   alphaCSR[ 43 ][ 324 ],
   alphaCSR[ 43 ][ 325 ],
   alphaCSR[ 43 ][ 326 ],
   alphaCSR[ 43 ][ 327 ],
   alphaCSR[ 43 ][ 328 ],
   alphaCSR[ 43 ][ 329 ],
   alphaCSR[ 43 ][ 330 ],
   alphaCSR[ 43 ][ 331 ],
   alphaCSR[ 43 ][ 332 ],
   alphaCSR[ 43 ][ 333 ],
   alphaCSR[ 43 ][ 334 ],
   alphaCSR[ 43 ][ 335 ],
   alphaCSR[ 43 ][ 336 ],
   alphaCSR[ 43 ][ 337 ],
   alphaCSR[ 43 ][ 338 ],
   alphaCSR[ 43 ][ 339 ],
   alphaCSR[ 43 ][ 340 ],
   alphaCSR[ 43 ][ 341 ],
   alphaCSR[ 43 ][ 342 ],
   alphaCSR[ 43 ][ 343 ],
   alphaCSR[ 43 ][ 344 ],
   alphaCSR[ 43 ][ 345 ],
   alphaCSR[ 43 ][ 346 ],
   alphaCSR[ 43 ][ 347 ],
   alphaCSR[ 43 ][ 348 ],
   alphaCSR[ 43 ][ 349 ],
   alphaCSR[ 43 ][ 350 ],
   alphaCSR[ 43 ][ 351 ],
   alphaCSR[ 43 ][ 352 ],
   alphaCSR[ 43 ][ 353 ],
   alphaCSR[ 43 ][ 354 ],
   alphaCSR[ 43 ][ 355 ],
   alphaCSR[ 43 ][ 356 ],
   alphaCSR[ 43 ][ 357 ],
   alphaCSR[ 43 ][ 358 ],
   alphaCSR[ 43 ][ 359 ],
   alphaCSR[ 43 ][ 360 ],
   alphaCSR[ 43 ][ 361 ],
   alphaCSR[ 43 ][ 362 ],
   alphaCSR[ 43 ][ 363 ],
   alphaCSR[ 43 ][ 364 ],
   alphaCSR[ 43 ][ 365 ],
   alphaCSR[ 43 ][ 366 ],
   alphaCSR[ 43 ][ 367 ],
   alphaCSR[ 43 ][ 368 ],
   alphaCSR[ 43 ][ 369 ],
   alphaCSR[ 43 ][ 370 ],
   alphaCSR[ 43 ][ 371 ],
   alphaCSR[ 43 ][ 372 ],
   alphaCSR[ 43 ][ 373 ],
   alphaCSR[ 43 ][ 374 ],
   alphaCSR[ 43 ][ 375 ],
   alphaCSR[ 43 ][ 376 ],
   alphaCSR[ 43 ][ 377 ],
   alphaCSR[ 43 ][ 378 ],
   alphaCSR[ 43 ][ 379 ],
   alphaCSR[ 43 ][ 380 ],
   alphaCSR[ 43 ][ 381 ],
   alphaCSR[ 43 ][ 382 ],
   alphaCSR[ 43 ][ 383 ],
   alphaCSR[ 44 ][ 0 ],
   alphaCSR[ 44 ][ 1 ],
   alphaCSR[ 44 ][ 2 ],
   alphaCSR[ 44 ][ 3 ],
   alphaCSR[ 44 ][ 4 ],
   alphaCSR[ 44 ][ 5 ],
   alphaCSR[ 44 ][ 6 ],
   alphaCSR[ 44 ][ 7 ],
   alphaCSR[ 44 ][ 8 ],
   alphaCSR[ 44 ][ 9 ],
   alphaCSR[ 44 ][ 10 ],
   alphaCSR[ 44 ][ 11 ],
   alphaCSR[ 44 ][ 12 ],
   alphaCSR[ 44 ][ 13 ],
   alphaCSR[ 44 ][ 14 ],
   alphaCSR[ 44 ][ 15 ],
   alphaCSR[ 44 ][ 16 ],
   alphaCSR[ 44 ][ 17 ],
   alphaCSR[ 44 ][ 18 ],
   alphaCSR[ 44 ][ 19 ],
   alphaCSR[ 44 ][ 20 ],
   alphaCSR[ 44 ][ 21 ],
   alphaCSR[ 44 ][ 22 ],
   alphaCSR[ 44 ][ 23 ],
   alphaCSR[ 44 ][ 24 ],
   alphaCSR[ 44 ][ 25 ],
   alphaCSR[ 44 ][ 26 ],
   alphaCSR[ 44 ][ 27 ],
   alphaCSR[ 44 ][ 28 ],
   alphaCSR[ 44 ][ 29 ],
   alphaCSR[ 44 ][ 30 ],
   alphaCSR[ 44 ][ 31 ],
   alphaCSR[ 44 ][ 32 ],
   alphaCSR[ 44 ][ 33 ],
   alphaCSR[ 44 ][ 34 ],
   alphaCSR[ 44 ][ 35 ],
   alphaCSR[ 44 ][ 36 ],
   alphaCSR[ 44 ][ 37 ],
   alphaCSR[ 44 ][ 38 ],
   alphaCSR[ 44 ][ 39 ],
   alphaCSR[ 44 ][ 40 ],
   alphaCSR[ 44 ][ 41 ],
   alphaCSR[ 44 ][ 42 ],
   alphaCSR[ 44 ][ 43 ],
   alphaCSR[ 44 ][ 44 ],
   alphaCSR[ 44 ][ 45 ],
   alphaCSR[ 44 ][ 46 ],
   alphaCSR[ 44 ][ 47 ],
   alphaCSR[ 44 ][ 48 ],
   alphaCSR[ 44 ][ 49 ],
   alphaCSR[ 44 ][ 50 ],
   alphaCSR[ 44 ][ 51 ],
   alphaCSR[ 44 ][ 52 ],
   alphaCSR[ 44 ][ 53 ],
   alphaCSR[ 44 ][ 54 ],
   alphaCSR[ 44 ][ 55 ],
   alphaCSR[ 44 ][ 56 ],
   alphaCSR[ 44 ][ 57 ],
   alphaCSR[ 44 ][ 58 ],
   alphaCSR[ 44 ][ 59 ],
   alphaCSR[ 44 ][ 60 ],
   alphaCSR[ 44 ][ 61 ],
   alphaCSR[ 44 ][ 62 ],
   alphaCSR[ 44 ][ 63 ],
   alphaCSR[ 44 ][ 64 ],
   alphaCSR[ 44 ][ 65 ],
   alphaCSR[ 44 ][ 66 ],
   alphaCSR[ 44 ][ 67 ],
   alphaCSR[ 44 ][ 68 ],
   alphaCSR[ 44 ][ 69 ],
   alphaCSR[ 44 ][ 70 ],
   alphaCSR[ 44 ][ 71 ],
   alphaCSR[ 44 ][ 72 ],
   alphaCSR[ 44 ][ 73 ],
   alphaCSR[ 44 ][ 74 ],
   alphaCSR[ 44 ][ 75 ],
   alphaCSR[ 44 ][ 76 ],
   alphaCSR[ 44 ][ 77 ],
   alphaCSR[ 44 ][ 78 ],
   alphaCSR[ 44 ][ 79 ],
   alphaCSR[ 44 ][ 80 ],
   alphaCSR[ 44 ][ 81 ],
   alphaCSR[ 44 ][ 82 ],
   alphaCSR[ 44 ][ 83 ],
   alphaCSR[ 44 ][ 84 ],
   alphaCSR[ 44 ][ 85 ],
   alphaCSR[ 44 ][ 86 ],
   alphaCSR[ 44 ][ 87 ],
   alphaCSR[ 44 ][ 88 ],
   alphaCSR[ 44 ][ 89 ],
   alphaCSR[ 44 ][ 90 ],
   alphaCSR[ 44 ][ 91 ],
   alphaCSR[ 44 ][ 92 ],
   alphaCSR[ 44 ][ 93 ],
   alphaCSR[ 44 ][ 94 ],
   alphaCSR[ 44 ][ 95 ],
   alphaCSR[ 44 ][ 96 ],
   alphaCSR[ 44 ][ 97 ],
   alphaCSR[ 44 ][ 98 ],
   alphaCSR[ 44 ][ 99 ],
   alphaCSR[ 44 ][ 100 ],
   alphaCSR[ 44 ][ 101 ],
   alphaCSR[ 44 ][ 102 ],
   alphaCSR[ 44 ][ 103 ],
   alphaCSR[ 44 ][ 104 ],
   alphaCSR[ 44 ][ 105 ],
   alphaCSR[ 44 ][ 106 ],
   alphaCSR[ 44 ][ 107 ],
   alphaCSR[ 44 ][ 108 ],
   alphaCSR[ 44 ][ 109 ],
   alphaCSR[ 44 ][ 110 ],
   alphaCSR[ 44 ][ 111 ],
   alphaCSR[ 44 ][ 112 ],
   alphaCSR[ 44 ][ 113 ],
   alphaCSR[ 44 ][ 114 ],
   alphaCSR[ 44 ][ 115 ],
   alphaCSR[ 44 ][ 116 ],
   alphaCSR[ 44 ][ 117 ],
   alphaCSR[ 44 ][ 118 ],
   alphaCSR[ 44 ][ 119 ],
   alphaCSR[ 44 ][ 120 ],
   alphaCSR[ 44 ][ 121 ],
   alphaCSR[ 44 ][ 122 ],
   alphaCSR[ 44 ][ 123 ],
   alphaCSR[ 44 ][ 124 ],
   alphaCSR[ 44 ][ 125 ],
   alphaCSR[ 44 ][ 126 ],
   alphaCSR[ 44 ][ 127 ],
   alphaCSR[ 44 ][ 128 ],
   alphaCSR[ 44 ][ 129 ],
   alphaCSR[ 44 ][ 130 ],
   alphaCSR[ 44 ][ 131 ],
   alphaCSR[ 44 ][ 132 ],
   alphaCSR[ 44 ][ 133 ],
   alphaCSR[ 44 ][ 134 ],
   alphaCSR[ 44 ][ 135 ],
   alphaCSR[ 44 ][ 136 ],
   alphaCSR[ 44 ][ 137 ],
   alphaCSR[ 44 ][ 138 ],
   alphaCSR[ 44 ][ 139 ],
   alphaCSR[ 44 ][ 140 ],
   alphaCSR[ 44 ][ 141 ],
   alphaCSR[ 44 ][ 142 ],
   alphaCSR[ 44 ][ 143 ],
   alphaCSR[ 44 ][ 144 ],
   alphaCSR[ 44 ][ 145 ],
   alphaCSR[ 44 ][ 146 ],
   alphaCSR[ 44 ][ 147 ],
   alphaCSR[ 44 ][ 148 ],
   alphaCSR[ 44 ][ 149 ],
   alphaCSR[ 44 ][ 150 ],
   alphaCSR[ 44 ][ 151 ],
   alphaCSR[ 44 ][ 152 ],
   alphaCSR[ 44 ][ 153 ],
   alphaCSR[ 44 ][ 154 ],
   alphaCSR[ 44 ][ 155 ],
   alphaCSR[ 44 ][ 156 ],
   alphaCSR[ 44 ][ 157 ],
   alphaCSR[ 44 ][ 158 ],
   alphaCSR[ 44 ][ 159 ],
   alphaCSR[ 44 ][ 160 ],
   alphaCSR[ 44 ][ 161 ],
   alphaCSR[ 44 ][ 162 ],
   alphaCSR[ 44 ][ 163 ],
   alphaCSR[ 44 ][ 164 ],
   alphaCSR[ 44 ][ 165 ],
   alphaCSR[ 44 ][ 166 ],
   alphaCSR[ 44 ][ 167 ],
   alphaCSR[ 44 ][ 168 ],
   alphaCSR[ 44 ][ 169 ],
   alphaCSR[ 44 ][ 170 ],
   alphaCSR[ 44 ][ 171 ],
   alphaCSR[ 44 ][ 172 ],
   alphaCSR[ 44 ][ 173 ],
   alphaCSR[ 44 ][ 174 ],
   alphaCSR[ 44 ][ 175 ],
   alphaCSR[ 44 ][ 176 ],
   alphaCSR[ 44 ][ 177 ],
   alphaCSR[ 44 ][ 178 ],
   alphaCSR[ 44 ][ 179 ],
   alphaCSR[ 44 ][ 180 ],
   alphaCSR[ 44 ][ 181 ],
   alphaCSR[ 44 ][ 182 ],
   alphaCSR[ 44 ][ 183 ],
   alphaCSR[ 44 ][ 184 ],
   alphaCSR[ 44 ][ 185 ],
   alphaCSR[ 44 ][ 186 ],
   alphaCSR[ 44 ][ 187 ],
   alphaCSR[ 44 ][ 188 ],
   alphaCSR[ 44 ][ 189 ],
   alphaCSR[ 44 ][ 190 ],
   alphaCSR[ 44 ][ 191 ],
   alphaCSR[ 44 ][ 192 ],
   alphaCSR[ 44 ][ 193 ],
   alphaCSR[ 44 ][ 194 ],
   alphaCSR[ 44 ][ 195 ],
   alphaCSR[ 44 ][ 196 ],
   alphaCSR[ 44 ][ 197 ],
   alphaCSR[ 44 ][ 198 ],
   alphaCSR[ 44 ][ 199 ],
   alphaCSR[ 44 ][ 200 ],
   alphaCSR[ 44 ][ 201 ],
   alphaCSR[ 44 ][ 202 ],
   alphaCSR[ 44 ][ 203 ],
   alphaCSR[ 44 ][ 204 ],
   alphaCSR[ 44 ][ 205 ],
   alphaCSR[ 44 ][ 206 ],
   alphaCSR[ 44 ][ 207 ],
   alphaCSR[ 44 ][ 208 ],
   alphaCSR[ 44 ][ 209 ],
   alphaCSR[ 44 ][ 210 ],
   alphaCSR[ 44 ][ 211 ],
   alphaCSR[ 44 ][ 212 ],
   alphaCSR[ 44 ][ 213 ],
   alphaCSR[ 44 ][ 214 ],
   alphaCSR[ 44 ][ 215 ],
   alphaCSR[ 44 ][ 216 ],
   alphaCSR[ 44 ][ 217 ],
   alphaCSR[ 44 ][ 218 ],
   alphaCSR[ 44 ][ 219 ],
   alphaCSR[ 44 ][ 220 ],
   alphaCSR[ 44 ][ 221 ],
   alphaCSR[ 44 ][ 222 ],
   alphaCSR[ 44 ][ 223 ],
   alphaCSR[ 44 ][ 224 ],
   alphaCSR[ 44 ][ 225 ],
   alphaCSR[ 44 ][ 226 ],
   alphaCSR[ 44 ][ 227 ],
   alphaCSR[ 44 ][ 228 ],
   alphaCSR[ 44 ][ 229 ],
   alphaCSR[ 44 ][ 230 ],
   alphaCSR[ 44 ][ 231 ],
   alphaCSR[ 44 ][ 232 ],
   alphaCSR[ 44 ][ 233 ],
   alphaCSR[ 44 ][ 234 ],
   alphaCSR[ 44 ][ 235 ],
   alphaCSR[ 44 ][ 236 ],
   alphaCSR[ 44 ][ 237 ],
   alphaCSR[ 44 ][ 238 ],
   alphaCSR[ 44 ][ 239 ],
   alphaCSR[ 44 ][ 240 ],
   alphaCSR[ 44 ][ 241 ],
   alphaCSR[ 44 ][ 242 ],
   alphaCSR[ 44 ][ 243 ],
   alphaCSR[ 44 ][ 244 ],
   alphaCSR[ 44 ][ 245 ],
   alphaCSR[ 44 ][ 246 ],
   alphaCSR[ 44 ][ 247 ],
   alphaCSR[ 44 ][ 248 ],
   alphaCSR[ 44 ][ 249 ],
   alphaCSR[ 44 ][ 250 ],
   alphaCSR[ 44 ][ 251 ],
   alphaCSR[ 44 ][ 252 ],
   alphaCSR[ 44 ][ 253 ],
   alphaCSR[ 44 ][ 254 ],
   alphaCSR[ 44 ][ 255 ],
   alphaCSR[ 44 ][ 256 ],
   alphaCSR[ 44 ][ 257 ],
   alphaCSR[ 44 ][ 258 ],
   alphaCSR[ 44 ][ 259 ],
   alphaCSR[ 44 ][ 260 ],
   alphaCSR[ 44 ][ 261 ],
   alphaCSR[ 44 ][ 262 ],
   alphaCSR[ 44 ][ 263 ],
   alphaCSR[ 44 ][ 264 ],
   alphaCSR[ 44 ][ 265 ],
   alphaCSR[ 44 ][ 266 ],
   alphaCSR[ 44 ][ 267 ],
   alphaCSR[ 44 ][ 268 ],
   alphaCSR[ 44 ][ 269 ],
   alphaCSR[ 44 ][ 270 ],
   alphaCSR[ 44 ][ 271 ],
   alphaCSR[ 44 ][ 272 ],
   alphaCSR[ 44 ][ 273 ],
   alphaCSR[ 44 ][ 274 ],
   alphaCSR[ 44 ][ 275 ],
   alphaCSR[ 44 ][ 276 ],
   alphaCSR[ 44 ][ 277 ],
   alphaCSR[ 44 ][ 278 ],
   alphaCSR[ 44 ][ 279 ],
   alphaCSR[ 44 ][ 280 ],
   alphaCSR[ 44 ][ 281 ],
   alphaCSR[ 44 ][ 282 ],
   alphaCSR[ 44 ][ 283 ],
   alphaCSR[ 44 ][ 284 ],
   alphaCSR[ 44 ][ 285 ],
   alphaCSR[ 44 ][ 286 ],
   alphaCSR[ 44 ][ 287 ],
   alphaCSR[ 44 ][ 288 ],
   alphaCSR[ 44 ][ 289 ],
   alphaCSR[ 44 ][ 290 ],
   alphaCSR[ 44 ][ 291 ],
   alphaCSR[ 44 ][ 292 ],
   alphaCSR[ 44 ][ 293 ],
   alphaCSR[ 44 ][ 294 ],
   alphaCSR[ 44 ][ 295 ],
   alphaCSR[ 44 ][ 296 ],
   alphaCSR[ 44 ][ 297 ],
   alphaCSR[ 44 ][ 298 ],
   alphaCSR[ 44 ][ 299 ],
   alphaCSR[ 44 ][ 300 ],
   alphaCSR[ 44 ][ 301 ],
   alphaCSR[ 44 ][ 302 ],
   alphaCSR[ 44 ][ 303 ],
   alphaCSR[ 44 ][ 304 ],
   alphaCSR[ 44 ][ 305 ],
   alphaCSR[ 44 ][ 306 ],
   alphaCSR[ 44 ][ 307 ],
   alphaCSR[ 44 ][ 308 ],
   alphaCSR[ 44 ][ 309 ],
   alphaCSR[ 44 ][ 310 ],
   alphaCSR[ 44 ][ 311 ],
   alphaCSR[ 44 ][ 312 ],
   alphaCSR[ 44 ][ 313 ],
   alphaCSR[ 44 ][ 314 ],
   alphaCSR[ 44 ][ 315 ],
   alphaCSR[ 44 ][ 316 ],
   alphaCSR[ 44 ][ 317 ],
   alphaCSR[ 44 ][ 318 ],
   alphaCSR[ 44 ][ 319 ],
   alphaCSR[ 44 ][ 320 ],
   alphaCSR[ 44 ][ 321 ],
   alphaCSR[ 44 ][ 322 ],
   alphaCSR[ 44 ][ 323 ],
   alphaCSR[ 44 ][ 324 ],
   alphaCSR[ 44 ][ 325 ],
   alphaCSR[ 44 ][ 326 ],
   alphaCSR[ 44 ][ 327 ],
   alphaCSR[ 44 ][ 328 ],
   alphaCSR[ 44 ][ 329 ],
   alphaCSR[ 44 ][ 330 ],
   alphaCSR[ 44 ][ 331 ],
   alphaCSR[ 44 ][ 332 ],
   alphaCSR[ 44 ][ 333 ],
   alphaCSR[ 44 ][ 334 ],
   alphaCSR[ 44 ][ 335 ],
   alphaCSR[ 44 ][ 336 ],
   alphaCSR[ 44 ][ 337 ],
   alphaCSR[ 44 ][ 338 ],
   alphaCSR[ 44 ][ 339 ],
   alphaCSR[ 44 ][ 340 ],
   alphaCSR[ 44 ][ 341 ],
   alphaCSR[ 44 ][ 342 ],
   alphaCSR[ 44 ][ 343 ],
   alphaCSR[ 44 ][ 344 ],
   alphaCSR[ 44 ][ 345 ],
   alphaCSR[ 44 ][ 346 ],
   alphaCSR[ 44 ][ 347 ],
   alphaCSR[ 44 ][ 348 ],
   alphaCSR[ 44 ][ 349 ],
   alphaCSR[ 44 ][ 350 ],
   alphaCSR[ 44 ][ 351 ],
   alphaCSR[ 44 ][ 352 ],
   alphaCSR[ 44 ][ 353 ],
   alphaCSR[ 44 ][ 354 ],
   alphaCSR[ 44 ][ 355 ],
   alphaCSR[ 44 ][ 356 ],
   alphaCSR[ 44 ][ 357 ],
   alphaCSR[ 44 ][ 358 ],
   alphaCSR[ 44 ][ 359 ],
   alphaCSR[ 44 ][ 360 ],
   alphaCSR[ 44 ][ 361 ],
   alphaCSR[ 44 ][ 362 ],
   alphaCSR[ 44 ][ 363 ],
   alphaCSR[ 44 ][ 364 ],
   alphaCSR[ 44 ][ 365 ],
   alphaCSR[ 44 ][ 366 ],
   alphaCSR[ 44 ][ 367 ],
   alphaCSR[ 44 ][ 368 ],
   alphaCSR[ 44 ][ 369 ],
   alphaCSR[ 44 ][ 370 ],
   alphaCSR[ 44 ][ 371 ],
   alphaCSR[ 44 ][ 372 ],
   alphaCSR[ 44 ][ 373 ],
   alphaCSR[ 44 ][ 374 ],
   alphaCSR[ 44 ][ 375 ],
   alphaCSR[ 44 ][ 376 ],
   alphaCSR[ 44 ][ 377 ],
   alphaCSR[ 44 ][ 378 ],
   alphaCSR[ 44 ][ 379 ],
   alphaCSR[ 44 ][ 380 ],
   alphaCSR[ 44 ][ 381 ],
   alphaCSR[ 44 ][ 382 ],
   alphaCSR[ 44 ][ 383 ],
   alphaCSR[ 45 ][ 0 ],
   alphaCSR[ 45 ][ 1 ],
   alphaCSR[ 45 ][ 2 ],
   alphaCSR[ 45 ][ 3 ],
   alphaCSR[ 45 ][ 4 ],
   alphaCSR[ 45 ][ 5 ],
   alphaCSR[ 45 ][ 6 ],
   alphaCSR[ 45 ][ 7 ],
   alphaCSR[ 45 ][ 8 ],
   alphaCSR[ 45 ][ 9 ],
   alphaCSR[ 45 ][ 10 ],
   alphaCSR[ 45 ][ 11 ],
   alphaCSR[ 45 ][ 12 ],
   alphaCSR[ 45 ][ 13 ],
   alphaCSR[ 45 ][ 14 ],
   alphaCSR[ 45 ][ 15 ],
   alphaCSR[ 45 ][ 16 ],
   alphaCSR[ 45 ][ 17 ],
   alphaCSR[ 45 ][ 18 ],
   alphaCSR[ 45 ][ 19 ],
   alphaCSR[ 45 ][ 20 ],
   alphaCSR[ 45 ][ 21 ],
   alphaCSR[ 45 ][ 22 ],
   alphaCSR[ 45 ][ 23 ],
   alphaCSR[ 45 ][ 24 ],
   alphaCSR[ 45 ][ 25 ],
   alphaCSR[ 45 ][ 26 ],
   alphaCSR[ 45 ][ 27 ],
   alphaCSR[ 45 ][ 28 ],
   alphaCSR[ 45 ][ 29 ],
   alphaCSR[ 45 ][ 30 ],
   alphaCSR[ 45 ][ 31 ],
   alphaCSR[ 45 ][ 32 ],
   alphaCSR[ 45 ][ 33 ],
   alphaCSR[ 45 ][ 34 ],
   alphaCSR[ 45 ][ 35 ],
   alphaCSR[ 45 ][ 36 ],
   alphaCSR[ 45 ][ 37 ],
   alphaCSR[ 45 ][ 38 ],
   alphaCSR[ 45 ][ 39 ],
   alphaCSR[ 45 ][ 40 ],
   alphaCSR[ 45 ][ 41 ],
   alphaCSR[ 45 ][ 42 ],
   alphaCSR[ 45 ][ 43 ],
   alphaCSR[ 45 ][ 44 ],
   alphaCSR[ 45 ][ 45 ],
   alphaCSR[ 45 ][ 46 ],
   alphaCSR[ 45 ][ 47 ],
   alphaCSR[ 45 ][ 48 ],
   alphaCSR[ 45 ][ 49 ],
   alphaCSR[ 45 ][ 50 ],
   alphaCSR[ 45 ][ 51 ],
   alphaCSR[ 45 ][ 52 ],
   alphaCSR[ 45 ][ 53 ],
   alphaCSR[ 45 ][ 54 ],
   alphaCSR[ 45 ][ 55 ],
   alphaCSR[ 45 ][ 56 ],
   alphaCSR[ 45 ][ 57 ],
   alphaCSR[ 45 ][ 58 ],
   alphaCSR[ 45 ][ 59 ],
   alphaCSR[ 45 ][ 60 ],
   alphaCSR[ 45 ][ 61 ],
   alphaCSR[ 45 ][ 62 ],
   alphaCSR[ 45 ][ 63 ],
   alphaCSR[ 45 ][ 64 ],
   alphaCSR[ 45 ][ 65 ],
   alphaCSR[ 45 ][ 66 ],
   alphaCSR[ 45 ][ 67 ],
   alphaCSR[ 45 ][ 68 ],
   alphaCSR[ 45 ][ 69 ],
   alphaCSR[ 45 ][ 70 ],
   alphaCSR[ 45 ][ 71 ],
   alphaCSR[ 45 ][ 72 ],
   alphaCSR[ 45 ][ 73 ],
   alphaCSR[ 45 ][ 74 ],
   alphaCSR[ 45 ][ 75 ],
   alphaCSR[ 45 ][ 76 ],
   alphaCSR[ 45 ][ 77 ],
   alphaCSR[ 45 ][ 78 ],
   alphaCSR[ 45 ][ 79 ],
   alphaCSR[ 45 ][ 80 ],
   alphaCSR[ 45 ][ 81 ],
   alphaCSR[ 45 ][ 82 ],
   alphaCSR[ 45 ][ 83 ],
   alphaCSR[ 45 ][ 84 ],
   alphaCSR[ 45 ][ 85 ],
   alphaCSR[ 45 ][ 86 ],
   alphaCSR[ 45 ][ 87 ],
   alphaCSR[ 45 ][ 88 ],
   alphaCSR[ 45 ][ 89 ],
   alphaCSR[ 45 ][ 90 ],
   alphaCSR[ 45 ][ 91 ],
   alphaCSR[ 45 ][ 92 ],
   alphaCSR[ 45 ][ 93 ],
   alphaCSR[ 45 ][ 94 ],
   alphaCSR[ 45 ][ 95 ],
   alphaCSR[ 45 ][ 96 ],
   alphaCSR[ 45 ][ 97 ],
   alphaCSR[ 45 ][ 98 ],
   alphaCSR[ 45 ][ 99 ],
   alphaCSR[ 45 ][ 100 ],
   alphaCSR[ 45 ][ 101 ],
   alphaCSR[ 45 ][ 102 ],
   alphaCSR[ 45 ][ 103 ],
   alphaCSR[ 45 ][ 104 ],
   alphaCSR[ 45 ][ 105 ],
   alphaCSR[ 45 ][ 106 ],
   alphaCSR[ 45 ][ 107 ],
   alphaCSR[ 45 ][ 108 ],
   alphaCSR[ 45 ][ 109 ],
   alphaCSR[ 45 ][ 110 ],
   alphaCSR[ 45 ][ 111 ],
   alphaCSR[ 45 ][ 112 ],
   alphaCSR[ 45 ][ 113 ],
   alphaCSR[ 45 ][ 114 ],
   alphaCSR[ 45 ][ 115 ],
   alphaCSR[ 45 ][ 116 ],
   alphaCSR[ 45 ][ 117 ],
   alphaCSR[ 45 ][ 118 ],
   alphaCSR[ 45 ][ 119 ],
   alphaCSR[ 45 ][ 120 ],
   alphaCSR[ 45 ][ 121 ],
   alphaCSR[ 45 ][ 122 ],
   alphaCSR[ 45 ][ 123 ],
   alphaCSR[ 45 ][ 124 ],
   alphaCSR[ 45 ][ 125 ],
   alphaCSR[ 45 ][ 126 ],
   alphaCSR[ 45 ][ 127 ],
   alphaCSR[ 45 ][ 128 ],
   alphaCSR[ 45 ][ 129 ],
   alphaCSR[ 45 ][ 130 ],
   alphaCSR[ 45 ][ 131 ],
   alphaCSR[ 45 ][ 132 ],
   alphaCSR[ 45 ][ 133 ],
   alphaCSR[ 45 ][ 134 ],
   alphaCSR[ 45 ][ 135 ],
   alphaCSR[ 45 ][ 136 ],
   alphaCSR[ 45 ][ 137 ],
   alphaCSR[ 45 ][ 138 ],
   alphaCSR[ 45 ][ 139 ],
   alphaCSR[ 45 ][ 140 ],
   alphaCSR[ 45 ][ 141 ],
   alphaCSR[ 45 ][ 142 ],
   alphaCSR[ 45 ][ 143 ],
   alphaCSR[ 45 ][ 144 ],
   alphaCSR[ 45 ][ 145 ],
   alphaCSR[ 45 ][ 146 ],
   alphaCSR[ 45 ][ 147 ],
   alphaCSR[ 45 ][ 148 ],
   alphaCSR[ 45 ][ 149 ],
   alphaCSR[ 45 ][ 150 ],
   alphaCSR[ 45 ][ 151 ],
   alphaCSR[ 45 ][ 152 ],
   alphaCSR[ 45 ][ 153 ],
   alphaCSR[ 45 ][ 154 ],
   alphaCSR[ 45 ][ 155 ],
   alphaCSR[ 45 ][ 156 ],
   alphaCSR[ 45 ][ 157 ],
   alphaCSR[ 45 ][ 158 ],
   alphaCSR[ 45 ][ 159 ],
   alphaCSR[ 45 ][ 160 ],
   alphaCSR[ 45 ][ 161 ],
   alphaCSR[ 45 ][ 162 ],
   alphaCSR[ 45 ][ 163 ],
   alphaCSR[ 45 ][ 164 ],
   alphaCSR[ 45 ][ 165 ],
   alphaCSR[ 45 ][ 166 ],
   alphaCSR[ 45 ][ 167 ],
   alphaCSR[ 45 ][ 168 ],
   alphaCSR[ 45 ][ 169 ],
   alphaCSR[ 45 ][ 170 ],
   alphaCSR[ 45 ][ 171 ],
   alphaCSR[ 45 ][ 172 ],
   alphaCSR[ 45 ][ 173 ],
   alphaCSR[ 45 ][ 174 ],
   alphaCSR[ 45 ][ 175 ],
   alphaCSR[ 45 ][ 176 ],
   alphaCSR[ 45 ][ 177 ],
   alphaCSR[ 45 ][ 178 ],
   alphaCSR[ 45 ][ 179 ],
   alphaCSR[ 45 ][ 180 ],
   alphaCSR[ 45 ][ 181 ],
   alphaCSR[ 45 ][ 182 ],
   alphaCSR[ 45 ][ 183 ],
   alphaCSR[ 45 ][ 184 ],
   alphaCSR[ 45 ][ 185 ],
   alphaCSR[ 45 ][ 186 ],
   alphaCSR[ 45 ][ 187 ],
   alphaCSR[ 45 ][ 188 ],
   alphaCSR[ 45 ][ 189 ],
   alphaCSR[ 45 ][ 190 ],
   alphaCSR[ 45 ][ 191 ],
   alphaCSR[ 45 ][ 192 ],
   alphaCSR[ 45 ][ 193 ],
   alphaCSR[ 45 ][ 194 ],
   alphaCSR[ 45 ][ 195 ],
   alphaCSR[ 45 ][ 196 ],
   alphaCSR[ 45 ][ 197 ],
   alphaCSR[ 45 ][ 198 ],
   alphaCSR[ 45 ][ 199 ],
   alphaCSR[ 45 ][ 200 ],
   alphaCSR[ 45 ][ 201 ],
   alphaCSR[ 45 ][ 202 ],
   alphaCSR[ 45 ][ 203 ],
   alphaCSR[ 45 ][ 204 ],
   alphaCSR[ 45 ][ 205 ],
   alphaCSR[ 45 ][ 206 ],
   alphaCSR[ 45 ][ 207 ],
   alphaCSR[ 45 ][ 208 ],
   alphaCSR[ 45 ][ 209 ],
   alphaCSR[ 45 ][ 210 ],
   alphaCSR[ 45 ][ 211 ],
   alphaCSR[ 45 ][ 212 ],
   alphaCSR[ 45 ][ 213 ],
   alphaCSR[ 45 ][ 214 ],
   alphaCSR[ 45 ][ 215 ],
   alphaCSR[ 45 ][ 216 ],
   alphaCSR[ 45 ][ 217 ],
   alphaCSR[ 45 ][ 218 ],
   alphaCSR[ 45 ][ 219 ],
   alphaCSR[ 45 ][ 220 ],
   alphaCSR[ 45 ][ 221 ],
   alphaCSR[ 45 ][ 222 ],
   alphaCSR[ 45 ][ 223 ],
   alphaCSR[ 45 ][ 224 ],
   alphaCSR[ 45 ][ 225 ],
   alphaCSR[ 45 ][ 226 ],
   alphaCSR[ 45 ][ 227 ],
   alphaCSR[ 45 ][ 228 ],
   alphaCSR[ 45 ][ 229 ],
   alphaCSR[ 45 ][ 230 ],
   alphaCSR[ 45 ][ 231 ],
   alphaCSR[ 45 ][ 232 ],
   alphaCSR[ 45 ][ 233 ],
   alphaCSR[ 45 ][ 234 ],
   alphaCSR[ 45 ][ 235 ],
   alphaCSR[ 45 ][ 236 ],
   alphaCSR[ 45 ][ 237 ],
   alphaCSR[ 45 ][ 238 ],
   alphaCSR[ 45 ][ 239 ],
   alphaCSR[ 45 ][ 240 ],
   alphaCSR[ 45 ][ 241 ],
   alphaCSR[ 45 ][ 242 ],
   alphaCSR[ 45 ][ 243 ],
   alphaCSR[ 45 ][ 244 ],
   alphaCSR[ 45 ][ 245 ],
   alphaCSR[ 45 ][ 246 ],
   alphaCSR[ 45 ][ 247 ],
   alphaCSR[ 45 ][ 248 ],
   alphaCSR[ 45 ][ 249 ],
   alphaCSR[ 45 ][ 250 ],
   alphaCSR[ 45 ][ 251 ],
   alphaCSR[ 45 ][ 252 ],
   alphaCSR[ 45 ][ 253 ],
   alphaCSR[ 45 ][ 254 ],
   alphaCSR[ 45 ][ 255 ],
   alphaCSR[ 45 ][ 256 ],
   alphaCSR[ 45 ][ 257 ],
   alphaCSR[ 45 ][ 258 ],
   alphaCSR[ 45 ][ 259 ],
   alphaCSR[ 45 ][ 260 ],
   alphaCSR[ 45 ][ 261 ],
   alphaCSR[ 45 ][ 262 ],
   alphaCSR[ 45 ][ 263 ],
   alphaCSR[ 45 ][ 264 ],
   alphaCSR[ 45 ][ 265 ],
   alphaCSR[ 45 ][ 266 ],
   alphaCSR[ 45 ][ 267 ],
   alphaCSR[ 45 ][ 268 ],
   alphaCSR[ 45 ][ 269 ],
   alphaCSR[ 45 ][ 270 ],
   alphaCSR[ 45 ][ 271 ],
   alphaCSR[ 45 ][ 272 ],
   alphaCSR[ 45 ][ 273 ],
   alphaCSR[ 45 ][ 274 ],
   alphaCSR[ 45 ][ 275 ],
   alphaCSR[ 45 ][ 276 ],
   alphaCSR[ 45 ][ 277 ],
   alphaCSR[ 45 ][ 278 ],
   alphaCSR[ 45 ][ 279 ],
   alphaCSR[ 45 ][ 280 ],
   alphaCSR[ 45 ][ 281 ],
   alphaCSR[ 45 ][ 282 ],
   alphaCSR[ 45 ][ 283 ],
   alphaCSR[ 45 ][ 284 ],
   alphaCSR[ 45 ][ 285 ],
   alphaCSR[ 45 ][ 286 ],
   alphaCSR[ 45 ][ 287 ],
   alphaCSR[ 45 ][ 288 ],
   alphaCSR[ 45 ][ 289 ],
   alphaCSR[ 45 ][ 290 ],
   alphaCSR[ 45 ][ 291 ],
   alphaCSR[ 45 ][ 292 ],
   alphaCSR[ 45 ][ 293 ],
   alphaCSR[ 45 ][ 294 ],
   alphaCSR[ 45 ][ 295 ],
   alphaCSR[ 45 ][ 296 ],
   alphaCSR[ 45 ][ 297 ],
   alphaCSR[ 45 ][ 298 ],
   alphaCSR[ 45 ][ 299 ],
   alphaCSR[ 45 ][ 300 ],
   alphaCSR[ 45 ][ 301 ],
   alphaCSR[ 45 ][ 302 ],
   alphaCSR[ 45 ][ 303 ],
   alphaCSR[ 45 ][ 304 ],
   alphaCSR[ 45 ][ 305 ],
   alphaCSR[ 45 ][ 306 ],
   alphaCSR[ 45 ][ 307 ],
   alphaCSR[ 45 ][ 308 ],
   alphaCSR[ 45 ][ 309 ],
   alphaCSR[ 45 ][ 310 ],
   alphaCSR[ 45 ][ 311 ],
   alphaCSR[ 45 ][ 312 ],
   alphaCSR[ 45 ][ 313 ],
   alphaCSR[ 45 ][ 314 ],
   alphaCSR[ 45 ][ 315 ],
   alphaCSR[ 45 ][ 316 ],
   alphaCSR[ 45 ][ 317 ],
   alphaCSR[ 45 ][ 318 ],
   alphaCSR[ 45 ][ 319 ],
   alphaCSR[ 45 ][ 320 ],
   alphaCSR[ 45 ][ 321 ],
   alphaCSR[ 45 ][ 322 ],
   alphaCSR[ 45 ][ 323 ],
   alphaCSR[ 45 ][ 324 ],
   alphaCSR[ 45 ][ 325 ],
   alphaCSR[ 45 ][ 326 ],
   alphaCSR[ 45 ][ 327 ],
   alphaCSR[ 45 ][ 328 ],
   alphaCSR[ 45 ][ 329 ],
   alphaCSR[ 45 ][ 330 ],
   alphaCSR[ 45 ][ 331 ],
   alphaCSR[ 45 ][ 332 ],
   alphaCSR[ 45 ][ 333 ],
   alphaCSR[ 45 ][ 334 ],
   alphaCSR[ 45 ][ 335 ],
   alphaCSR[ 45 ][ 336 ],
   alphaCSR[ 45 ][ 337 ],
   alphaCSR[ 45 ][ 338 ],
   alphaCSR[ 45 ][ 339 ],
   alphaCSR[ 45 ][ 340 ],
   alphaCSR[ 45 ][ 341 ],
   alphaCSR[ 45 ][ 342 ],
   alphaCSR[ 45 ][ 343 ],
   alphaCSR[ 45 ][ 344 ],
   alphaCSR[ 45 ][ 345 ],
   alphaCSR[ 45 ][ 346 ],
   alphaCSR[ 45 ][ 347 ],
   alphaCSR[ 45 ][ 348 ],
   alphaCSR[ 45 ][ 349 ],
   alphaCSR[ 45 ][ 350 ],
   alphaCSR[ 45 ][ 351 ],
   alphaCSR[ 45 ][ 352 ],
   alphaCSR[ 45 ][ 353 ],
   alphaCSR[ 45 ][ 354 ],
   alphaCSR[ 45 ][ 355 ],
   alphaCSR[ 45 ][ 356 ],
   alphaCSR[ 45 ][ 357 ],
   alphaCSR[ 45 ][ 358 ],
   alphaCSR[ 45 ][ 359 ],
   alphaCSR[ 45 ][ 360 ],
   alphaCSR[ 45 ][ 361 ],
   alphaCSR[ 45 ][ 362 ],
   alphaCSR[ 45 ][ 363 ],
   alphaCSR[ 45 ][ 364 ],
   alphaCSR[ 45 ][ 365 ],
   alphaCSR[ 45 ][ 366 ],
   alphaCSR[ 45 ][ 367 ],
   alphaCSR[ 45 ][ 368 ],
   alphaCSR[ 45 ][ 369 ],
   alphaCSR[ 45 ][ 370 ],
   alphaCSR[ 45 ][ 371 ],
   alphaCSR[ 45 ][ 372 ],
   alphaCSR[ 45 ][ 373 ],
   alphaCSR[ 45 ][ 374 ],
   alphaCSR[ 45 ][ 375 ],
   alphaCSR[ 45 ][ 376 ],
   alphaCSR[ 45 ][ 377 ],
   alphaCSR[ 45 ][ 378 ],
   alphaCSR[ 45 ][ 379 ],
   alphaCSR[ 45 ][ 380 ],
   alphaCSR[ 45 ][ 381 ],
   alphaCSR[ 45 ][ 382 ],
   alphaCSR[ 45 ][ 383 ],
   alphaCSR[ 46 ][ 0 ],
   alphaCSR[ 46 ][ 1 ],
   alphaCSR[ 46 ][ 2 ],
   alphaCSR[ 46 ][ 3 ],
   alphaCSR[ 46 ][ 4 ],
   alphaCSR[ 46 ][ 5 ],
   alphaCSR[ 46 ][ 6 ],
   alphaCSR[ 46 ][ 7 ],
   alphaCSR[ 46 ][ 8 ],
   alphaCSR[ 46 ][ 9 ],
   alphaCSR[ 46 ][ 10 ],
   alphaCSR[ 46 ][ 11 ],
   alphaCSR[ 46 ][ 12 ],
   alphaCSR[ 46 ][ 13 ],
   alphaCSR[ 46 ][ 14 ],
   alphaCSR[ 46 ][ 15 ],
   alphaCSR[ 46 ][ 16 ],
   alphaCSR[ 46 ][ 17 ],
   alphaCSR[ 46 ][ 18 ],
   alphaCSR[ 46 ][ 19 ],
   alphaCSR[ 46 ][ 20 ],
   alphaCSR[ 46 ][ 21 ],
   alphaCSR[ 46 ][ 22 ],
   alphaCSR[ 46 ][ 23 ],
   alphaCSR[ 46 ][ 24 ],
   alphaCSR[ 46 ][ 25 ],
   alphaCSR[ 46 ][ 26 ],
   alphaCSR[ 46 ][ 27 ],
   alphaCSR[ 46 ][ 28 ],
   alphaCSR[ 46 ][ 29 ],
   alphaCSR[ 46 ][ 30 ],
   alphaCSR[ 46 ][ 31 ],
   alphaCSR[ 46 ][ 32 ],
   alphaCSR[ 46 ][ 33 ],
   alphaCSR[ 46 ][ 34 ],
   alphaCSR[ 46 ][ 35 ],
   alphaCSR[ 46 ][ 36 ],
   alphaCSR[ 46 ][ 37 ],
   alphaCSR[ 46 ][ 38 ],
   alphaCSR[ 46 ][ 39 ],
   alphaCSR[ 46 ][ 40 ],
   alphaCSR[ 46 ][ 41 ],
   alphaCSR[ 46 ][ 42 ],
   alphaCSR[ 46 ][ 43 ],
   alphaCSR[ 46 ][ 44 ],
   alphaCSR[ 46 ][ 45 ],
   alphaCSR[ 46 ][ 46 ],
   alphaCSR[ 46 ][ 47 ],
   alphaCSR[ 46 ][ 48 ],
   alphaCSR[ 46 ][ 49 ],
   alphaCSR[ 46 ][ 50 ],
   alphaCSR[ 46 ][ 51 ],
   alphaCSR[ 46 ][ 52 ],
   alphaCSR[ 46 ][ 53 ],
   alphaCSR[ 46 ][ 54 ],
   alphaCSR[ 46 ][ 55 ],
   alphaCSR[ 46 ][ 56 ],
   alphaCSR[ 46 ][ 57 ],
   alphaCSR[ 46 ][ 58 ],
   alphaCSR[ 46 ][ 59 ],
   alphaCSR[ 46 ][ 60 ],
   alphaCSR[ 46 ][ 61 ],
   alphaCSR[ 46 ][ 62 ],
   alphaCSR[ 46 ][ 63 ],
   alphaCSR[ 46 ][ 64 ],
   alphaCSR[ 46 ][ 65 ],
   alphaCSR[ 46 ][ 66 ],
   alphaCSR[ 46 ][ 67 ],
   alphaCSR[ 46 ][ 68 ],
   alphaCSR[ 46 ][ 69 ],
   alphaCSR[ 46 ][ 70 ],
   alphaCSR[ 46 ][ 71 ],
   alphaCSR[ 46 ][ 72 ],
   alphaCSR[ 46 ][ 73 ],
   alphaCSR[ 46 ][ 74 ],
   alphaCSR[ 46 ][ 75 ],
   alphaCSR[ 46 ][ 76 ],
   alphaCSR[ 46 ][ 77 ],
   alphaCSR[ 46 ][ 78 ],
   alphaCSR[ 46 ][ 79 ],
   alphaCSR[ 46 ][ 80 ],
   alphaCSR[ 46 ][ 81 ],
   alphaCSR[ 46 ][ 82 ],
   alphaCSR[ 46 ][ 83 ],
   alphaCSR[ 46 ][ 84 ],
   alphaCSR[ 46 ][ 85 ],
   alphaCSR[ 46 ][ 86 ],
   alphaCSR[ 46 ][ 87 ],
   alphaCSR[ 46 ][ 88 ],
   alphaCSR[ 46 ][ 89 ],
   alphaCSR[ 46 ][ 90 ],
   alphaCSR[ 46 ][ 91 ],
   alphaCSR[ 46 ][ 92 ],
   alphaCSR[ 46 ][ 93 ],
   alphaCSR[ 46 ][ 94 ],
   alphaCSR[ 46 ][ 95 ],
   alphaCSR[ 46 ][ 96 ],
   alphaCSR[ 46 ][ 97 ],
   alphaCSR[ 46 ][ 98 ],
   alphaCSR[ 46 ][ 99 ],
   alphaCSR[ 46 ][ 100 ],
   alphaCSR[ 46 ][ 101 ],
   alphaCSR[ 46 ][ 102 ],
   alphaCSR[ 46 ][ 103 ],
   alphaCSR[ 46 ][ 104 ],
   alphaCSR[ 46 ][ 105 ],
   alphaCSR[ 46 ][ 106 ],
   alphaCSR[ 46 ][ 107 ],
   alphaCSR[ 46 ][ 108 ],
   alphaCSR[ 46 ][ 109 ],
   alphaCSR[ 46 ][ 110 ],
   alphaCSR[ 46 ][ 111 ],
   alphaCSR[ 46 ][ 112 ],
   alphaCSR[ 46 ][ 113 ],
   alphaCSR[ 46 ][ 114 ],
   alphaCSR[ 46 ][ 115 ],
   alphaCSR[ 46 ][ 116 ],
   alphaCSR[ 46 ][ 117 ],
   alphaCSR[ 46 ][ 118 ],
   alphaCSR[ 46 ][ 119 ],
   alphaCSR[ 46 ][ 120 ],
   alphaCSR[ 46 ][ 121 ],
   alphaCSR[ 46 ][ 122 ],
   alphaCSR[ 46 ][ 123 ],
   alphaCSR[ 46 ][ 124 ],
   alphaCSR[ 46 ][ 125 ],
   alphaCSR[ 46 ][ 126 ],
   alphaCSR[ 46 ][ 127 ],
   alphaCSR[ 46 ][ 128 ],
   alphaCSR[ 46 ][ 129 ],
   alphaCSR[ 46 ][ 130 ],
   alphaCSR[ 46 ][ 131 ],
   alphaCSR[ 46 ][ 132 ],
   alphaCSR[ 46 ][ 133 ],
   alphaCSR[ 46 ][ 134 ],
   alphaCSR[ 46 ][ 135 ],
   alphaCSR[ 46 ][ 136 ],
   alphaCSR[ 46 ][ 137 ],
   alphaCSR[ 46 ][ 138 ],
   alphaCSR[ 46 ][ 139 ],
   alphaCSR[ 46 ][ 140 ],
   alphaCSR[ 46 ][ 141 ],
   alphaCSR[ 46 ][ 142 ],
   alphaCSR[ 46 ][ 143 ],
   alphaCSR[ 46 ][ 144 ],
   alphaCSR[ 46 ][ 145 ],
   alphaCSR[ 46 ][ 146 ],
   alphaCSR[ 46 ][ 147 ],
   alphaCSR[ 46 ][ 148 ],
   alphaCSR[ 46 ][ 149 ],
   alphaCSR[ 46 ][ 150 ],
   alphaCSR[ 46 ][ 151 ],
   alphaCSR[ 46 ][ 152 ],
   alphaCSR[ 46 ][ 153 ],
   alphaCSR[ 46 ][ 154 ],
   alphaCSR[ 46 ][ 155 ],
   alphaCSR[ 46 ][ 156 ],
   alphaCSR[ 46 ][ 157 ],
   alphaCSR[ 46 ][ 158 ],
   alphaCSR[ 46 ][ 159 ],
   alphaCSR[ 46 ][ 160 ],
   alphaCSR[ 46 ][ 161 ],
   alphaCSR[ 46 ][ 162 ],
   alphaCSR[ 46 ][ 163 ],
   alphaCSR[ 46 ][ 164 ],
   alphaCSR[ 46 ][ 165 ],
   alphaCSR[ 46 ][ 166 ],
   alphaCSR[ 46 ][ 167 ],
   alphaCSR[ 46 ][ 168 ],
   alphaCSR[ 46 ][ 169 ],
   alphaCSR[ 46 ][ 170 ],
   alphaCSR[ 46 ][ 171 ],
   alphaCSR[ 46 ][ 172 ],
   alphaCSR[ 46 ][ 173 ],
   alphaCSR[ 46 ][ 174 ],
   alphaCSR[ 46 ][ 175 ],
   alphaCSR[ 46 ][ 176 ],
   alphaCSR[ 46 ][ 177 ],
   alphaCSR[ 46 ][ 178 ],
   alphaCSR[ 46 ][ 179 ],
   alphaCSR[ 46 ][ 180 ],
   alphaCSR[ 46 ][ 181 ],
   alphaCSR[ 46 ][ 182 ],
   alphaCSR[ 46 ][ 183 ],
   alphaCSR[ 46 ][ 184 ],
   alphaCSR[ 46 ][ 185 ],
   alphaCSR[ 46 ][ 186 ],
   alphaCSR[ 46 ][ 187 ],
   alphaCSR[ 46 ][ 188 ],
   alphaCSR[ 46 ][ 189 ],
   alphaCSR[ 46 ][ 190 ],
   alphaCSR[ 46 ][ 191 ],
   alphaCSR[ 46 ][ 192 ],
   alphaCSR[ 46 ][ 193 ],
   alphaCSR[ 46 ][ 194 ],
   alphaCSR[ 46 ][ 195 ],
   alphaCSR[ 46 ][ 196 ],
   alphaCSR[ 46 ][ 197 ],
   alphaCSR[ 46 ][ 198 ],
   alphaCSR[ 46 ][ 199 ],
   alphaCSR[ 46 ][ 200 ],
   alphaCSR[ 46 ][ 201 ],
   alphaCSR[ 46 ][ 202 ],
   alphaCSR[ 46 ][ 203 ],
   alphaCSR[ 46 ][ 204 ],
   alphaCSR[ 46 ][ 205 ],
   alphaCSR[ 46 ][ 206 ],
   alphaCSR[ 46 ][ 207 ],
   alphaCSR[ 46 ][ 208 ],
   alphaCSR[ 46 ][ 209 ],
   alphaCSR[ 46 ][ 210 ],
   alphaCSR[ 46 ][ 211 ],
   alphaCSR[ 46 ][ 212 ],
   alphaCSR[ 46 ][ 213 ],
   alphaCSR[ 46 ][ 214 ],
   alphaCSR[ 46 ][ 215 ],
   alphaCSR[ 46 ][ 216 ],
   alphaCSR[ 46 ][ 217 ],
   alphaCSR[ 46 ][ 218 ],
   alphaCSR[ 46 ][ 219 ],
   alphaCSR[ 46 ][ 220 ],
   alphaCSR[ 46 ][ 221 ],
   alphaCSR[ 46 ][ 222 ],
   alphaCSR[ 46 ][ 223 ],
   alphaCSR[ 46 ][ 224 ],
   alphaCSR[ 46 ][ 225 ],
   alphaCSR[ 46 ][ 226 ],
   alphaCSR[ 46 ][ 227 ],
   alphaCSR[ 46 ][ 228 ],
   alphaCSR[ 46 ][ 229 ],
   alphaCSR[ 46 ][ 230 ],
   alphaCSR[ 46 ][ 231 ],
   alphaCSR[ 46 ][ 232 ],
   alphaCSR[ 46 ][ 233 ],
   alphaCSR[ 46 ][ 234 ],
   alphaCSR[ 46 ][ 235 ],
   alphaCSR[ 46 ][ 236 ],
   alphaCSR[ 46 ][ 237 ],
   alphaCSR[ 46 ][ 238 ],
   alphaCSR[ 46 ][ 239 ],
   alphaCSR[ 46 ][ 240 ],
   alphaCSR[ 46 ][ 241 ],
   alphaCSR[ 46 ][ 242 ],
   alphaCSR[ 46 ][ 243 ],
   alphaCSR[ 46 ][ 244 ],
   alphaCSR[ 46 ][ 245 ],
   alphaCSR[ 46 ][ 246 ],
   alphaCSR[ 46 ][ 247 ],
   alphaCSR[ 46 ][ 248 ],
   alphaCSR[ 46 ][ 249 ],
   alphaCSR[ 46 ][ 250 ],
   alphaCSR[ 46 ][ 251 ],
   alphaCSR[ 46 ][ 252 ],
   alphaCSR[ 46 ][ 253 ],
   alphaCSR[ 46 ][ 254 ],
   alphaCSR[ 46 ][ 255 ],
   alphaCSR[ 46 ][ 256 ],
   alphaCSR[ 46 ][ 257 ],
   alphaCSR[ 46 ][ 258 ],
   alphaCSR[ 46 ][ 259 ],
   alphaCSR[ 46 ][ 260 ],
   alphaCSR[ 46 ][ 261 ],
   alphaCSR[ 46 ][ 262 ],
   alphaCSR[ 46 ][ 263 ],
   alphaCSR[ 46 ][ 264 ],
   alphaCSR[ 46 ][ 265 ],
   alphaCSR[ 46 ][ 266 ],
   alphaCSR[ 46 ][ 267 ],
   alphaCSR[ 46 ][ 268 ],
   alphaCSR[ 46 ][ 269 ],
   alphaCSR[ 46 ][ 270 ],
   alphaCSR[ 46 ][ 271 ],
   alphaCSR[ 46 ][ 272 ],
   alphaCSR[ 46 ][ 273 ],
   alphaCSR[ 46 ][ 274 ],
   alphaCSR[ 46 ][ 275 ],
   alphaCSR[ 46 ][ 276 ],
   alphaCSR[ 46 ][ 277 ],
   alphaCSR[ 46 ][ 278 ],
   alphaCSR[ 46 ][ 279 ],
   alphaCSR[ 46 ][ 280 ],
   alphaCSR[ 46 ][ 281 ],
   alphaCSR[ 46 ][ 282 ],
   alphaCSR[ 46 ][ 283 ],
   alphaCSR[ 46 ][ 284 ],
   alphaCSR[ 46 ][ 285 ],
   alphaCSR[ 46 ][ 286 ],
   alphaCSR[ 46 ][ 287 ],
   alphaCSR[ 46 ][ 288 ],
   alphaCSR[ 46 ][ 289 ],
   alphaCSR[ 46 ][ 290 ],
   alphaCSR[ 46 ][ 291 ],
   alphaCSR[ 46 ][ 292 ],
   alphaCSR[ 46 ][ 293 ],
   alphaCSR[ 46 ][ 294 ],
   alphaCSR[ 46 ][ 295 ],
   alphaCSR[ 46 ][ 296 ],
   alphaCSR[ 46 ][ 297 ],
   alphaCSR[ 46 ][ 298 ],
   alphaCSR[ 46 ][ 299 ],
   alphaCSR[ 46 ][ 300 ],
   alphaCSR[ 46 ][ 301 ],
   alphaCSR[ 46 ][ 302 ],
   alphaCSR[ 46 ][ 303 ],
   alphaCSR[ 46 ][ 304 ],
   alphaCSR[ 46 ][ 305 ],
   alphaCSR[ 46 ][ 306 ],
   alphaCSR[ 46 ][ 307 ],
   alphaCSR[ 46 ][ 308 ],
   alphaCSR[ 46 ][ 309 ],
   alphaCSR[ 46 ][ 310 ],
   alphaCSR[ 46 ][ 311 ],
   alphaCSR[ 46 ][ 312 ],
   alphaCSR[ 46 ][ 313 ],
   alphaCSR[ 46 ][ 314 ],
   alphaCSR[ 46 ][ 315 ],
   alphaCSR[ 46 ][ 316 ],
   alphaCSR[ 46 ][ 317 ],
   alphaCSR[ 46 ][ 318 ],
   alphaCSR[ 46 ][ 319 ],
   alphaCSR[ 46 ][ 320 ],
   alphaCSR[ 46 ][ 321 ],
   alphaCSR[ 46 ][ 322 ],
   alphaCSR[ 46 ][ 323 ],
   alphaCSR[ 46 ][ 324 ],
   alphaCSR[ 46 ][ 325 ],
   alphaCSR[ 46 ][ 326 ],
   alphaCSR[ 46 ][ 327 ],
   alphaCSR[ 46 ][ 328 ],
   alphaCSR[ 46 ][ 329 ],
   alphaCSR[ 46 ][ 330 ],
   alphaCSR[ 46 ][ 331 ],
   alphaCSR[ 46 ][ 332 ],
   alphaCSR[ 46 ][ 333 ],
   alphaCSR[ 46 ][ 334 ],
   alphaCSR[ 46 ][ 335 ],
   alphaCSR[ 46 ][ 336 ],
   alphaCSR[ 46 ][ 337 ],
   alphaCSR[ 46 ][ 338 ],
   alphaCSR[ 46 ][ 339 ],
   alphaCSR[ 46 ][ 340 ],
   alphaCSR[ 46 ][ 341 ],
   alphaCSR[ 46 ][ 342 ],
   alphaCSR[ 46 ][ 343 ],
   alphaCSR[ 46 ][ 344 ],
   alphaCSR[ 46 ][ 345 ],
   alphaCSR[ 46 ][ 346 ],
   alphaCSR[ 46 ][ 347 ],
   alphaCSR[ 46 ][ 348 ],
   alphaCSR[ 46 ][ 349 ],
   alphaCSR[ 46 ][ 350 ],
   alphaCSR[ 46 ][ 351 ],
   alphaCSR[ 46 ][ 352 ],
   alphaCSR[ 46 ][ 353 ],
   alphaCSR[ 46 ][ 354 ],
   alphaCSR[ 46 ][ 355 ],
   alphaCSR[ 46 ][ 356 ],
   alphaCSR[ 46 ][ 357 ],
   alphaCSR[ 46 ][ 358 ],
   alphaCSR[ 46 ][ 359 ],
   alphaCSR[ 46 ][ 360 ],
   alphaCSR[ 46 ][ 361 ],
   alphaCSR[ 46 ][ 362 ],
   alphaCSR[ 46 ][ 363 ],
   alphaCSR[ 46 ][ 364 ],
   alphaCSR[ 46 ][ 365 ],
   alphaCSR[ 46 ][ 366 ],
   alphaCSR[ 46 ][ 367 ],
   alphaCSR[ 46 ][ 368 ],
   alphaCSR[ 46 ][ 369 ],
   alphaCSR[ 46 ][ 370 ],
   alphaCSR[ 46 ][ 371 ],
   alphaCSR[ 46 ][ 372 ],
   alphaCSR[ 46 ][ 373 ],
   alphaCSR[ 46 ][ 374 ],
   alphaCSR[ 46 ][ 375 ],
   alphaCSR[ 46 ][ 376 ],
   alphaCSR[ 46 ][ 377 ],
   alphaCSR[ 46 ][ 378 ],
   alphaCSR[ 46 ][ 379 ],
   alphaCSR[ 46 ][ 380 ],
   alphaCSR[ 46 ][ 381 ],
   alphaCSR[ 46 ][ 382 ],
   alphaCSR[ 46 ][ 383 ],
   alphaCSR[ 47 ][ 0 ],
   alphaCSR[ 47 ][ 1 ],
   alphaCSR[ 47 ][ 2 ],
   alphaCSR[ 47 ][ 3 ],
   alphaCSR[ 47 ][ 4 ],
   alphaCSR[ 47 ][ 5 ],
   alphaCSR[ 47 ][ 6 ],
   alphaCSR[ 47 ][ 7 ],
   alphaCSR[ 47 ][ 8 ],
   alphaCSR[ 47 ][ 9 ],
   alphaCSR[ 47 ][ 10 ],
   alphaCSR[ 47 ][ 11 ],
   alphaCSR[ 47 ][ 12 ],
   alphaCSR[ 47 ][ 13 ],
   alphaCSR[ 47 ][ 14 ],
   alphaCSR[ 47 ][ 15 ],
   alphaCSR[ 47 ][ 16 ],
   alphaCSR[ 47 ][ 17 ],
   alphaCSR[ 47 ][ 18 ],
   alphaCSR[ 47 ][ 19 ],
   alphaCSR[ 47 ][ 20 ],
   alphaCSR[ 47 ][ 21 ],
   alphaCSR[ 47 ][ 22 ],
   alphaCSR[ 47 ][ 23 ],
   alphaCSR[ 47 ][ 24 ],
   alphaCSR[ 47 ][ 25 ],
   alphaCSR[ 47 ][ 26 ],
   alphaCSR[ 47 ][ 27 ],
   alphaCSR[ 47 ][ 28 ],
   alphaCSR[ 47 ][ 29 ],
   alphaCSR[ 47 ][ 30 ],
   alphaCSR[ 47 ][ 31 ],
   alphaCSR[ 47 ][ 32 ],
   alphaCSR[ 47 ][ 33 ],
   alphaCSR[ 47 ][ 34 ],
   alphaCSR[ 47 ][ 35 ],
   alphaCSR[ 47 ][ 36 ],
   alphaCSR[ 47 ][ 37 ],
   alphaCSR[ 47 ][ 38 ],
   alphaCSR[ 47 ][ 39 ],
   alphaCSR[ 47 ][ 40 ],
   alphaCSR[ 47 ][ 41 ],
   alphaCSR[ 47 ][ 42 ],
   alphaCSR[ 47 ][ 43 ],
   alphaCSR[ 47 ][ 44 ],
   alphaCSR[ 47 ][ 45 ],
   alphaCSR[ 47 ][ 46 ],
   alphaCSR[ 47 ][ 47 ],
   alphaCSR[ 47 ][ 48 ],
   alphaCSR[ 47 ][ 49 ],
   alphaCSR[ 47 ][ 50 ],
   alphaCSR[ 47 ][ 51 ],
   alphaCSR[ 47 ][ 52 ],
   alphaCSR[ 47 ][ 53 ],
   alphaCSR[ 47 ][ 54 ],
   alphaCSR[ 47 ][ 55 ],
   alphaCSR[ 47 ][ 56 ],
   alphaCSR[ 47 ][ 57 ],
   alphaCSR[ 47 ][ 58 ],
   alphaCSR[ 47 ][ 59 ],
   alphaCSR[ 47 ][ 60 ],
   alphaCSR[ 47 ][ 61 ],
   alphaCSR[ 47 ][ 62 ],
   alphaCSR[ 47 ][ 63 ],
   alphaCSR[ 47 ][ 64 ],
   alphaCSR[ 47 ][ 65 ],
   alphaCSR[ 47 ][ 66 ],
   alphaCSR[ 47 ][ 67 ],
   alphaCSR[ 47 ][ 68 ],
   alphaCSR[ 47 ][ 69 ],
   alphaCSR[ 47 ][ 70 ],
   alphaCSR[ 47 ][ 71 ],
   alphaCSR[ 47 ][ 72 ],
   alphaCSR[ 47 ][ 73 ],
   alphaCSR[ 47 ][ 74 ],
   alphaCSR[ 47 ][ 75 ],
   alphaCSR[ 47 ][ 76 ],
   alphaCSR[ 47 ][ 77 ],
   alphaCSR[ 47 ][ 78 ],
   alphaCSR[ 47 ][ 79 ],
   alphaCSR[ 47 ][ 80 ],
   alphaCSR[ 47 ][ 81 ],
   alphaCSR[ 47 ][ 82 ],
   alphaCSR[ 47 ][ 83 ],
   alphaCSR[ 47 ][ 84 ],
   alphaCSR[ 47 ][ 85 ],
   alphaCSR[ 47 ][ 86 ],
   alphaCSR[ 47 ][ 87 ],
   alphaCSR[ 47 ][ 88 ],
   alphaCSR[ 47 ][ 89 ],
   alphaCSR[ 47 ][ 90 ],
   alphaCSR[ 47 ][ 91 ],
   alphaCSR[ 47 ][ 92 ],
   alphaCSR[ 47 ][ 93 ],
   alphaCSR[ 47 ][ 94 ],
   alphaCSR[ 47 ][ 95 ],
   alphaCSR[ 47 ][ 96 ],
   alphaCSR[ 47 ][ 97 ],
   alphaCSR[ 47 ][ 98 ],
   alphaCSR[ 47 ][ 99 ],
   alphaCSR[ 47 ][ 100 ],
   alphaCSR[ 47 ][ 101 ],
   alphaCSR[ 47 ][ 102 ],
   alphaCSR[ 47 ][ 103 ],
   alphaCSR[ 47 ][ 104 ],
   alphaCSR[ 47 ][ 105 ],
   alphaCSR[ 47 ][ 106 ],
   alphaCSR[ 47 ][ 107 ],
   alphaCSR[ 47 ][ 108 ],
   alphaCSR[ 47 ][ 109 ],
   alphaCSR[ 47 ][ 110 ],
   alphaCSR[ 47 ][ 111 ],
   alphaCSR[ 47 ][ 112 ],
   alphaCSR[ 47 ][ 113 ],
   alphaCSR[ 47 ][ 114 ],
   alphaCSR[ 47 ][ 115 ],
   alphaCSR[ 47 ][ 116 ],
   alphaCSR[ 47 ][ 117 ],
   alphaCSR[ 47 ][ 118 ],
   alphaCSR[ 47 ][ 119 ],
   alphaCSR[ 47 ][ 120 ],
   alphaCSR[ 47 ][ 121 ],
   alphaCSR[ 47 ][ 122 ],
   alphaCSR[ 47 ][ 123 ],
   alphaCSR[ 47 ][ 124 ],
   alphaCSR[ 47 ][ 125 ],
   alphaCSR[ 47 ][ 126 ],
   alphaCSR[ 47 ][ 127 ],
   alphaCSR[ 47 ][ 128 ],
   alphaCSR[ 47 ][ 129 ],
   alphaCSR[ 47 ][ 130 ],
   alphaCSR[ 47 ][ 131 ],
   alphaCSR[ 47 ][ 132 ],
   alphaCSR[ 47 ][ 133 ],
   alphaCSR[ 47 ][ 134 ],
   alphaCSR[ 47 ][ 135 ],
   alphaCSR[ 47 ][ 136 ],
   alphaCSR[ 47 ][ 137 ],
   alphaCSR[ 47 ][ 138 ],
   alphaCSR[ 47 ][ 139 ],
   alphaCSR[ 47 ][ 140 ],
   alphaCSR[ 47 ][ 141 ],
   alphaCSR[ 47 ][ 142 ],
   alphaCSR[ 47 ][ 143 ],
   alphaCSR[ 47 ][ 144 ],
   alphaCSR[ 47 ][ 145 ],
   alphaCSR[ 47 ][ 146 ],
   alphaCSR[ 47 ][ 147 ],
   alphaCSR[ 47 ][ 148 ],
   alphaCSR[ 47 ][ 149 ],
   alphaCSR[ 47 ][ 150 ],
   alphaCSR[ 47 ][ 151 ],
   alphaCSR[ 47 ][ 152 ],
   alphaCSR[ 47 ][ 153 ],
   alphaCSR[ 47 ][ 154 ],
   alphaCSR[ 47 ][ 155 ],
   alphaCSR[ 47 ][ 156 ],
   alphaCSR[ 47 ][ 157 ],
   alphaCSR[ 47 ][ 158 ],
   alphaCSR[ 47 ][ 159 ],
   alphaCSR[ 47 ][ 160 ],
   alphaCSR[ 47 ][ 161 ],
   alphaCSR[ 47 ][ 162 ],
   alphaCSR[ 47 ][ 163 ],
   alphaCSR[ 47 ][ 164 ],
   alphaCSR[ 47 ][ 165 ],
   alphaCSR[ 47 ][ 166 ],
   alphaCSR[ 47 ][ 167 ],
   alphaCSR[ 47 ][ 168 ],
   alphaCSR[ 47 ][ 169 ],
   alphaCSR[ 47 ][ 170 ],
   alphaCSR[ 47 ][ 171 ],
   alphaCSR[ 47 ][ 172 ],
   alphaCSR[ 47 ][ 173 ],
   alphaCSR[ 47 ][ 174 ],
   alphaCSR[ 47 ][ 175 ],
   alphaCSR[ 47 ][ 176 ],
   alphaCSR[ 47 ][ 177 ],
   alphaCSR[ 47 ][ 178 ],
   alphaCSR[ 47 ][ 179 ],
   alphaCSR[ 47 ][ 180 ],
   alphaCSR[ 47 ][ 181 ],
   alphaCSR[ 47 ][ 182 ],
   alphaCSR[ 47 ][ 183 ],
   alphaCSR[ 47 ][ 184 ],
   alphaCSR[ 47 ][ 185 ],
   alphaCSR[ 47 ][ 186 ],
   alphaCSR[ 47 ][ 187 ],
   alphaCSR[ 47 ][ 188 ],
   alphaCSR[ 47 ][ 189 ],
   alphaCSR[ 47 ][ 190 ],
   alphaCSR[ 47 ][ 191 ],
   alphaCSR[ 47 ][ 192 ],
   alphaCSR[ 47 ][ 193 ],
   alphaCSR[ 47 ][ 194 ],
   alphaCSR[ 47 ][ 195 ],
   alphaCSR[ 47 ][ 196 ],
   alphaCSR[ 47 ][ 197 ],
   alphaCSR[ 47 ][ 198 ],
   alphaCSR[ 47 ][ 199 ],
   alphaCSR[ 47 ][ 200 ],
   alphaCSR[ 47 ][ 201 ],
   alphaCSR[ 47 ][ 202 ],
   alphaCSR[ 47 ][ 203 ],
   alphaCSR[ 47 ][ 204 ],
   alphaCSR[ 47 ][ 205 ],
   alphaCSR[ 47 ][ 206 ],
   alphaCSR[ 47 ][ 207 ],
   alphaCSR[ 47 ][ 208 ],
   alphaCSR[ 47 ][ 209 ],
   alphaCSR[ 47 ][ 210 ],
   alphaCSR[ 47 ][ 211 ],
   alphaCSR[ 47 ][ 212 ],
   alphaCSR[ 47 ][ 213 ],
   alphaCSR[ 47 ][ 214 ],
   alphaCSR[ 47 ][ 215 ],
   alphaCSR[ 47 ][ 216 ],
   alphaCSR[ 47 ][ 217 ],
   alphaCSR[ 47 ][ 218 ],
   alphaCSR[ 47 ][ 219 ],
   alphaCSR[ 47 ][ 220 ],
   alphaCSR[ 47 ][ 221 ],
   alphaCSR[ 47 ][ 222 ],
   alphaCSR[ 47 ][ 223 ],
   alphaCSR[ 47 ][ 224 ],
   alphaCSR[ 47 ][ 225 ],
   alphaCSR[ 47 ][ 226 ],
   alphaCSR[ 47 ][ 227 ],
   alphaCSR[ 47 ][ 228 ],
   alphaCSR[ 47 ][ 229 ],
   alphaCSR[ 47 ][ 230 ],
   alphaCSR[ 47 ][ 231 ],
   alphaCSR[ 47 ][ 232 ],
   alphaCSR[ 47 ][ 233 ],
   alphaCSR[ 47 ][ 234 ],
   alphaCSR[ 47 ][ 235 ],
   alphaCSR[ 47 ][ 236 ],
   alphaCSR[ 47 ][ 237 ],
   alphaCSR[ 47 ][ 238 ],
   alphaCSR[ 47 ][ 239 ],
   alphaCSR[ 47 ][ 240 ],
   alphaCSR[ 47 ][ 241 ],
   alphaCSR[ 47 ][ 242 ],
   alphaCSR[ 47 ][ 243 ],
   alphaCSR[ 47 ][ 244 ],
   alphaCSR[ 47 ][ 245 ],
   alphaCSR[ 47 ][ 246 ],
   alphaCSR[ 47 ][ 247 ],
   alphaCSR[ 47 ][ 248 ],
   alphaCSR[ 47 ][ 249 ],
   alphaCSR[ 47 ][ 250 ],
   alphaCSR[ 47 ][ 251 ],
   alphaCSR[ 47 ][ 252 ],
   alphaCSR[ 47 ][ 253 ],
   alphaCSR[ 47 ][ 254 ],
   alphaCSR[ 47 ][ 255 ],
   alphaCSR[ 47 ][ 256 ],
   alphaCSR[ 47 ][ 257 ],
   alphaCSR[ 47 ][ 258 ],
   alphaCSR[ 47 ][ 259 ],
   alphaCSR[ 47 ][ 260 ],
   alphaCSR[ 47 ][ 261 ],
   alphaCSR[ 47 ][ 262 ],
   alphaCSR[ 47 ][ 263 ],
   alphaCSR[ 47 ][ 264 ],
   alphaCSR[ 47 ][ 265 ],
   alphaCSR[ 47 ][ 266 ],
   alphaCSR[ 47 ][ 267 ],
   alphaCSR[ 47 ][ 268 ],
   alphaCSR[ 47 ][ 269 ],
   alphaCSR[ 47 ][ 270 ],
   alphaCSR[ 47 ][ 271 ],
   alphaCSR[ 47 ][ 272 ],
   alphaCSR[ 47 ][ 273 ],
   alphaCSR[ 47 ][ 274 ],
   alphaCSR[ 47 ][ 275 ],
   alphaCSR[ 47 ][ 276 ],
   alphaCSR[ 47 ][ 277 ],
   alphaCSR[ 47 ][ 278 ],
   alphaCSR[ 47 ][ 279 ],
   alphaCSR[ 47 ][ 280 ],
   alphaCSR[ 47 ][ 281 ],
   alphaCSR[ 47 ][ 282 ],
   alphaCSR[ 47 ][ 283 ],
   alphaCSR[ 47 ][ 284 ],
   alphaCSR[ 47 ][ 285 ],
   alphaCSR[ 47 ][ 286 ],
   alphaCSR[ 47 ][ 287 ],
   alphaCSR[ 47 ][ 288 ],
   alphaCSR[ 47 ][ 289 ],
   alphaCSR[ 47 ][ 290 ],
   alphaCSR[ 47 ][ 291 ],
   alphaCSR[ 47 ][ 292 ],
   alphaCSR[ 47 ][ 293 ],
   alphaCSR[ 47 ][ 294 ],
   alphaCSR[ 47 ][ 295 ],
   alphaCSR[ 47 ][ 296 ],
   alphaCSR[ 47 ][ 297 ],
   alphaCSR[ 47 ][ 298 ],
   alphaCSR[ 47 ][ 299 ],
   alphaCSR[ 47 ][ 300 ],
   alphaCSR[ 47 ][ 301 ],
   alphaCSR[ 47 ][ 302 ],
   alphaCSR[ 47 ][ 303 ],
   alphaCSR[ 47 ][ 304 ],
   alphaCSR[ 47 ][ 305 ],
   alphaCSR[ 47 ][ 306 ],
   alphaCSR[ 47 ][ 307 ],
   alphaCSR[ 47 ][ 308 ],
   alphaCSR[ 47 ][ 309 ],
   alphaCSR[ 47 ][ 310 ],
   alphaCSR[ 47 ][ 311 ],
   alphaCSR[ 47 ][ 312 ],
   alphaCSR[ 47 ][ 313 ],
   alphaCSR[ 47 ][ 314 ],
   alphaCSR[ 47 ][ 315 ],
   alphaCSR[ 47 ][ 316 ],
   alphaCSR[ 47 ][ 317 ],
   alphaCSR[ 47 ][ 318 ],
   alphaCSR[ 47 ][ 319 ],
   alphaCSR[ 47 ][ 320 ],
   alphaCSR[ 47 ][ 321 ],
   alphaCSR[ 47 ][ 322 ],
   alphaCSR[ 47 ][ 323 ],
   alphaCSR[ 47 ][ 324 ],
   alphaCSR[ 47 ][ 325 ],
   alphaCSR[ 47 ][ 326 ],
   alphaCSR[ 47 ][ 327 ],
   alphaCSR[ 47 ][ 328 ],
   alphaCSR[ 47 ][ 329 ],
   alphaCSR[ 47 ][ 330 ],
   alphaCSR[ 47 ][ 331 ],
   alphaCSR[ 47 ][ 332 ],
   alphaCSR[ 47 ][ 333 ],
   alphaCSR[ 47 ][ 334 ],
   alphaCSR[ 47 ][ 335 ],
   alphaCSR[ 47 ][ 336 ],
   alphaCSR[ 47 ][ 337 ],
   alphaCSR[ 47 ][ 338 ],
   alphaCSR[ 47 ][ 339 ],
   alphaCSR[ 47 ][ 340 ],
   alphaCSR[ 47 ][ 341 ],
   alphaCSR[ 47 ][ 342 ],
   alphaCSR[ 47 ][ 343 ],
   alphaCSR[ 47 ][ 344 ],
   alphaCSR[ 47 ][ 345 ],
   alphaCSR[ 47 ][ 346 ],
   alphaCSR[ 47 ][ 347 ],
   alphaCSR[ 47 ][ 348 ],
   alphaCSR[ 47 ][ 349 ],
   alphaCSR[ 47 ][ 350 ],
   alphaCSR[ 47 ][ 351 ],
   alphaCSR[ 47 ][ 352 ],
   alphaCSR[ 47 ][ 353 ],
   alphaCSR[ 47 ][ 354 ],
   alphaCSR[ 47 ][ 355 ],
   alphaCSR[ 47 ][ 356 ],
   alphaCSR[ 47 ][ 357 ],
   alphaCSR[ 47 ][ 358 ],
   alphaCSR[ 47 ][ 359 ],
   alphaCSR[ 47 ][ 360 ],
   alphaCSR[ 47 ][ 361 ],
   alphaCSR[ 47 ][ 362 ],
   alphaCSR[ 47 ][ 363 ],
   alphaCSR[ 47 ][ 364 ],
   alphaCSR[ 47 ][ 365 ],
   alphaCSR[ 47 ][ 366 ],
   alphaCSR[ 47 ][ 367 ],
   alphaCSR[ 47 ][ 368 ],
   alphaCSR[ 47 ][ 369 ],
   alphaCSR[ 47 ][ 370 ],
   alphaCSR[ 47 ][ 371 ],
   alphaCSR[ 47 ][ 372 ],
   alphaCSR[ 47 ][ 373 ],
   alphaCSR[ 47 ][ 374 ],
   alphaCSR[ 47 ][ 375 ],
   alphaCSR[ 47 ][ 376 ],
   alphaCSR[ 47 ][ 377 ],
   alphaCSR[ 47 ][ 378 ],
   alphaCSR[ 47 ][ 379 ],
   alphaCSR[ 47 ][ 380 ],
   alphaCSR[ 47 ][ 381 ],
   alphaCSR[ 47 ][ 382 ],
   alphaCSR[ 47 ][ 383 ],
   alphaCSR[ 48 ][ 0 ],
   alphaCSR[ 48 ][ 1 ],
   alphaCSR[ 48 ][ 2 ],
   alphaCSR[ 48 ][ 3 ],
   alphaCSR[ 48 ][ 4 ],
   alphaCSR[ 48 ][ 5 ],
   alphaCSR[ 48 ][ 6 ],
   alphaCSR[ 48 ][ 7 ],
   alphaCSR[ 48 ][ 8 ],
   alphaCSR[ 48 ][ 9 ],
   alphaCSR[ 48 ][ 10 ],
   alphaCSR[ 48 ][ 11 ],
   alphaCSR[ 48 ][ 12 ],
   alphaCSR[ 48 ][ 13 ],
   alphaCSR[ 48 ][ 14 ],
   alphaCSR[ 48 ][ 15 ],
   alphaCSR[ 48 ][ 16 ],
   alphaCSR[ 48 ][ 17 ],
   alphaCSR[ 48 ][ 18 ],
   alphaCSR[ 48 ][ 19 ],
   alphaCSR[ 48 ][ 20 ],
   alphaCSR[ 48 ][ 21 ],
   alphaCSR[ 48 ][ 22 ],
   alphaCSR[ 48 ][ 23 ],
   alphaCSR[ 48 ][ 24 ],
   alphaCSR[ 48 ][ 25 ],
   alphaCSR[ 48 ][ 26 ],
   alphaCSR[ 48 ][ 27 ],
   alphaCSR[ 48 ][ 28 ],
   alphaCSR[ 48 ][ 29 ],
   alphaCSR[ 48 ][ 30 ],
   alphaCSR[ 48 ][ 31 ],
   alphaCSR[ 48 ][ 32 ],
   alphaCSR[ 48 ][ 33 ],
   alphaCSR[ 48 ][ 34 ],
   alphaCSR[ 48 ][ 35 ],
   alphaCSR[ 48 ][ 36 ],
   alphaCSR[ 48 ][ 37 ],
   alphaCSR[ 48 ][ 38 ],
   alphaCSR[ 48 ][ 39 ],
   alphaCSR[ 48 ][ 40 ],
   alphaCSR[ 48 ][ 41 ],
   alphaCSR[ 48 ][ 42 ],
   alphaCSR[ 48 ][ 43 ],
   alphaCSR[ 48 ][ 44 ],
   alphaCSR[ 48 ][ 45 ],
   alphaCSR[ 48 ][ 46 ],
   alphaCSR[ 48 ][ 47 ],
   alphaCSR[ 48 ][ 48 ],
   alphaCSR[ 48 ][ 49 ],
   alphaCSR[ 48 ][ 50 ],
   alphaCSR[ 48 ][ 51 ],
   alphaCSR[ 48 ][ 52 ],
   alphaCSR[ 48 ][ 53 ],
   alphaCSR[ 48 ][ 54 ],
   alphaCSR[ 48 ][ 55 ],
   alphaCSR[ 48 ][ 56 ],
   alphaCSR[ 48 ][ 57 ],
   alphaCSR[ 48 ][ 58 ],
   alphaCSR[ 48 ][ 59 ],
   alphaCSR[ 48 ][ 60 ],
   alphaCSR[ 48 ][ 61 ],
   alphaCSR[ 48 ][ 62 ],
   alphaCSR[ 48 ][ 63 ],
   alphaCSR[ 48 ][ 64 ],
   alphaCSR[ 48 ][ 65 ],
   alphaCSR[ 48 ][ 66 ],
   alphaCSR[ 48 ][ 67 ],
   alphaCSR[ 48 ][ 68 ],
   alphaCSR[ 48 ][ 69 ],
   alphaCSR[ 48 ][ 70 ],
   alphaCSR[ 48 ][ 71 ],
   alphaCSR[ 48 ][ 72 ],
   alphaCSR[ 48 ][ 73 ],
   alphaCSR[ 48 ][ 74 ],
   alphaCSR[ 48 ][ 75 ],
   alphaCSR[ 48 ][ 76 ],
   alphaCSR[ 48 ][ 77 ],
   alphaCSR[ 48 ][ 78 ],
   alphaCSR[ 48 ][ 79 ],
   alphaCSR[ 48 ][ 80 ],
   alphaCSR[ 48 ][ 81 ],
   alphaCSR[ 48 ][ 82 ],
   alphaCSR[ 48 ][ 83 ],
   alphaCSR[ 48 ][ 84 ],
   alphaCSR[ 48 ][ 85 ],
   alphaCSR[ 48 ][ 86 ],
   alphaCSR[ 48 ][ 87 ],
   alphaCSR[ 48 ][ 88 ],
   alphaCSR[ 48 ][ 89 ],
   alphaCSR[ 48 ][ 90 ],
   alphaCSR[ 48 ][ 91 ],
   alphaCSR[ 48 ][ 92 ],
   alphaCSR[ 48 ][ 93 ],
   alphaCSR[ 48 ][ 94 ],
   alphaCSR[ 48 ][ 95 ],
   alphaCSR[ 48 ][ 96 ],
   alphaCSR[ 48 ][ 97 ],
   alphaCSR[ 48 ][ 98 ],
   alphaCSR[ 48 ][ 99 ],
   alphaCSR[ 48 ][ 100 ],
   alphaCSR[ 48 ][ 101 ],
   alphaCSR[ 48 ][ 102 ],
   alphaCSR[ 48 ][ 103 ],
   alphaCSR[ 48 ][ 104 ],
   alphaCSR[ 48 ][ 105 ],
   alphaCSR[ 48 ][ 106 ],
   alphaCSR[ 48 ][ 107 ],
   alphaCSR[ 48 ][ 108 ],
   alphaCSR[ 48 ][ 109 ],
   alphaCSR[ 48 ][ 110 ],
   alphaCSR[ 48 ][ 111 ],
   alphaCSR[ 48 ][ 112 ],
   alphaCSR[ 48 ][ 113 ],
   alphaCSR[ 48 ][ 114 ],
   alphaCSR[ 48 ][ 115 ],
   alphaCSR[ 48 ][ 116 ],
   alphaCSR[ 48 ][ 117 ],
   alphaCSR[ 48 ][ 118 ],
   alphaCSR[ 48 ][ 119 ],
   alphaCSR[ 48 ][ 120 ],
   alphaCSR[ 48 ][ 121 ],
   alphaCSR[ 48 ][ 122 ],
   alphaCSR[ 48 ][ 123 ],
   alphaCSR[ 48 ][ 124 ],
   alphaCSR[ 48 ][ 125 ],
   alphaCSR[ 48 ][ 126 ],
   alphaCSR[ 48 ][ 127 ],
   alphaCSR[ 48 ][ 128 ],
   alphaCSR[ 48 ][ 129 ],
   alphaCSR[ 48 ][ 130 ],
   alphaCSR[ 48 ][ 131 ],
   alphaCSR[ 48 ][ 132 ],
   alphaCSR[ 48 ][ 133 ],
   alphaCSR[ 48 ][ 134 ],
   alphaCSR[ 48 ][ 135 ],
   alphaCSR[ 48 ][ 136 ],
   alphaCSR[ 48 ][ 137 ],
   alphaCSR[ 48 ][ 138 ],
   alphaCSR[ 48 ][ 139 ],
   alphaCSR[ 48 ][ 140 ],
   alphaCSR[ 48 ][ 141 ],
   alphaCSR[ 48 ][ 142 ],
   alphaCSR[ 48 ][ 143 ],
   alphaCSR[ 48 ][ 144 ],
   alphaCSR[ 48 ][ 145 ],
   alphaCSR[ 48 ][ 146 ],
   alphaCSR[ 48 ][ 147 ],
   alphaCSR[ 48 ][ 148 ],
   alphaCSR[ 48 ][ 149 ],
   alphaCSR[ 48 ][ 150 ],
   alphaCSR[ 48 ][ 151 ],
   alphaCSR[ 48 ][ 152 ],
   alphaCSR[ 48 ][ 153 ],
   alphaCSR[ 48 ][ 154 ],
   alphaCSR[ 48 ][ 155 ],
   alphaCSR[ 48 ][ 156 ],
   alphaCSR[ 48 ][ 157 ],
   alphaCSR[ 48 ][ 158 ],
   alphaCSR[ 48 ][ 159 ],
   alphaCSR[ 48 ][ 160 ],
   alphaCSR[ 48 ][ 161 ],
   alphaCSR[ 48 ][ 162 ],
   alphaCSR[ 48 ][ 163 ],
   alphaCSR[ 48 ][ 164 ],
   alphaCSR[ 48 ][ 165 ],
   alphaCSR[ 48 ][ 166 ],
   alphaCSR[ 48 ][ 167 ],
   alphaCSR[ 48 ][ 168 ],
   alphaCSR[ 48 ][ 169 ],
   alphaCSR[ 48 ][ 170 ],
   alphaCSR[ 48 ][ 171 ],
   alphaCSR[ 48 ][ 172 ],
   alphaCSR[ 48 ][ 173 ],
   alphaCSR[ 48 ][ 174 ],
   alphaCSR[ 48 ][ 175 ],
   alphaCSR[ 48 ][ 176 ],
   alphaCSR[ 48 ][ 177 ],
   alphaCSR[ 48 ][ 178 ],
   alphaCSR[ 48 ][ 179 ],
   alphaCSR[ 48 ][ 180 ],
   alphaCSR[ 48 ][ 181 ],
   alphaCSR[ 48 ][ 182 ],
   alphaCSR[ 48 ][ 183 ],
   alphaCSR[ 48 ][ 184 ],
   alphaCSR[ 48 ][ 185 ],
   alphaCSR[ 48 ][ 186 ],
   alphaCSR[ 48 ][ 187 ],
   alphaCSR[ 48 ][ 188 ],
   alphaCSR[ 48 ][ 189 ],
   alphaCSR[ 48 ][ 190 ],
   alphaCSR[ 48 ][ 191 ],
   alphaCSR[ 48 ][ 192 ],
   alphaCSR[ 48 ][ 193 ],
   alphaCSR[ 48 ][ 194 ],
   alphaCSR[ 48 ][ 195 ],
   alphaCSR[ 48 ][ 196 ],
   alphaCSR[ 48 ][ 197 ],
   alphaCSR[ 48 ][ 198 ],
   alphaCSR[ 48 ][ 199 ],
   alphaCSR[ 48 ][ 200 ],
   alphaCSR[ 48 ][ 201 ],
   alphaCSR[ 48 ][ 202 ],
   alphaCSR[ 48 ][ 203 ],
   alphaCSR[ 48 ][ 204 ],
   alphaCSR[ 48 ][ 205 ],
   alphaCSR[ 48 ][ 206 ],
   alphaCSR[ 48 ][ 207 ],
   alphaCSR[ 48 ][ 208 ],
   alphaCSR[ 48 ][ 209 ],
   alphaCSR[ 48 ][ 210 ],
   alphaCSR[ 48 ][ 211 ],
   alphaCSR[ 48 ][ 212 ],
   alphaCSR[ 48 ][ 213 ],
   alphaCSR[ 48 ][ 214 ],
   alphaCSR[ 48 ][ 215 ],
   alphaCSR[ 48 ][ 216 ],
   alphaCSR[ 48 ][ 217 ],
   alphaCSR[ 48 ][ 218 ],
   alphaCSR[ 48 ][ 219 ],
   alphaCSR[ 48 ][ 220 ],
   alphaCSR[ 48 ][ 221 ],
   alphaCSR[ 48 ][ 222 ],
   alphaCSR[ 48 ][ 223 ],
   alphaCSR[ 48 ][ 224 ],
   alphaCSR[ 48 ][ 225 ],
   alphaCSR[ 48 ][ 226 ],
   alphaCSR[ 48 ][ 227 ],
   alphaCSR[ 48 ][ 228 ],
   alphaCSR[ 48 ][ 229 ],
   alphaCSR[ 48 ][ 230 ],
   alphaCSR[ 48 ][ 231 ],
   alphaCSR[ 48 ][ 232 ],
   alphaCSR[ 48 ][ 233 ],
   alphaCSR[ 48 ][ 234 ],
   alphaCSR[ 48 ][ 235 ],
   alphaCSR[ 48 ][ 236 ],
   alphaCSR[ 48 ][ 237 ],
   alphaCSR[ 48 ][ 238 ],
   alphaCSR[ 48 ][ 239 ],
   alphaCSR[ 48 ][ 240 ],
   alphaCSR[ 48 ][ 241 ],
   alphaCSR[ 48 ][ 242 ],
   alphaCSR[ 48 ][ 243 ],
   alphaCSR[ 48 ][ 244 ],
   alphaCSR[ 48 ][ 245 ],
   alphaCSR[ 48 ][ 246 ],
   alphaCSR[ 48 ][ 247 ],
   alphaCSR[ 48 ][ 248 ],
   alphaCSR[ 48 ][ 249 ],
   alphaCSR[ 48 ][ 250 ],
   alphaCSR[ 48 ][ 251 ],
   alphaCSR[ 48 ][ 252 ],
   alphaCSR[ 48 ][ 253 ],
   alphaCSR[ 48 ][ 254 ],
   alphaCSR[ 48 ][ 255 ],
   alphaCSR[ 48 ][ 256 ],
   alphaCSR[ 48 ][ 257 ],
   alphaCSR[ 48 ][ 258 ],
   alphaCSR[ 48 ][ 259 ],
   alphaCSR[ 48 ][ 260 ],
   alphaCSR[ 48 ][ 261 ],
   alphaCSR[ 48 ][ 262 ],
   alphaCSR[ 48 ][ 263 ],
   alphaCSR[ 48 ][ 264 ],
   alphaCSR[ 48 ][ 265 ],
   alphaCSR[ 48 ][ 266 ],
   alphaCSR[ 48 ][ 267 ],
   alphaCSR[ 48 ][ 268 ],
   alphaCSR[ 48 ][ 269 ],
   alphaCSR[ 48 ][ 270 ],
   alphaCSR[ 48 ][ 271 ],
   alphaCSR[ 48 ][ 272 ],
   alphaCSR[ 48 ][ 273 ],
   alphaCSR[ 48 ][ 274 ],
   alphaCSR[ 48 ][ 275 ],
   alphaCSR[ 48 ][ 276 ],
   alphaCSR[ 48 ][ 277 ],
   alphaCSR[ 48 ][ 278 ],
   alphaCSR[ 48 ][ 279 ],
   alphaCSR[ 48 ][ 280 ],
   alphaCSR[ 48 ][ 281 ],
   alphaCSR[ 48 ][ 282 ],
   alphaCSR[ 48 ][ 283 ],
   alphaCSR[ 48 ][ 284 ],
   alphaCSR[ 48 ][ 285 ],
   alphaCSR[ 48 ][ 286 ],
   alphaCSR[ 48 ][ 287 ],
   alphaCSR[ 48 ][ 288 ],
   alphaCSR[ 48 ][ 289 ],
   alphaCSR[ 48 ][ 290 ],
   alphaCSR[ 48 ][ 291 ],
   alphaCSR[ 48 ][ 292 ],
   alphaCSR[ 48 ][ 293 ],
   alphaCSR[ 48 ][ 294 ],
   alphaCSR[ 48 ][ 295 ],
   alphaCSR[ 48 ][ 296 ],
   alphaCSR[ 48 ][ 297 ],
   alphaCSR[ 48 ][ 298 ],
   alphaCSR[ 48 ][ 299 ],
   alphaCSR[ 48 ][ 300 ],
   alphaCSR[ 48 ][ 301 ],
   alphaCSR[ 48 ][ 302 ],
   alphaCSR[ 48 ][ 303 ],
   alphaCSR[ 48 ][ 304 ],
   alphaCSR[ 48 ][ 305 ],
   alphaCSR[ 48 ][ 306 ],
   alphaCSR[ 48 ][ 307 ],
   alphaCSR[ 48 ][ 308 ],
   alphaCSR[ 48 ][ 309 ],
   alphaCSR[ 48 ][ 310 ],
   alphaCSR[ 48 ][ 311 ],
   alphaCSR[ 48 ][ 312 ],
   alphaCSR[ 48 ][ 313 ],
   alphaCSR[ 48 ][ 314 ],
   alphaCSR[ 48 ][ 315 ],
   alphaCSR[ 48 ][ 316 ],
   alphaCSR[ 48 ][ 317 ],
   alphaCSR[ 48 ][ 318 ],
   alphaCSR[ 48 ][ 319 ],
   alphaCSR[ 48 ][ 320 ],
   alphaCSR[ 48 ][ 321 ],
   alphaCSR[ 48 ][ 322 ],
   alphaCSR[ 48 ][ 323 ],
   alphaCSR[ 48 ][ 324 ],
   alphaCSR[ 48 ][ 325 ],
   alphaCSR[ 48 ][ 326 ],
   alphaCSR[ 48 ][ 327 ],
   alphaCSR[ 48 ][ 328 ],
   alphaCSR[ 48 ][ 329 ],
   alphaCSR[ 48 ][ 330 ],
   alphaCSR[ 48 ][ 331 ],
   alphaCSR[ 48 ][ 332 ],
   alphaCSR[ 48 ][ 333 ],
   alphaCSR[ 48 ][ 334 ],
   alphaCSR[ 48 ][ 335 ],
   alphaCSR[ 48 ][ 336 ],
   alphaCSR[ 48 ][ 337 ],
   alphaCSR[ 48 ][ 338 ],
   alphaCSR[ 48 ][ 339 ],
   alphaCSR[ 48 ][ 340 ],
   alphaCSR[ 48 ][ 341 ],
   alphaCSR[ 48 ][ 342 ],
   alphaCSR[ 48 ][ 343 ],
   alphaCSR[ 48 ][ 344 ],
   alphaCSR[ 48 ][ 345 ],
   alphaCSR[ 48 ][ 346 ],
   alphaCSR[ 48 ][ 347 ],
   alphaCSR[ 48 ][ 348 ],
   alphaCSR[ 48 ][ 349 ],
   alphaCSR[ 48 ][ 350 ],
   alphaCSR[ 48 ][ 351 ],
   alphaCSR[ 48 ][ 352 ],
   alphaCSR[ 48 ][ 353 ],
   alphaCSR[ 48 ][ 354 ],
   alphaCSR[ 48 ][ 355 ],
   alphaCSR[ 48 ][ 356 ],
   alphaCSR[ 48 ][ 357 ],
   alphaCSR[ 48 ][ 358 ],
   alphaCSR[ 48 ][ 359 ],
   alphaCSR[ 48 ][ 360 ],
   alphaCSR[ 48 ][ 361 ],
   alphaCSR[ 48 ][ 362 ],
   alphaCSR[ 48 ][ 363 ],
   alphaCSR[ 48 ][ 364 ],
   alphaCSR[ 48 ][ 365 ],
   alphaCSR[ 48 ][ 366 ],
   alphaCSR[ 48 ][ 367 ],
   alphaCSR[ 48 ][ 368 ],
   alphaCSR[ 48 ][ 369 ],
   alphaCSR[ 48 ][ 370 ],
   alphaCSR[ 48 ][ 371 ],
   alphaCSR[ 48 ][ 372 ],
   alphaCSR[ 48 ][ 373 ],
   alphaCSR[ 48 ][ 374 ],
   alphaCSR[ 48 ][ 375 ],
   alphaCSR[ 48 ][ 376 ],
   alphaCSR[ 48 ][ 377 ],
   alphaCSR[ 48 ][ 378 ],
   alphaCSR[ 48 ][ 379 ],
   alphaCSR[ 48 ][ 380 ],
   alphaCSR[ 48 ][ 381 ],
   alphaCSR[ 48 ][ 382 ],
   alphaCSR[ 48 ][ 383 ],
   alphaCSR[ 49 ][ 0 ],
   alphaCSR[ 49 ][ 1 ],
   alphaCSR[ 49 ][ 2 ],
   alphaCSR[ 49 ][ 3 ],
   alphaCSR[ 49 ][ 4 ],
   alphaCSR[ 49 ][ 5 ],
   alphaCSR[ 49 ][ 6 ],
   alphaCSR[ 49 ][ 7 ],
   alphaCSR[ 49 ][ 8 ],
   alphaCSR[ 49 ][ 9 ],
   alphaCSR[ 49 ][ 10 ],
   alphaCSR[ 49 ][ 11 ],
   alphaCSR[ 49 ][ 12 ],
   alphaCSR[ 49 ][ 13 ],
   alphaCSR[ 49 ][ 14 ],
   alphaCSR[ 49 ][ 15 ],
   alphaCSR[ 49 ][ 16 ],
   alphaCSR[ 49 ][ 17 ],
   alphaCSR[ 49 ][ 18 ],
   alphaCSR[ 49 ][ 19 ],
   alphaCSR[ 49 ][ 20 ],
   alphaCSR[ 49 ][ 21 ],
   alphaCSR[ 49 ][ 22 ],
   alphaCSR[ 49 ][ 23 ],
   alphaCSR[ 49 ][ 24 ],
   alphaCSR[ 49 ][ 25 ],
   alphaCSR[ 49 ][ 26 ],
   alphaCSR[ 49 ][ 27 ],
   alphaCSR[ 49 ][ 28 ],
   alphaCSR[ 49 ][ 29 ],
   alphaCSR[ 49 ][ 30 ],
   alphaCSR[ 49 ][ 31 ],
   alphaCSR[ 49 ][ 32 ],
   alphaCSR[ 49 ][ 33 ],
   alphaCSR[ 49 ][ 34 ],
   alphaCSR[ 49 ][ 35 ],
   alphaCSR[ 49 ][ 36 ],
   alphaCSR[ 49 ][ 37 ],
   alphaCSR[ 49 ][ 38 ],
   alphaCSR[ 49 ][ 39 ],
   alphaCSR[ 49 ][ 40 ],
   alphaCSR[ 49 ][ 41 ],
   alphaCSR[ 49 ][ 42 ],
   alphaCSR[ 49 ][ 43 ],
   alphaCSR[ 49 ][ 44 ],
   alphaCSR[ 49 ][ 45 ],
   alphaCSR[ 49 ][ 46 ],
   alphaCSR[ 49 ][ 47 ],
   alphaCSR[ 49 ][ 48 ],
   alphaCSR[ 49 ][ 49 ],
   alphaCSR[ 49 ][ 50 ],
   alphaCSR[ 49 ][ 51 ],
   alphaCSR[ 49 ][ 52 ],
   alphaCSR[ 49 ][ 53 ],
   alphaCSR[ 49 ][ 54 ],
   alphaCSR[ 49 ][ 55 ],
   alphaCSR[ 49 ][ 56 ],
   alphaCSR[ 49 ][ 57 ],
   alphaCSR[ 49 ][ 58 ],
   alphaCSR[ 49 ][ 59 ],
   alphaCSR[ 49 ][ 60 ],
   alphaCSR[ 49 ][ 61 ],
   alphaCSR[ 49 ][ 62 ],
   alphaCSR[ 49 ][ 63 ],
   alphaCSR[ 49 ][ 64 ],
   alphaCSR[ 49 ][ 65 ],
   alphaCSR[ 49 ][ 66 ],
   alphaCSR[ 49 ][ 67 ],
   alphaCSR[ 49 ][ 68 ],
   alphaCSR[ 49 ][ 69 ],
   alphaCSR[ 49 ][ 70 ],
   alphaCSR[ 49 ][ 71 ],
   alphaCSR[ 49 ][ 72 ],
   alphaCSR[ 49 ][ 73 ],
   alphaCSR[ 49 ][ 74 ],
   alphaCSR[ 49 ][ 75 ],
   alphaCSR[ 49 ][ 76 ],
   alphaCSR[ 49 ][ 77 ],
   alphaCSR[ 49 ][ 78 ],
   alphaCSR[ 49 ][ 79 ],
   alphaCSR[ 49 ][ 80 ],
   alphaCSR[ 49 ][ 81 ],
   alphaCSR[ 49 ][ 82 ],
   alphaCSR[ 49 ][ 83 ],
   alphaCSR[ 49 ][ 84 ],
   alphaCSR[ 49 ][ 85 ],
   alphaCSR[ 49 ][ 86 ],
   alphaCSR[ 49 ][ 87 ],
   alphaCSR[ 49 ][ 88 ],
   alphaCSR[ 49 ][ 89 ],
   alphaCSR[ 49 ][ 90 ],
   alphaCSR[ 49 ][ 91 ],
   alphaCSR[ 49 ][ 92 ],
   alphaCSR[ 49 ][ 93 ],
   alphaCSR[ 49 ][ 94 ],
   alphaCSR[ 49 ][ 95 ],
   alphaCSR[ 49 ][ 96 ],
   alphaCSR[ 49 ][ 97 ],
   alphaCSR[ 49 ][ 98 ],
   alphaCSR[ 49 ][ 99 ],
   alphaCSR[ 49 ][ 100 ],
   alphaCSR[ 49 ][ 101 ],
   alphaCSR[ 49 ][ 102 ],
   alphaCSR[ 49 ][ 103 ],
   alphaCSR[ 49 ][ 104 ],
   alphaCSR[ 49 ][ 105 ],
   alphaCSR[ 49 ][ 106 ],
   alphaCSR[ 49 ][ 107 ],
   alphaCSR[ 49 ][ 108 ],
   alphaCSR[ 49 ][ 109 ],
   alphaCSR[ 49 ][ 110 ],
   alphaCSR[ 49 ][ 111 ],
   alphaCSR[ 49 ][ 112 ],
   alphaCSR[ 49 ][ 113 ],
   alphaCSR[ 49 ][ 114 ],
   alphaCSR[ 49 ][ 115 ],
   alphaCSR[ 49 ][ 116 ],
   alphaCSR[ 49 ][ 117 ],
   alphaCSR[ 49 ][ 118 ],
   alphaCSR[ 49 ][ 119 ],
   alphaCSR[ 49 ][ 120 ],
   alphaCSR[ 49 ][ 121 ],
   alphaCSR[ 49 ][ 122 ],
   alphaCSR[ 49 ][ 123 ],
   alphaCSR[ 49 ][ 124 ],
   alphaCSR[ 49 ][ 125 ],
   alphaCSR[ 49 ][ 126 ],
   alphaCSR[ 49 ][ 127 ],
   alphaCSR[ 49 ][ 128 ],
   alphaCSR[ 49 ][ 129 ],
   alphaCSR[ 49 ][ 130 ],
   alphaCSR[ 49 ][ 131 ],
   alphaCSR[ 49 ][ 132 ],
   alphaCSR[ 49 ][ 133 ],
   alphaCSR[ 49 ][ 134 ],
   alphaCSR[ 49 ][ 135 ],
   alphaCSR[ 49 ][ 136 ],
   alphaCSR[ 49 ][ 137 ],
   alphaCSR[ 49 ][ 138 ],
   alphaCSR[ 49 ][ 139 ],
   alphaCSR[ 49 ][ 140 ],
   alphaCSR[ 49 ][ 141 ],
   alphaCSR[ 49 ][ 142 ],
   alphaCSR[ 49 ][ 143 ],
   alphaCSR[ 49 ][ 144 ],
   alphaCSR[ 49 ][ 145 ],
   alphaCSR[ 49 ][ 146 ],
   alphaCSR[ 49 ][ 147 ],
   alphaCSR[ 49 ][ 148 ],
   alphaCSR[ 49 ][ 149 ],
   alphaCSR[ 49 ][ 150 ],
   alphaCSR[ 49 ][ 151 ],
   alphaCSR[ 49 ][ 152 ],
   alphaCSR[ 49 ][ 153 ],
   alphaCSR[ 49 ][ 154 ],
   alphaCSR[ 49 ][ 155 ],
   alphaCSR[ 49 ][ 156 ],
   alphaCSR[ 49 ][ 157 ],
   alphaCSR[ 49 ][ 158 ],
   alphaCSR[ 49 ][ 159 ],
   alphaCSR[ 49 ][ 160 ],
   alphaCSR[ 49 ][ 161 ],
   alphaCSR[ 49 ][ 162 ],
   alphaCSR[ 49 ][ 163 ],
   alphaCSR[ 49 ][ 164 ],
   alphaCSR[ 49 ][ 165 ],
   alphaCSR[ 49 ][ 166 ],
   alphaCSR[ 49 ][ 167 ],
   alphaCSR[ 49 ][ 168 ],
   alphaCSR[ 49 ][ 169 ],
   alphaCSR[ 49 ][ 170 ],
   alphaCSR[ 49 ][ 171 ],
   alphaCSR[ 49 ][ 172 ],
   alphaCSR[ 49 ][ 173 ],
   alphaCSR[ 49 ][ 174 ],
   alphaCSR[ 49 ][ 175 ],
   alphaCSR[ 49 ][ 176 ],
   alphaCSR[ 49 ][ 177 ],
   alphaCSR[ 49 ][ 178 ],
   alphaCSR[ 49 ][ 179 ],
   alphaCSR[ 49 ][ 180 ],
   alphaCSR[ 49 ][ 181 ],
   alphaCSR[ 49 ][ 182 ],
   alphaCSR[ 49 ][ 183 ],
   alphaCSR[ 49 ][ 184 ],
   alphaCSR[ 49 ][ 185 ],
   alphaCSR[ 49 ][ 186 ],
   alphaCSR[ 49 ][ 187 ],
   alphaCSR[ 49 ][ 188 ],
   alphaCSR[ 49 ][ 189 ],
   alphaCSR[ 49 ][ 190 ],
   alphaCSR[ 49 ][ 191 ],
   alphaCSR[ 49 ][ 192 ],
   alphaCSR[ 49 ][ 193 ],
   alphaCSR[ 49 ][ 194 ],
   alphaCSR[ 49 ][ 195 ],
   alphaCSR[ 49 ][ 196 ],
   alphaCSR[ 49 ][ 197 ],
   alphaCSR[ 49 ][ 198 ],
   alphaCSR[ 49 ][ 199 ],
   alphaCSR[ 49 ][ 200 ],
   alphaCSR[ 49 ][ 201 ],
   alphaCSR[ 49 ][ 202 ],
   alphaCSR[ 49 ][ 203 ],
   alphaCSR[ 49 ][ 204 ],
   alphaCSR[ 49 ][ 205 ],
   alphaCSR[ 49 ][ 206 ],
   alphaCSR[ 49 ][ 207 ],
   alphaCSR[ 49 ][ 208 ],
   alphaCSR[ 49 ][ 209 ],
   alphaCSR[ 49 ][ 210 ],
   alphaCSR[ 49 ][ 211 ],
   alphaCSR[ 49 ][ 212 ],
   alphaCSR[ 49 ][ 213 ],
   alphaCSR[ 49 ][ 214 ],
   alphaCSR[ 49 ][ 215 ],
   alphaCSR[ 49 ][ 216 ],
   alphaCSR[ 49 ][ 217 ],
   alphaCSR[ 49 ][ 218 ],
   alphaCSR[ 49 ][ 219 ],
   alphaCSR[ 49 ][ 220 ],
   alphaCSR[ 49 ][ 221 ],
   alphaCSR[ 49 ][ 222 ],
   alphaCSR[ 49 ][ 223 ],
   alphaCSR[ 49 ][ 224 ],
   alphaCSR[ 49 ][ 225 ],
   alphaCSR[ 49 ][ 226 ],
   alphaCSR[ 49 ][ 227 ],
   alphaCSR[ 49 ][ 228 ],
   alphaCSR[ 49 ][ 229 ],
   alphaCSR[ 49 ][ 230 ],
   alphaCSR[ 49 ][ 231 ],
   alphaCSR[ 49 ][ 232 ],
   alphaCSR[ 49 ][ 233 ],
   alphaCSR[ 49 ][ 234 ],
   alphaCSR[ 49 ][ 235 ],
   alphaCSR[ 49 ][ 236 ],
   alphaCSR[ 49 ][ 237 ],
   alphaCSR[ 49 ][ 238 ],
   alphaCSR[ 49 ][ 239 ],
   alphaCSR[ 49 ][ 240 ],
   alphaCSR[ 49 ][ 241 ],
   alphaCSR[ 49 ][ 242 ],
   alphaCSR[ 49 ][ 243 ],
   alphaCSR[ 49 ][ 244 ],
   alphaCSR[ 49 ][ 245 ],
   alphaCSR[ 49 ][ 246 ],
   alphaCSR[ 49 ][ 247 ],
   alphaCSR[ 49 ][ 248 ],
   alphaCSR[ 49 ][ 249 ],
   alphaCSR[ 49 ][ 250 ],
   alphaCSR[ 49 ][ 251 ],
   alphaCSR[ 49 ][ 252 ],
   alphaCSR[ 49 ][ 253 ],
   alphaCSR[ 49 ][ 254 ],
   alphaCSR[ 49 ][ 255 ],
   alphaCSR[ 49 ][ 256 ],
   alphaCSR[ 49 ][ 257 ],
   alphaCSR[ 49 ][ 258 ],
   alphaCSR[ 49 ][ 259 ],
   alphaCSR[ 49 ][ 260 ],
   alphaCSR[ 49 ][ 261 ],
   alphaCSR[ 49 ][ 262 ],
   alphaCSR[ 49 ][ 263 ],
   alphaCSR[ 49 ][ 264 ],
   alphaCSR[ 49 ][ 265 ],
   alphaCSR[ 49 ][ 266 ],
   alphaCSR[ 49 ][ 267 ],
   alphaCSR[ 49 ][ 268 ],
   alphaCSR[ 49 ][ 269 ],
   alphaCSR[ 49 ][ 270 ],
   alphaCSR[ 49 ][ 271 ],
   alphaCSR[ 49 ][ 272 ],
   alphaCSR[ 49 ][ 273 ],
   alphaCSR[ 49 ][ 274 ],
   alphaCSR[ 49 ][ 275 ],
   alphaCSR[ 49 ][ 276 ],
   alphaCSR[ 49 ][ 277 ],
   alphaCSR[ 49 ][ 278 ],
   alphaCSR[ 49 ][ 279 ],
   alphaCSR[ 49 ][ 280 ],
   alphaCSR[ 49 ][ 281 ],
   alphaCSR[ 49 ][ 282 ],
   alphaCSR[ 49 ][ 283 ],
   alphaCSR[ 49 ][ 284 ],
   alphaCSR[ 49 ][ 285 ],
   alphaCSR[ 49 ][ 286 ],
   alphaCSR[ 49 ][ 287 ],
   alphaCSR[ 49 ][ 288 ],
   alphaCSR[ 49 ][ 289 ],
   alphaCSR[ 49 ][ 290 ],
   alphaCSR[ 49 ][ 291 ],
   alphaCSR[ 49 ][ 292 ],
   alphaCSR[ 49 ][ 293 ],
   alphaCSR[ 49 ][ 294 ],
   alphaCSR[ 49 ][ 295 ],
   alphaCSR[ 49 ][ 296 ],
   alphaCSR[ 49 ][ 297 ],
   alphaCSR[ 49 ][ 298 ],
   alphaCSR[ 49 ][ 299 ],
   alphaCSR[ 49 ][ 300 ],
   alphaCSR[ 49 ][ 301 ],
   alphaCSR[ 49 ][ 302 ],
   alphaCSR[ 49 ][ 303 ],
   alphaCSR[ 49 ][ 304 ],
   alphaCSR[ 49 ][ 305 ],
   alphaCSR[ 49 ][ 306 ],
   alphaCSR[ 49 ][ 307 ],
   alphaCSR[ 49 ][ 308 ],
   alphaCSR[ 49 ][ 309 ],
   alphaCSR[ 49 ][ 310 ],
   alphaCSR[ 49 ][ 311 ],
   alphaCSR[ 49 ][ 312 ],
   alphaCSR[ 49 ][ 313 ],
   alphaCSR[ 49 ][ 314 ],
   alphaCSR[ 49 ][ 315 ],
   alphaCSR[ 49 ][ 316 ],
   alphaCSR[ 49 ][ 317 ],
   alphaCSR[ 49 ][ 318 ],
   alphaCSR[ 49 ][ 319 ],
   alphaCSR[ 49 ][ 320 ],
   alphaCSR[ 49 ][ 321 ],
   alphaCSR[ 49 ][ 322 ],
   alphaCSR[ 49 ][ 323 ],
   alphaCSR[ 49 ][ 324 ],
   alphaCSR[ 49 ][ 325 ],
   alphaCSR[ 49 ][ 326 ],
   alphaCSR[ 49 ][ 327 ],
   alphaCSR[ 49 ][ 328 ],
   alphaCSR[ 49 ][ 329 ],
   alphaCSR[ 49 ][ 330 ],
   alphaCSR[ 49 ][ 331 ],
   alphaCSR[ 49 ][ 332 ],
   alphaCSR[ 49 ][ 333 ],
   alphaCSR[ 49 ][ 334 ],
   alphaCSR[ 49 ][ 335 ],
   alphaCSR[ 49 ][ 336 ],
   alphaCSR[ 49 ][ 337 ],
   alphaCSR[ 49 ][ 338 ],
   alphaCSR[ 49 ][ 339 ],
   alphaCSR[ 49 ][ 340 ],
   alphaCSR[ 49 ][ 341 ],
   alphaCSR[ 49 ][ 342 ],
   alphaCSR[ 49 ][ 343 ],
   alphaCSR[ 49 ][ 344 ],
   alphaCSR[ 49 ][ 345 ],
   alphaCSR[ 49 ][ 346 ],
   alphaCSR[ 49 ][ 347 ],
   alphaCSR[ 49 ][ 348 ],
   alphaCSR[ 49 ][ 349 ],
   alphaCSR[ 49 ][ 350 ],
   alphaCSR[ 49 ][ 351 ],
   alphaCSR[ 49 ][ 352 ],
   alphaCSR[ 49 ][ 353 ],
   alphaCSR[ 49 ][ 354 ],
   alphaCSR[ 49 ][ 355 ],
   alphaCSR[ 49 ][ 356 ],
   alphaCSR[ 49 ][ 357 ],
   alphaCSR[ 49 ][ 358 ],
   alphaCSR[ 49 ][ 359 ],
   alphaCSR[ 49 ][ 360 ],
   alphaCSR[ 49 ][ 361 ],
   alphaCSR[ 49 ][ 362 ],
   alphaCSR[ 49 ][ 363 ],
   alphaCSR[ 49 ][ 364 ],
   alphaCSR[ 49 ][ 365 ],
   alphaCSR[ 49 ][ 366 ],
   alphaCSR[ 49 ][ 367 ],
   alphaCSR[ 49 ][ 368 ],
   alphaCSR[ 49 ][ 369 ],
   alphaCSR[ 49 ][ 370 ],
   alphaCSR[ 49 ][ 371 ],
   alphaCSR[ 49 ][ 372 ],
   alphaCSR[ 49 ][ 373 ],
   alphaCSR[ 49 ][ 374 ],
   alphaCSR[ 49 ][ 375 ],
   alphaCSR[ 49 ][ 376 ],
   alphaCSR[ 49 ][ 377 ],
   alphaCSR[ 49 ][ 378 ],
   alphaCSR[ 49 ][ 379 ],
   alphaCSR[ 49 ][ 380 ],
   alphaCSR[ 49 ][ 381 ],
   alphaCSR[ 49 ][ 382 ],
   alphaCSR[ 49 ][ 383 ],
   alphaCSR[ 50 ][ 0 ],
   alphaCSR[ 50 ][ 1 ],
   alphaCSR[ 50 ][ 2 ],
   alphaCSR[ 50 ][ 3 ],
   alphaCSR[ 50 ][ 4 ],
   alphaCSR[ 50 ][ 5 ],
   alphaCSR[ 50 ][ 6 ],
   alphaCSR[ 50 ][ 7 ],
   alphaCSR[ 50 ][ 8 ],
   alphaCSR[ 50 ][ 9 ],
   alphaCSR[ 50 ][ 10 ],
   alphaCSR[ 50 ][ 11 ],
   alphaCSR[ 50 ][ 12 ],
   alphaCSR[ 50 ][ 13 ],
   alphaCSR[ 50 ][ 14 ],
   alphaCSR[ 50 ][ 15 ],
   alphaCSR[ 50 ][ 16 ],
   alphaCSR[ 50 ][ 17 ],
   alphaCSR[ 50 ][ 18 ],
   alphaCSR[ 50 ][ 19 ],
   alphaCSR[ 50 ][ 20 ],
   alphaCSR[ 50 ][ 21 ],
   alphaCSR[ 50 ][ 22 ],
   alphaCSR[ 50 ][ 23 ],
   alphaCSR[ 50 ][ 24 ],
   alphaCSR[ 50 ][ 25 ],
   alphaCSR[ 50 ][ 26 ],
   alphaCSR[ 50 ][ 27 ],
   alphaCSR[ 50 ][ 28 ],
   alphaCSR[ 50 ][ 29 ],
   alphaCSR[ 50 ][ 30 ],
   alphaCSR[ 50 ][ 31 ],
   alphaCSR[ 50 ][ 32 ],
   alphaCSR[ 50 ][ 33 ],
   alphaCSR[ 50 ][ 34 ],
   alphaCSR[ 50 ][ 35 ],
   alphaCSR[ 50 ][ 36 ],
   alphaCSR[ 50 ][ 37 ],
   alphaCSR[ 50 ][ 38 ],
   alphaCSR[ 50 ][ 39 ],
   alphaCSR[ 50 ][ 40 ],
   alphaCSR[ 50 ][ 41 ],
   alphaCSR[ 50 ][ 42 ],
   alphaCSR[ 50 ][ 43 ],
   alphaCSR[ 50 ][ 44 ],
   alphaCSR[ 50 ][ 45 ],
   alphaCSR[ 50 ][ 46 ],
   alphaCSR[ 50 ][ 47 ],
   alphaCSR[ 50 ][ 48 ],
   alphaCSR[ 50 ][ 49 ],
   alphaCSR[ 50 ][ 50 ],
   alphaCSR[ 50 ][ 51 ],
   alphaCSR[ 50 ][ 52 ],
   alphaCSR[ 50 ][ 53 ],
   alphaCSR[ 50 ][ 54 ],
   alphaCSR[ 50 ][ 55 ],
   alphaCSR[ 50 ][ 56 ],
   alphaCSR[ 50 ][ 57 ],
   alphaCSR[ 50 ][ 58 ],
   alphaCSR[ 50 ][ 59 ],
   alphaCSR[ 50 ][ 60 ],
   alphaCSR[ 50 ][ 61 ],
   alphaCSR[ 50 ][ 62 ],
   alphaCSR[ 50 ][ 63 ],
   alphaCSR[ 50 ][ 64 ],
   alphaCSR[ 50 ][ 65 ],
   alphaCSR[ 50 ][ 66 ],
   alphaCSR[ 50 ][ 67 ],
   alphaCSR[ 50 ][ 68 ],
   alphaCSR[ 50 ][ 69 ],
   alphaCSR[ 50 ][ 70 ],
   alphaCSR[ 50 ][ 71 ],
   alphaCSR[ 50 ][ 72 ],
   alphaCSR[ 50 ][ 73 ],
   alphaCSR[ 50 ][ 74 ],
   alphaCSR[ 50 ][ 75 ],
   alphaCSR[ 50 ][ 76 ],
   alphaCSR[ 50 ][ 77 ],
   alphaCSR[ 50 ][ 78 ],
   alphaCSR[ 50 ][ 79 ],
   alphaCSR[ 50 ][ 80 ],
   alphaCSR[ 50 ][ 81 ],
   alphaCSR[ 50 ][ 82 ],
   alphaCSR[ 50 ][ 83 ],
   alphaCSR[ 50 ][ 84 ],
   alphaCSR[ 50 ][ 85 ],
   alphaCSR[ 50 ][ 86 ],
   alphaCSR[ 50 ][ 87 ],
   alphaCSR[ 50 ][ 88 ],
   alphaCSR[ 50 ][ 89 ],
   alphaCSR[ 50 ][ 90 ],
   alphaCSR[ 50 ][ 91 ],
   alphaCSR[ 50 ][ 92 ],
   alphaCSR[ 50 ][ 93 ],
   alphaCSR[ 50 ][ 94 ],
   alphaCSR[ 50 ][ 95 ],
   alphaCSR[ 50 ][ 96 ],
   alphaCSR[ 50 ][ 97 ],
   alphaCSR[ 50 ][ 98 ],
   alphaCSR[ 50 ][ 99 ],
   alphaCSR[ 50 ][ 100 ],
   alphaCSR[ 50 ][ 101 ],
   alphaCSR[ 50 ][ 102 ],
   alphaCSR[ 50 ][ 103 ],
   alphaCSR[ 50 ][ 104 ],
   alphaCSR[ 50 ][ 105 ],
   alphaCSR[ 50 ][ 106 ],
   alphaCSR[ 50 ][ 107 ],
   alphaCSR[ 50 ][ 108 ],
   alphaCSR[ 50 ][ 109 ],
   alphaCSR[ 50 ][ 110 ],
   alphaCSR[ 50 ][ 111 ],
   alphaCSR[ 50 ][ 112 ],
   alphaCSR[ 50 ][ 113 ],
   alphaCSR[ 50 ][ 114 ],
   alphaCSR[ 50 ][ 115 ],
   alphaCSR[ 50 ][ 116 ],
   alphaCSR[ 50 ][ 117 ],
   alphaCSR[ 50 ][ 118 ],
   alphaCSR[ 50 ][ 119 ],
   alphaCSR[ 50 ][ 120 ],
   alphaCSR[ 50 ][ 121 ],
   alphaCSR[ 50 ][ 122 ],
   alphaCSR[ 50 ][ 123 ],
   alphaCSR[ 50 ][ 124 ],
   alphaCSR[ 50 ][ 125 ],
   alphaCSR[ 50 ][ 126 ],
   alphaCSR[ 50 ][ 127 ],
   alphaCSR[ 50 ][ 128 ],
   alphaCSR[ 50 ][ 129 ],
   alphaCSR[ 50 ][ 130 ],
   alphaCSR[ 50 ][ 131 ],
   alphaCSR[ 50 ][ 132 ],
   alphaCSR[ 50 ][ 133 ],
   alphaCSR[ 50 ][ 134 ],
   alphaCSR[ 50 ][ 135 ],
   alphaCSR[ 50 ][ 136 ],
   alphaCSR[ 50 ][ 137 ],
   alphaCSR[ 50 ][ 138 ],
   alphaCSR[ 50 ][ 139 ],
   alphaCSR[ 50 ][ 140 ],
   alphaCSR[ 50 ][ 141 ],
   alphaCSR[ 50 ][ 142 ],
   alphaCSR[ 50 ][ 143 ],
   alphaCSR[ 50 ][ 144 ],
   alphaCSR[ 50 ][ 145 ],
   alphaCSR[ 50 ][ 146 ],
   alphaCSR[ 50 ][ 147 ],
   alphaCSR[ 50 ][ 148 ],
   alphaCSR[ 50 ][ 149 ],
   alphaCSR[ 50 ][ 150 ],
   alphaCSR[ 50 ][ 151 ],
   alphaCSR[ 50 ][ 152 ],
   alphaCSR[ 50 ][ 153 ],
   alphaCSR[ 50 ][ 154 ],
   alphaCSR[ 50 ][ 155 ],
   alphaCSR[ 50 ][ 156 ],
   alphaCSR[ 50 ][ 157 ],
   alphaCSR[ 50 ][ 158 ],
   alphaCSR[ 50 ][ 159 ],
   alphaCSR[ 50 ][ 160 ],
   alphaCSR[ 50 ][ 161 ],
   alphaCSR[ 50 ][ 162 ],
   alphaCSR[ 50 ][ 163 ],
   alphaCSR[ 50 ][ 164 ],
   alphaCSR[ 50 ][ 165 ],
   alphaCSR[ 50 ][ 166 ],
   alphaCSR[ 50 ][ 167 ],
   alphaCSR[ 50 ][ 168 ],
   alphaCSR[ 50 ][ 169 ],
   alphaCSR[ 50 ][ 170 ],
   alphaCSR[ 50 ][ 171 ],
   alphaCSR[ 50 ][ 172 ],
   alphaCSR[ 50 ][ 173 ],
   alphaCSR[ 50 ][ 174 ],
   alphaCSR[ 50 ][ 175 ],
   alphaCSR[ 50 ][ 176 ],
   alphaCSR[ 50 ][ 177 ],
   alphaCSR[ 50 ][ 178 ],
   alphaCSR[ 50 ][ 179 ],
   alphaCSR[ 50 ][ 180 ],
   alphaCSR[ 50 ][ 181 ],
   alphaCSR[ 50 ][ 182 ],
   alphaCSR[ 50 ][ 183 ],
   alphaCSR[ 50 ][ 184 ],
   alphaCSR[ 50 ][ 185 ],
   alphaCSR[ 50 ][ 186 ],
   alphaCSR[ 50 ][ 187 ],
   alphaCSR[ 50 ][ 188 ],
   alphaCSR[ 50 ][ 189 ],
   alphaCSR[ 50 ][ 190 ],
   alphaCSR[ 50 ][ 191 ],
   alphaCSR[ 50 ][ 192 ],
   alphaCSR[ 50 ][ 193 ],
   alphaCSR[ 50 ][ 194 ],
   alphaCSR[ 50 ][ 195 ],
   alphaCSR[ 50 ][ 196 ],
   alphaCSR[ 50 ][ 197 ],
   alphaCSR[ 50 ][ 198 ],
   alphaCSR[ 50 ][ 199 ],
   alphaCSR[ 50 ][ 200 ],
   alphaCSR[ 50 ][ 201 ],
   alphaCSR[ 50 ][ 202 ],
   alphaCSR[ 50 ][ 203 ],
   alphaCSR[ 50 ][ 204 ],
   alphaCSR[ 50 ][ 205 ],
   alphaCSR[ 50 ][ 206 ],
   alphaCSR[ 50 ][ 207 ],
   alphaCSR[ 50 ][ 208 ],
   alphaCSR[ 50 ][ 209 ],
   alphaCSR[ 50 ][ 210 ],
   alphaCSR[ 50 ][ 211 ],
   alphaCSR[ 50 ][ 212 ],
   alphaCSR[ 50 ][ 213 ],
   alphaCSR[ 50 ][ 214 ],
   alphaCSR[ 50 ][ 215 ],
   alphaCSR[ 50 ][ 216 ],
   alphaCSR[ 50 ][ 217 ],
   alphaCSR[ 50 ][ 218 ],
   alphaCSR[ 50 ][ 219 ],
   alphaCSR[ 50 ][ 220 ],
   alphaCSR[ 50 ][ 221 ],
   alphaCSR[ 50 ][ 222 ],
   alphaCSR[ 50 ][ 223 ],
   alphaCSR[ 50 ][ 224 ],
   alphaCSR[ 50 ][ 225 ],
   alphaCSR[ 50 ][ 226 ],
   alphaCSR[ 50 ][ 227 ],
   alphaCSR[ 50 ][ 228 ],
   alphaCSR[ 50 ][ 229 ],
   alphaCSR[ 50 ][ 230 ],
   alphaCSR[ 50 ][ 231 ],
   alphaCSR[ 50 ][ 232 ],
   alphaCSR[ 50 ][ 233 ],
   alphaCSR[ 50 ][ 234 ],
   alphaCSR[ 50 ][ 235 ],
   alphaCSR[ 50 ][ 236 ],
   alphaCSR[ 50 ][ 237 ],
   alphaCSR[ 50 ][ 238 ],
   alphaCSR[ 50 ][ 239 ],
   alphaCSR[ 50 ][ 240 ],
   alphaCSR[ 50 ][ 241 ],
   alphaCSR[ 50 ][ 242 ],
   alphaCSR[ 50 ][ 243 ],
   alphaCSR[ 50 ][ 244 ],
   alphaCSR[ 50 ][ 245 ],
   alphaCSR[ 50 ][ 246 ],
   alphaCSR[ 50 ][ 247 ],
   alphaCSR[ 50 ][ 248 ],
   alphaCSR[ 50 ][ 249 ],
   alphaCSR[ 50 ][ 250 ],
   alphaCSR[ 50 ][ 251 ],
   alphaCSR[ 50 ][ 252 ],
   alphaCSR[ 50 ][ 253 ],
   alphaCSR[ 50 ][ 254 ],
   alphaCSR[ 50 ][ 255 ],
   alphaCSR[ 50 ][ 256 ],
   alphaCSR[ 50 ][ 257 ],
   alphaCSR[ 50 ][ 258 ],
   alphaCSR[ 50 ][ 259 ],
   alphaCSR[ 50 ][ 260 ],
   alphaCSR[ 50 ][ 261 ],
   alphaCSR[ 50 ][ 262 ],
   alphaCSR[ 50 ][ 263 ],
   alphaCSR[ 50 ][ 264 ],
   alphaCSR[ 50 ][ 265 ],
   alphaCSR[ 50 ][ 266 ],
   alphaCSR[ 50 ][ 267 ],
   alphaCSR[ 50 ][ 268 ],
   alphaCSR[ 50 ][ 269 ],
   alphaCSR[ 50 ][ 270 ],
   alphaCSR[ 50 ][ 271 ],
   alphaCSR[ 50 ][ 272 ],
   alphaCSR[ 50 ][ 273 ],
   alphaCSR[ 50 ][ 274 ],
   alphaCSR[ 50 ][ 275 ],
   alphaCSR[ 50 ][ 276 ],
   alphaCSR[ 50 ][ 277 ],
   alphaCSR[ 50 ][ 278 ],
   alphaCSR[ 50 ][ 279 ],
   alphaCSR[ 50 ][ 280 ],
   alphaCSR[ 50 ][ 281 ],
   alphaCSR[ 50 ][ 282 ],
   alphaCSR[ 50 ][ 283 ],
   alphaCSR[ 50 ][ 284 ],
   alphaCSR[ 50 ][ 285 ],
   alphaCSR[ 50 ][ 286 ],
   alphaCSR[ 50 ][ 287 ],
   alphaCSR[ 50 ][ 288 ],
   alphaCSR[ 50 ][ 289 ],
   alphaCSR[ 50 ][ 290 ],
   alphaCSR[ 50 ][ 291 ],
   alphaCSR[ 50 ][ 292 ],
   alphaCSR[ 50 ][ 293 ],
   alphaCSR[ 50 ][ 294 ],
   alphaCSR[ 50 ][ 295 ],
   alphaCSR[ 50 ][ 296 ],
   alphaCSR[ 50 ][ 297 ],
   alphaCSR[ 50 ][ 298 ],
   alphaCSR[ 50 ][ 299 ],
   alphaCSR[ 50 ][ 300 ],
   alphaCSR[ 50 ][ 301 ],
   alphaCSR[ 50 ][ 302 ],
   alphaCSR[ 50 ][ 303 ],
   alphaCSR[ 50 ][ 304 ],
   alphaCSR[ 50 ][ 305 ],
   alphaCSR[ 50 ][ 306 ],
   alphaCSR[ 50 ][ 307 ],
   alphaCSR[ 50 ][ 308 ],
   alphaCSR[ 50 ][ 309 ],
   alphaCSR[ 50 ][ 310 ],
   alphaCSR[ 50 ][ 311 ],
   alphaCSR[ 50 ][ 312 ],
   alphaCSR[ 50 ][ 313 ],
   alphaCSR[ 50 ][ 314 ],
   alphaCSR[ 50 ][ 315 ],
   alphaCSR[ 50 ][ 316 ],
   alphaCSR[ 50 ][ 317 ],
   alphaCSR[ 50 ][ 318 ],
   alphaCSR[ 50 ][ 319 ],
   alphaCSR[ 50 ][ 320 ],
   alphaCSR[ 50 ][ 321 ],
   alphaCSR[ 50 ][ 322 ],
   alphaCSR[ 50 ][ 323 ],
   alphaCSR[ 50 ][ 324 ],
   alphaCSR[ 50 ][ 325 ],
   alphaCSR[ 50 ][ 326 ],
   alphaCSR[ 50 ][ 327 ],
   alphaCSR[ 50 ][ 328 ],
   alphaCSR[ 50 ][ 329 ],
   alphaCSR[ 50 ][ 330 ],
   alphaCSR[ 50 ][ 331 ],
   alphaCSR[ 50 ][ 332 ],
   alphaCSR[ 50 ][ 333 ],
   alphaCSR[ 50 ][ 334 ],
   alphaCSR[ 50 ][ 335 ],
   alphaCSR[ 50 ][ 336 ],
   alphaCSR[ 50 ][ 337 ],
   alphaCSR[ 50 ][ 338 ],
   alphaCSR[ 50 ][ 339 ],
   alphaCSR[ 50 ][ 340 ],
   alphaCSR[ 50 ][ 341 ],
   alphaCSR[ 50 ][ 342 ],
   alphaCSR[ 50 ][ 343 ],
   alphaCSR[ 50 ][ 344 ],
   alphaCSR[ 50 ][ 345 ],
   alphaCSR[ 50 ][ 346 ],
   alphaCSR[ 50 ][ 347 ],
   alphaCSR[ 50 ][ 348 ],
   alphaCSR[ 50 ][ 349 ],
   alphaCSR[ 50 ][ 350 ],
   alphaCSR[ 50 ][ 351 ],
   alphaCSR[ 50 ][ 352 ],
   alphaCSR[ 50 ][ 353 ],
   alphaCSR[ 50 ][ 354 ],
   alphaCSR[ 50 ][ 355 ],
   alphaCSR[ 50 ][ 356 ],
   alphaCSR[ 50 ][ 357 ],
   alphaCSR[ 50 ][ 358 ],
   alphaCSR[ 50 ][ 359 ],
   alphaCSR[ 50 ][ 360 ],
   alphaCSR[ 50 ][ 361 ],
   alphaCSR[ 50 ][ 362 ],
   alphaCSR[ 50 ][ 363 ],
   alphaCSR[ 50 ][ 364 ],
   alphaCSR[ 50 ][ 365 ],
   alphaCSR[ 50 ][ 366 ],
   alphaCSR[ 50 ][ 367 ],
   alphaCSR[ 50 ][ 368 ],
   alphaCSR[ 50 ][ 369 ],
   alphaCSR[ 50 ][ 370 ],
   alphaCSR[ 50 ][ 371 ],
   alphaCSR[ 50 ][ 372 ],
   alphaCSR[ 50 ][ 373 ],
   alphaCSR[ 50 ][ 374 ],
   alphaCSR[ 50 ][ 375 ],
   alphaCSR[ 50 ][ 376 ],
   alphaCSR[ 50 ][ 377 ],
   alphaCSR[ 50 ][ 378 ],
   alphaCSR[ 50 ][ 379 ],
   alphaCSR[ 50 ][ 380 ],
   alphaCSR[ 50 ][ 381 ],
   alphaCSR[ 50 ][ 382 ],
   alphaCSR[ 50 ][ 383 ],
   alphaCSR[ 51 ][ 0 ],
   alphaCSR[ 51 ][ 1 ],
   alphaCSR[ 51 ][ 2 ],
   alphaCSR[ 51 ][ 3 ],
   alphaCSR[ 51 ][ 4 ],
   alphaCSR[ 51 ][ 5 ],
   alphaCSR[ 51 ][ 6 ],
   alphaCSR[ 51 ][ 7 ],
   alphaCSR[ 51 ][ 8 ],
   alphaCSR[ 51 ][ 9 ],
   alphaCSR[ 51 ][ 10 ],
   alphaCSR[ 51 ][ 11 ],
   alphaCSR[ 51 ][ 12 ],
   alphaCSR[ 51 ][ 13 ],
   alphaCSR[ 51 ][ 14 ],
   alphaCSR[ 51 ][ 15 ],
   alphaCSR[ 51 ][ 16 ],
   alphaCSR[ 51 ][ 17 ],
   alphaCSR[ 51 ][ 18 ],
   alphaCSR[ 51 ][ 19 ],
   alphaCSR[ 51 ][ 20 ],
   alphaCSR[ 51 ][ 21 ],
   alphaCSR[ 51 ][ 22 ],
   alphaCSR[ 51 ][ 23 ],
   alphaCSR[ 51 ][ 24 ],
   alphaCSR[ 51 ][ 25 ],
   alphaCSR[ 51 ][ 26 ],
   alphaCSR[ 51 ][ 27 ],
   alphaCSR[ 51 ][ 28 ],
   alphaCSR[ 51 ][ 29 ],
   alphaCSR[ 51 ][ 30 ],
   alphaCSR[ 51 ][ 31 ],
   alphaCSR[ 51 ][ 32 ],
   alphaCSR[ 51 ][ 33 ],
   alphaCSR[ 51 ][ 34 ],
   alphaCSR[ 51 ][ 35 ],
   alphaCSR[ 51 ][ 36 ],
   alphaCSR[ 51 ][ 37 ],
   alphaCSR[ 51 ][ 38 ],
   alphaCSR[ 51 ][ 39 ],
   alphaCSR[ 51 ][ 40 ],
   alphaCSR[ 51 ][ 41 ],
   alphaCSR[ 51 ][ 42 ],
   alphaCSR[ 51 ][ 43 ],
   alphaCSR[ 51 ][ 44 ],
   alphaCSR[ 51 ][ 45 ],
   alphaCSR[ 51 ][ 46 ],
   alphaCSR[ 51 ][ 47 ],
   alphaCSR[ 51 ][ 48 ],
   alphaCSR[ 51 ][ 49 ],
   alphaCSR[ 51 ][ 50 ],
   alphaCSR[ 51 ][ 51 ],
   alphaCSR[ 51 ][ 52 ],
   alphaCSR[ 51 ][ 53 ],
   alphaCSR[ 51 ][ 54 ],
   alphaCSR[ 51 ][ 55 ],
   alphaCSR[ 51 ][ 56 ],
   alphaCSR[ 51 ][ 57 ],
   alphaCSR[ 51 ][ 58 ],
   alphaCSR[ 51 ][ 59 ],
   alphaCSR[ 51 ][ 60 ],
   alphaCSR[ 51 ][ 61 ],
   alphaCSR[ 51 ][ 62 ],
   alphaCSR[ 51 ][ 63 ],
   alphaCSR[ 51 ][ 64 ],
   alphaCSR[ 51 ][ 65 ],
   alphaCSR[ 51 ][ 66 ],
   alphaCSR[ 51 ][ 67 ],
   alphaCSR[ 51 ][ 68 ],
   alphaCSR[ 51 ][ 69 ],
   alphaCSR[ 51 ][ 70 ],
   alphaCSR[ 51 ][ 71 ],
   alphaCSR[ 51 ][ 72 ],
   alphaCSR[ 51 ][ 73 ],
   alphaCSR[ 51 ][ 74 ],
   alphaCSR[ 51 ][ 75 ],
   alphaCSR[ 51 ][ 76 ],
   alphaCSR[ 51 ][ 77 ],
   alphaCSR[ 51 ][ 78 ],
   alphaCSR[ 51 ][ 79 ],
   alphaCSR[ 51 ][ 80 ],
   alphaCSR[ 51 ][ 81 ],
   alphaCSR[ 51 ][ 82 ],
   alphaCSR[ 51 ][ 83 ],
   alphaCSR[ 51 ][ 84 ],
   alphaCSR[ 51 ][ 85 ],
   alphaCSR[ 51 ][ 86 ],
   alphaCSR[ 51 ][ 87 ],
   alphaCSR[ 51 ][ 88 ],
   alphaCSR[ 51 ][ 89 ],
   alphaCSR[ 51 ][ 90 ],
   alphaCSR[ 51 ][ 91 ],
   alphaCSR[ 51 ][ 92 ],
   alphaCSR[ 51 ][ 93 ],
   alphaCSR[ 51 ][ 94 ],
   alphaCSR[ 51 ][ 95 ],
   alphaCSR[ 51 ][ 96 ],
   alphaCSR[ 51 ][ 97 ],
   alphaCSR[ 51 ][ 98 ],
   alphaCSR[ 51 ][ 99 ],
   alphaCSR[ 51 ][ 100 ],
   alphaCSR[ 51 ][ 101 ],
   alphaCSR[ 51 ][ 102 ],
   alphaCSR[ 51 ][ 103 ],
   alphaCSR[ 51 ][ 104 ],
   alphaCSR[ 51 ][ 105 ],
   alphaCSR[ 51 ][ 106 ],
   alphaCSR[ 51 ][ 107 ],
   alphaCSR[ 51 ][ 108 ],
   alphaCSR[ 51 ][ 109 ],
   alphaCSR[ 51 ][ 110 ],
   alphaCSR[ 51 ][ 111 ],
   alphaCSR[ 51 ][ 112 ],
   alphaCSR[ 51 ][ 113 ],
   alphaCSR[ 51 ][ 114 ],
   alphaCSR[ 51 ][ 115 ],
   alphaCSR[ 51 ][ 116 ],
   alphaCSR[ 51 ][ 117 ],
   alphaCSR[ 51 ][ 118 ],
   alphaCSR[ 51 ][ 119 ],
   alphaCSR[ 51 ][ 120 ],
   alphaCSR[ 51 ][ 121 ],
   alphaCSR[ 51 ][ 122 ],
   alphaCSR[ 51 ][ 123 ],
   alphaCSR[ 51 ][ 124 ],
   alphaCSR[ 51 ][ 125 ],
   alphaCSR[ 51 ][ 126 ],
   alphaCSR[ 51 ][ 127 ],
   alphaCSR[ 51 ][ 128 ],
   alphaCSR[ 51 ][ 129 ],
   alphaCSR[ 51 ][ 130 ],
   alphaCSR[ 51 ][ 131 ],
   alphaCSR[ 51 ][ 132 ],
   alphaCSR[ 51 ][ 133 ],
   alphaCSR[ 51 ][ 134 ],
   alphaCSR[ 51 ][ 135 ],
   alphaCSR[ 51 ][ 136 ],
   alphaCSR[ 51 ][ 137 ],
   alphaCSR[ 51 ][ 138 ],
   alphaCSR[ 51 ][ 139 ],
   alphaCSR[ 51 ][ 140 ],
   alphaCSR[ 51 ][ 141 ],
   alphaCSR[ 51 ][ 142 ],
   alphaCSR[ 51 ][ 143 ],
   alphaCSR[ 51 ][ 144 ],
   alphaCSR[ 51 ][ 145 ],
   alphaCSR[ 51 ][ 146 ],
   alphaCSR[ 51 ][ 147 ],
   alphaCSR[ 51 ][ 148 ],
   alphaCSR[ 51 ][ 149 ],
   alphaCSR[ 51 ][ 150 ],
   alphaCSR[ 51 ][ 151 ],
   alphaCSR[ 51 ][ 152 ],
   alphaCSR[ 51 ][ 153 ],
   alphaCSR[ 51 ][ 154 ],
   alphaCSR[ 51 ][ 155 ],
   alphaCSR[ 51 ][ 156 ],
   alphaCSR[ 51 ][ 157 ],
   alphaCSR[ 51 ][ 158 ],
   alphaCSR[ 51 ][ 159 ],
   alphaCSR[ 51 ][ 160 ],
   alphaCSR[ 51 ][ 161 ],
   alphaCSR[ 51 ][ 162 ],
   alphaCSR[ 51 ][ 163 ],
   alphaCSR[ 51 ][ 164 ],
   alphaCSR[ 51 ][ 165 ],
   alphaCSR[ 51 ][ 166 ],
   alphaCSR[ 51 ][ 167 ],
   alphaCSR[ 51 ][ 168 ],
   alphaCSR[ 51 ][ 169 ],
   alphaCSR[ 51 ][ 170 ],
   alphaCSR[ 51 ][ 171 ],
   alphaCSR[ 51 ][ 172 ],
   alphaCSR[ 51 ][ 173 ],
   alphaCSR[ 51 ][ 174 ],
   alphaCSR[ 51 ][ 175 ],
   alphaCSR[ 51 ][ 176 ],
   alphaCSR[ 51 ][ 177 ],
   alphaCSR[ 51 ][ 178 ],
   alphaCSR[ 51 ][ 179 ],
   alphaCSR[ 51 ][ 180 ],
   alphaCSR[ 51 ][ 181 ],
   alphaCSR[ 51 ][ 182 ],
   alphaCSR[ 51 ][ 183 ],
   alphaCSR[ 51 ][ 184 ],
   alphaCSR[ 51 ][ 185 ],
   alphaCSR[ 51 ][ 186 ],
   alphaCSR[ 51 ][ 187 ],
   alphaCSR[ 51 ][ 188 ],
   alphaCSR[ 51 ][ 189 ],
   alphaCSR[ 51 ][ 190 ],
   alphaCSR[ 51 ][ 191 ],
   alphaCSR[ 51 ][ 192 ],
   alphaCSR[ 51 ][ 193 ],
   alphaCSR[ 51 ][ 194 ],
   alphaCSR[ 51 ][ 195 ],
   alphaCSR[ 51 ][ 196 ],
   alphaCSR[ 51 ][ 197 ],
   alphaCSR[ 51 ][ 198 ],
   alphaCSR[ 51 ][ 199 ],
   alphaCSR[ 51 ][ 200 ],
   alphaCSR[ 51 ][ 201 ],
   alphaCSR[ 51 ][ 202 ],
   alphaCSR[ 51 ][ 203 ],
   alphaCSR[ 51 ][ 204 ],
   alphaCSR[ 51 ][ 205 ],
   alphaCSR[ 51 ][ 206 ],
   alphaCSR[ 51 ][ 207 ],
   alphaCSR[ 51 ][ 208 ],
   alphaCSR[ 51 ][ 209 ],
   alphaCSR[ 51 ][ 210 ],
   alphaCSR[ 51 ][ 211 ],
   alphaCSR[ 51 ][ 212 ],
   alphaCSR[ 51 ][ 213 ],
   alphaCSR[ 51 ][ 214 ],
   alphaCSR[ 51 ][ 215 ],
   alphaCSR[ 51 ][ 216 ],
   alphaCSR[ 51 ][ 217 ],
   alphaCSR[ 51 ][ 218 ],
   alphaCSR[ 51 ][ 219 ],
   alphaCSR[ 51 ][ 220 ],
   alphaCSR[ 51 ][ 221 ],
   alphaCSR[ 51 ][ 222 ],
   alphaCSR[ 51 ][ 223 ],
   alphaCSR[ 51 ][ 224 ],
   alphaCSR[ 51 ][ 225 ],
   alphaCSR[ 51 ][ 226 ],
   alphaCSR[ 51 ][ 227 ],
   alphaCSR[ 51 ][ 228 ],
   alphaCSR[ 51 ][ 229 ],
   alphaCSR[ 51 ][ 230 ],
   alphaCSR[ 51 ][ 231 ],
   alphaCSR[ 51 ][ 232 ],
   alphaCSR[ 51 ][ 233 ],
   alphaCSR[ 51 ][ 234 ],
   alphaCSR[ 51 ][ 235 ],
   alphaCSR[ 51 ][ 236 ],
   alphaCSR[ 51 ][ 237 ],
   alphaCSR[ 51 ][ 238 ],
   alphaCSR[ 51 ][ 239 ],
   alphaCSR[ 51 ][ 240 ],
   alphaCSR[ 51 ][ 241 ],
   alphaCSR[ 51 ][ 242 ],
   alphaCSR[ 51 ][ 243 ],
   alphaCSR[ 51 ][ 244 ],
   alphaCSR[ 51 ][ 245 ],
   alphaCSR[ 51 ][ 246 ],
   alphaCSR[ 51 ][ 247 ],
   alphaCSR[ 51 ][ 248 ],
   alphaCSR[ 51 ][ 249 ],
   alphaCSR[ 51 ][ 250 ],
   alphaCSR[ 51 ][ 251 ],
   alphaCSR[ 51 ][ 252 ],
   alphaCSR[ 51 ][ 253 ],
   alphaCSR[ 51 ][ 254 ],
   alphaCSR[ 51 ][ 255 ],
   alphaCSR[ 51 ][ 256 ],
   alphaCSR[ 51 ][ 257 ],
   alphaCSR[ 51 ][ 258 ],
   alphaCSR[ 51 ][ 259 ],
   alphaCSR[ 51 ][ 260 ],
   alphaCSR[ 51 ][ 261 ],
   alphaCSR[ 51 ][ 262 ],
   alphaCSR[ 51 ][ 263 ],
   alphaCSR[ 51 ][ 264 ],
   alphaCSR[ 51 ][ 265 ],
   alphaCSR[ 51 ][ 266 ],
   alphaCSR[ 51 ][ 267 ],
   alphaCSR[ 51 ][ 268 ],
   alphaCSR[ 51 ][ 269 ],
   alphaCSR[ 51 ][ 270 ],
   alphaCSR[ 51 ][ 271 ],
   alphaCSR[ 51 ][ 272 ],
   alphaCSR[ 51 ][ 273 ],
   alphaCSR[ 51 ][ 274 ],
   alphaCSR[ 51 ][ 275 ],
   alphaCSR[ 51 ][ 276 ],
   alphaCSR[ 51 ][ 277 ],
   alphaCSR[ 51 ][ 278 ],
   alphaCSR[ 51 ][ 279 ],
   alphaCSR[ 51 ][ 280 ],
   alphaCSR[ 51 ][ 281 ],
   alphaCSR[ 51 ][ 282 ],
   alphaCSR[ 51 ][ 283 ],
   alphaCSR[ 51 ][ 284 ],
   alphaCSR[ 51 ][ 285 ],
   alphaCSR[ 51 ][ 286 ],
   alphaCSR[ 51 ][ 287 ],
   alphaCSR[ 51 ][ 288 ],
   alphaCSR[ 51 ][ 289 ],
   alphaCSR[ 51 ][ 290 ],
   alphaCSR[ 51 ][ 291 ],
   alphaCSR[ 51 ][ 292 ],
   alphaCSR[ 51 ][ 293 ],
   alphaCSR[ 51 ][ 294 ],
   alphaCSR[ 51 ][ 295 ],
   alphaCSR[ 51 ][ 296 ],
   alphaCSR[ 51 ][ 297 ],
   alphaCSR[ 51 ][ 298 ],
   alphaCSR[ 51 ][ 299 ],
   alphaCSR[ 51 ][ 300 ],
   alphaCSR[ 51 ][ 301 ],
   alphaCSR[ 51 ][ 302 ],
   alphaCSR[ 51 ][ 303 ],
   alphaCSR[ 51 ][ 304 ],
   alphaCSR[ 51 ][ 305 ],
   alphaCSR[ 51 ][ 306 ],
   alphaCSR[ 51 ][ 307 ],
   alphaCSR[ 51 ][ 308 ],
   alphaCSR[ 51 ][ 309 ],
   alphaCSR[ 51 ][ 310 ],
   alphaCSR[ 51 ][ 311 ],
   alphaCSR[ 51 ][ 312 ],
   alphaCSR[ 51 ][ 313 ],
   alphaCSR[ 51 ][ 314 ],
   alphaCSR[ 51 ][ 315 ],
   alphaCSR[ 51 ][ 316 ],
   alphaCSR[ 51 ][ 317 ],
   alphaCSR[ 51 ][ 318 ],
   alphaCSR[ 51 ][ 319 ],
   alphaCSR[ 51 ][ 320 ],
   alphaCSR[ 51 ][ 321 ],
   alphaCSR[ 51 ][ 322 ],
   alphaCSR[ 51 ][ 323 ],
   alphaCSR[ 51 ][ 324 ],
   alphaCSR[ 51 ][ 325 ],
   alphaCSR[ 51 ][ 326 ],
   alphaCSR[ 51 ][ 327 ],
   alphaCSR[ 51 ][ 328 ],
   alphaCSR[ 51 ][ 329 ],
   alphaCSR[ 51 ][ 330 ],
   alphaCSR[ 51 ][ 331 ],
   alphaCSR[ 51 ][ 332 ],
   alphaCSR[ 51 ][ 333 ],
   alphaCSR[ 51 ][ 334 ],
   alphaCSR[ 51 ][ 335 ],
   alphaCSR[ 51 ][ 336 ],
   alphaCSR[ 51 ][ 337 ],
   alphaCSR[ 51 ][ 338 ],
   alphaCSR[ 51 ][ 339 ],
   alphaCSR[ 51 ][ 340 ],
   alphaCSR[ 51 ][ 341 ],
   alphaCSR[ 51 ][ 342 ],
   alphaCSR[ 51 ][ 343 ],
   alphaCSR[ 51 ][ 344 ],
   alphaCSR[ 51 ][ 345 ],
   alphaCSR[ 51 ][ 346 ],
   alphaCSR[ 51 ][ 347 ],
   alphaCSR[ 51 ][ 348 ],
   alphaCSR[ 51 ][ 349 ],
   alphaCSR[ 51 ][ 350 ],
   alphaCSR[ 51 ][ 351 ],
   alphaCSR[ 51 ][ 352 ],
   alphaCSR[ 51 ][ 353 ],
   alphaCSR[ 51 ][ 354 ],
   alphaCSR[ 51 ][ 355 ],
   alphaCSR[ 51 ][ 356 ],
   alphaCSR[ 51 ][ 357 ],
   alphaCSR[ 51 ][ 358 ],
   alphaCSR[ 51 ][ 359 ],
   alphaCSR[ 51 ][ 360 ],
   alphaCSR[ 51 ][ 361 ],
   alphaCSR[ 51 ][ 362 ],
   alphaCSR[ 51 ][ 363 ],
   alphaCSR[ 51 ][ 364 ],
   alphaCSR[ 51 ][ 365 ],
   alphaCSR[ 51 ][ 366 ],
   alphaCSR[ 51 ][ 367 ],
   alphaCSR[ 51 ][ 368 ],
   alphaCSR[ 51 ][ 369 ],
   alphaCSR[ 51 ][ 370 ],
   alphaCSR[ 51 ][ 371 ],
   alphaCSR[ 51 ][ 372 ],
   alphaCSR[ 51 ][ 373 ],
   alphaCSR[ 51 ][ 374 ],
   alphaCSR[ 51 ][ 375 ],
   alphaCSR[ 51 ][ 376 ],
   alphaCSR[ 51 ][ 377 ],
   alphaCSR[ 51 ][ 378 ],
   alphaCSR[ 51 ][ 379 ],
   alphaCSR[ 51 ][ 380 ],
   alphaCSR[ 51 ][ 381 ],
   alphaCSR[ 51 ][ 382 ],
   alphaCSR[ 51 ][ 383 ],
   alphaCSR[ 52 ][ 0 ],
   alphaCSR[ 52 ][ 1 ],
   alphaCSR[ 52 ][ 2 ],
   alphaCSR[ 52 ][ 3 ],
   alphaCSR[ 52 ][ 4 ],
   alphaCSR[ 52 ][ 5 ],
   alphaCSR[ 52 ][ 6 ],
   alphaCSR[ 52 ][ 7 ],
   alphaCSR[ 52 ][ 8 ],
   alphaCSR[ 52 ][ 9 ],
   alphaCSR[ 52 ][ 10 ],
   alphaCSR[ 52 ][ 11 ],
   alphaCSR[ 52 ][ 12 ],
   alphaCSR[ 52 ][ 13 ],
   alphaCSR[ 52 ][ 14 ],
   alphaCSR[ 52 ][ 15 ],
   alphaCSR[ 52 ][ 16 ],
   alphaCSR[ 52 ][ 17 ],
   alphaCSR[ 52 ][ 18 ],
   alphaCSR[ 52 ][ 19 ],
   alphaCSR[ 52 ][ 20 ],
   alphaCSR[ 52 ][ 21 ],
   alphaCSR[ 52 ][ 22 ],
   alphaCSR[ 52 ][ 23 ],
   alphaCSR[ 52 ][ 24 ],
   alphaCSR[ 52 ][ 25 ],
   alphaCSR[ 52 ][ 26 ],
   alphaCSR[ 52 ][ 27 ],
   alphaCSR[ 52 ][ 28 ],
   alphaCSR[ 52 ][ 29 ],
   alphaCSR[ 52 ][ 30 ],
   alphaCSR[ 52 ][ 31 ],
   alphaCSR[ 52 ][ 32 ],
   alphaCSR[ 52 ][ 33 ],
   alphaCSR[ 52 ][ 34 ],
   alphaCSR[ 52 ][ 35 ],
   alphaCSR[ 52 ][ 36 ],
   alphaCSR[ 52 ][ 37 ],
   alphaCSR[ 52 ][ 38 ],
   alphaCSR[ 52 ][ 39 ],
   alphaCSR[ 52 ][ 40 ],
   alphaCSR[ 52 ][ 41 ],
   alphaCSR[ 52 ][ 42 ],
   alphaCSR[ 52 ][ 43 ],
   alphaCSR[ 52 ][ 44 ],
   alphaCSR[ 52 ][ 45 ],
   alphaCSR[ 52 ][ 46 ],
   alphaCSR[ 52 ][ 47 ],
   alphaCSR[ 52 ][ 48 ],
   alphaCSR[ 52 ][ 49 ],
   alphaCSR[ 52 ][ 50 ],
   alphaCSR[ 52 ][ 51 ],
   alphaCSR[ 52 ][ 52 ],
   alphaCSR[ 52 ][ 53 ],
   alphaCSR[ 52 ][ 54 ],
   alphaCSR[ 52 ][ 55 ],
   alphaCSR[ 52 ][ 56 ],
   alphaCSR[ 52 ][ 57 ],
   alphaCSR[ 52 ][ 58 ],
   alphaCSR[ 52 ][ 59 ],
   alphaCSR[ 52 ][ 60 ],
   alphaCSR[ 52 ][ 61 ],
   alphaCSR[ 52 ][ 62 ],
   alphaCSR[ 52 ][ 63 ],
   alphaCSR[ 52 ][ 64 ],
   alphaCSR[ 52 ][ 65 ],
   alphaCSR[ 52 ][ 66 ],
   alphaCSR[ 52 ][ 67 ],
   alphaCSR[ 52 ][ 68 ],
   alphaCSR[ 52 ][ 69 ],
   alphaCSR[ 52 ][ 70 ],
   alphaCSR[ 52 ][ 71 ],
   alphaCSR[ 52 ][ 72 ],
   alphaCSR[ 52 ][ 73 ],
   alphaCSR[ 52 ][ 74 ],
   alphaCSR[ 52 ][ 75 ],
   alphaCSR[ 52 ][ 76 ],
   alphaCSR[ 52 ][ 77 ],
   alphaCSR[ 52 ][ 78 ],
   alphaCSR[ 52 ][ 79 ],
   alphaCSR[ 52 ][ 80 ],
   alphaCSR[ 52 ][ 81 ],
   alphaCSR[ 52 ][ 82 ],
   alphaCSR[ 52 ][ 83 ],
   alphaCSR[ 52 ][ 84 ],
   alphaCSR[ 52 ][ 85 ],
   alphaCSR[ 52 ][ 86 ],
   alphaCSR[ 52 ][ 87 ],
   alphaCSR[ 52 ][ 88 ],
   alphaCSR[ 52 ][ 89 ],
   alphaCSR[ 52 ][ 90 ],
   alphaCSR[ 52 ][ 91 ],
   alphaCSR[ 52 ][ 92 ],
   alphaCSR[ 52 ][ 93 ],
   alphaCSR[ 52 ][ 94 ],
   alphaCSR[ 52 ][ 95 ],
   alphaCSR[ 52 ][ 96 ],
   alphaCSR[ 52 ][ 97 ],
   alphaCSR[ 52 ][ 98 ],
   alphaCSR[ 52 ][ 99 ],
   alphaCSR[ 52 ][ 100 ],
   alphaCSR[ 52 ][ 101 ],
   alphaCSR[ 52 ][ 102 ],
   alphaCSR[ 52 ][ 103 ],
   alphaCSR[ 52 ][ 104 ],
   alphaCSR[ 52 ][ 105 ],
   alphaCSR[ 52 ][ 106 ],
   alphaCSR[ 52 ][ 107 ],
   alphaCSR[ 52 ][ 108 ],
   alphaCSR[ 52 ][ 109 ],
   alphaCSR[ 52 ][ 110 ],
   alphaCSR[ 52 ][ 111 ],
   alphaCSR[ 52 ][ 112 ],
   alphaCSR[ 52 ][ 113 ],
   alphaCSR[ 52 ][ 114 ],
   alphaCSR[ 52 ][ 115 ],
   alphaCSR[ 52 ][ 116 ],
   alphaCSR[ 52 ][ 117 ],
   alphaCSR[ 52 ][ 118 ],
   alphaCSR[ 52 ][ 119 ],
   alphaCSR[ 52 ][ 120 ],
   alphaCSR[ 52 ][ 121 ],
   alphaCSR[ 52 ][ 122 ],
   alphaCSR[ 52 ][ 123 ],
   alphaCSR[ 52 ][ 124 ],
   alphaCSR[ 52 ][ 125 ],
   alphaCSR[ 52 ][ 126 ],
   alphaCSR[ 52 ][ 127 ],
   alphaCSR[ 52 ][ 128 ],
   alphaCSR[ 52 ][ 129 ],
   alphaCSR[ 52 ][ 130 ],
   alphaCSR[ 52 ][ 131 ],
   alphaCSR[ 52 ][ 132 ],
   alphaCSR[ 52 ][ 133 ],
   alphaCSR[ 52 ][ 134 ],
   alphaCSR[ 52 ][ 135 ],
   alphaCSR[ 52 ][ 136 ],
   alphaCSR[ 52 ][ 137 ],
   alphaCSR[ 52 ][ 138 ],
   alphaCSR[ 52 ][ 139 ],
   alphaCSR[ 52 ][ 140 ],
   alphaCSR[ 52 ][ 141 ],
   alphaCSR[ 52 ][ 142 ],
   alphaCSR[ 52 ][ 143 ],
   alphaCSR[ 52 ][ 144 ],
   alphaCSR[ 52 ][ 145 ],
   alphaCSR[ 52 ][ 146 ],
   alphaCSR[ 52 ][ 147 ],
   alphaCSR[ 52 ][ 148 ],
   alphaCSR[ 52 ][ 149 ],
   alphaCSR[ 52 ][ 150 ],
   alphaCSR[ 52 ][ 151 ],
   alphaCSR[ 52 ][ 152 ],
   alphaCSR[ 52 ][ 153 ],
   alphaCSR[ 52 ][ 154 ],
   alphaCSR[ 52 ][ 155 ],
   alphaCSR[ 52 ][ 156 ],
   alphaCSR[ 52 ][ 157 ],
   alphaCSR[ 52 ][ 158 ],
   alphaCSR[ 52 ][ 159 ],
   alphaCSR[ 52 ][ 160 ],
   alphaCSR[ 52 ][ 161 ],
   alphaCSR[ 52 ][ 162 ],
   alphaCSR[ 52 ][ 163 ],
   alphaCSR[ 52 ][ 164 ],
   alphaCSR[ 52 ][ 165 ],
   alphaCSR[ 52 ][ 166 ],
   alphaCSR[ 52 ][ 167 ],
   alphaCSR[ 52 ][ 168 ],
   alphaCSR[ 52 ][ 169 ],
   alphaCSR[ 52 ][ 170 ],
   alphaCSR[ 52 ][ 171 ],
   alphaCSR[ 52 ][ 172 ],
   alphaCSR[ 52 ][ 173 ],
   alphaCSR[ 52 ][ 174 ],
   alphaCSR[ 52 ][ 175 ],
   alphaCSR[ 52 ][ 176 ],
   alphaCSR[ 52 ][ 177 ],
   alphaCSR[ 52 ][ 178 ],
   alphaCSR[ 52 ][ 179 ],
   alphaCSR[ 52 ][ 180 ],
   alphaCSR[ 52 ][ 181 ],
   alphaCSR[ 52 ][ 182 ],
   alphaCSR[ 52 ][ 183 ],
   alphaCSR[ 52 ][ 184 ],
   alphaCSR[ 52 ][ 185 ],
   alphaCSR[ 52 ][ 186 ],
   alphaCSR[ 52 ][ 187 ],
   alphaCSR[ 52 ][ 188 ],
   alphaCSR[ 52 ][ 189 ],
   alphaCSR[ 52 ][ 190 ],
   alphaCSR[ 52 ][ 191 ],
   alphaCSR[ 52 ][ 192 ],
   alphaCSR[ 52 ][ 193 ],
   alphaCSR[ 52 ][ 194 ],
   alphaCSR[ 52 ][ 195 ],
   alphaCSR[ 52 ][ 196 ],
   alphaCSR[ 52 ][ 197 ],
   alphaCSR[ 52 ][ 198 ],
   alphaCSR[ 52 ][ 199 ],
   alphaCSR[ 52 ][ 200 ],
   alphaCSR[ 52 ][ 201 ],
   alphaCSR[ 52 ][ 202 ],
   alphaCSR[ 52 ][ 203 ],
   alphaCSR[ 52 ][ 204 ],
   alphaCSR[ 52 ][ 205 ],
   alphaCSR[ 52 ][ 206 ],
   alphaCSR[ 52 ][ 207 ],
   alphaCSR[ 52 ][ 208 ],
   alphaCSR[ 52 ][ 209 ],
   alphaCSR[ 52 ][ 210 ],
   alphaCSR[ 52 ][ 211 ],
   alphaCSR[ 52 ][ 212 ],
   alphaCSR[ 52 ][ 213 ],
   alphaCSR[ 52 ][ 214 ],
   alphaCSR[ 52 ][ 215 ],
   alphaCSR[ 52 ][ 216 ],
   alphaCSR[ 52 ][ 217 ],
   alphaCSR[ 52 ][ 218 ],
   alphaCSR[ 52 ][ 219 ],
   alphaCSR[ 52 ][ 220 ],
   alphaCSR[ 52 ][ 221 ],
   alphaCSR[ 52 ][ 222 ],
   alphaCSR[ 52 ][ 223 ],
   alphaCSR[ 52 ][ 224 ],
   alphaCSR[ 52 ][ 225 ],
   alphaCSR[ 52 ][ 226 ],
   alphaCSR[ 52 ][ 227 ],
   alphaCSR[ 52 ][ 228 ],
   alphaCSR[ 52 ][ 229 ],
   alphaCSR[ 52 ][ 230 ],
   alphaCSR[ 52 ][ 231 ],
   alphaCSR[ 52 ][ 232 ],
   alphaCSR[ 52 ][ 233 ],
   alphaCSR[ 52 ][ 234 ],
   alphaCSR[ 52 ][ 235 ],
   alphaCSR[ 52 ][ 236 ],
   alphaCSR[ 52 ][ 237 ],
   alphaCSR[ 52 ][ 238 ],
   alphaCSR[ 52 ][ 239 ],
   alphaCSR[ 52 ][ 240 ],
   alphaCSR[ 52 ][ 241 ],
   alphaCSR[ 52 ][ 242 ],
   alphaCSR[ 52 ][ 243 ],
   alphaCSR[ 52 ][ 244 ],
   alphaCSR[ 52 ][ 245 ],
   alphaCSR[ 52 ][ 246 ],
   alphaCSR[ 52 ][ 247 ],
   alphaCSR[ 52 ][ 248 ],
   alphaCSR[ 52 ][ 249 ],
   alphaCSR[ 52 ][ 250 ],
   alphaCSR[ 52 ][ 251 ],
   alphaCSR[ 52 ][ 252 ],
   alphaCSR[ 52 ][ 253 ],
   alphaCSR[ 52 ][ 254 ],
   alphaCSR[ 52 ][ 255 ],
   alphaCSR[ 52 ][ 256 ],
   alphaCSR[ 52 ][ 257 ],
   alphaCSR[ 52 ][ 258 ],
   alphaCSR[ 52 ][ 259 ],
   alphaCSR[ 52 ][ 260 ],
   alphaCSR[ 52 ][ 261 ],
   alphaCSR[ 52 ][ 262 ],
   alphaCSR[ 52 ][ 263 ],
   alphaCSR[ 52 ][ 264 ],
   alphaCSR[ 52 ][ 265 ],
   alphaCSR[ 52 ][ 266 ],
   alphaCSR[ 52 ][ 267 ],
   alphaCSR[ 52 ][ 268 ],
   alphaCSR[ 52 ][ 269 ],
   alphaCSR[ 52 ][ 270 ],
   alphaCSR[ 52 ][ 271 ],
   alphaCSR[ 52 ][ 272 ],
   alphaCSR[ 52 ][ 273 ],
   alphaCSR[ 52 ][ 274 ],
   alphaCSR[ 52 ][ 275 ],
   alphaCSR[ 52 ][ 276 ],
   alphaCSR[ 52 ][ 277 ],
   alphaCSR[ 52 ][ 278 ],
   alphaCSR[ 52 ][ 279 ],
   alphaCSR[ 52 ][ 280 ],
   alphaCSR[ 52 ][ 281 ],
   alphaCSR[ 52 ][ 282 ],
   alphaCSR[ 52 ][ 283 ],
   alphaCSR[ 52 ][ 284 ],
   alphaCSR[ 52 ][ 285 ],
   alphaCSR[ 52 ][ 286 ],
   alphaCSR[ 52 ][ 287 ],
   alphaCSR[ 52 ][ 288 ],
   alphaCSR[ 52 ][ 289 ],
   alphaCSR[ 52 ][ 290 ],
   alphaCSR[ 52 ][ 291 ],
   alphaCSR[ 52 ][ 292 ],
   alphaCSR[ 52 ][ 293 ],
   alphaCSR[ 52 ][ 294 ],
   alphaCSR[ 52 ][ 295 ],
   alphaCSR[ 52 ][ 296 ],
   alphaCSR[ 52 ][ 297 ],
   alphaCSR[ 52 ][ 298 ],
   alphaCSR[ 52 ][ 299 ],
   alphaCSR[ 52 ][ 300 ],
   alphaCSR[ 52 ][ 301 ],
   alphaCSR[ 52 ][ 302 ],
   alphaCSR[ 52 ][ 303 ],
   alphaCSR[ 52 ][ 304 ],
   alphaCSR[ 52 ][ 305 ],
   alphaCSR[ 52 ][ 306 ],
   alphaCSR[ 52 ][ 307 ],
   alphaCSR[ 52 ][ 308 ],
   alphaCSR[ 52 ][ 309 ],
   alphaCSR[ 52 ][ 310 ],
   alphaCSR[ 52 ][ 311 ],
   alphaCSR[ 52 ][ 312 ],
   alphaCSR[ 52 ][ 313 ],
   alphaCSR[ 52 ][ 314 ],
   alphaCSR[ 52 ][ 315 ],
   alphaCSR[ 52 ][ 316 ],
   alphaCSR[ 52 ][ 317 ],
   alphaCSR[ 52 ][ 318 ],
   alphaCSR[ 52 ][ 319 ],
   alphaCSR[ 52 ][ 320 ],
   alphaCSR[ 52 ][ 321 ],
   alphaCSR[ 52 ][ 322 ],
   alphaCSR[ 52 ][ 323 ],
   alphaCSR[ 52 ][ 324 ],
   alphaCSR[ 52 ][ 325 ],
   alphaCSR[ 52 ][ 326 ],
   alphaCSR[ 52 ][ 327 ],
   alphaCSR[ 52 ][ 328 ],
   alphaCSR[ 52 ][ 329 ],
   alphaCSR[ 52 ][ 330 ],
   alphaCSR[ 52 ][ 331 ],
   alphaCSR[ 52 ][ 332 ],
   alphaCSR[ 52 ][ 333 ],
   alphaCSR[ 52 ][ 334 ],
   alphaCSR[ 52 ][ 335 ],
   alphaCSR[ 52 ][ 336 ],
   alphaCSR[ 52 ][ 337 ],
   alphaCSR[ 52 ][ 338 ],
   alphaCSR[ 52 ][ 339 ],
   alphaCSR[ 52 ][ 340 ],
   alphaCSR[ 52 ][ 341 ],
   alphaCSR[ 52 ][ 342 ],
   alphaCSR[ 52 ][ 343 ],
   alphaCSR[ 52 ][ 344 ],
   alphaCSR[ 52 ][ 345 ],
   alphaCSR[ 52 ][ 346 ],
   alphaCSR[ 52 ][ 347 ],
   alphaCSR[ 52 ][ 348 ],
   alphaCSR[ 52 ][ 349 ],
   alphaCSR[ 52 ][ 350 ],
   alphaCSR[ 52 ][ 351 ],
   alphaCSR[ 52 ][ 352 ],
   alphaCSR[ 52 ][ 353 ],
   alphaCSR[ 52 ][ 354 ],
   alphaCSR[ 52 ][ 355 ],
   alphaCSR[ 52 ][ 356 ],
   alphaCSR[ 52 ][ 357 ],
   alphaCSR[ 52 ][ 358 ],
   alphaCSR[ 52 ][ 359 ],
   alphaCSR[ 52 ][ 360 ],
   alphaCSR[ 52 ][ 361 ],
   alphaCSR[ 52 ][ 362 ],
   alphaCSR[ 52 ][ 363 ],
   alphaCSR[ 52 ][ 364 ],
   alphaCSR[ 52 ][ 365 ],
   alphaCSR[ 52 ][ 366 ],
   alphaCSR[ 52 ][ 367 ],
   alphaCSR[ 52 ][ 368 ],
   alphaCSR[ 52 ][ 369 ],
   alphaCSR[ 52 ][ 370 ],
   alphaCSR[ 52 ][ 371 ],
   alphaCSR[ 52 ][ 372 ],
   alphaCSR[ 52 ][ 373 ],
   alphaCSR[ 52 ][ 374 ],
   alphaCSR[ 52 ][ 375 ],
   alphaCSR[ 52 ][ 376 ],
   alphaCSR[ 52 ][ 377 ],
   alphaCSR[ 52 ][ 378 ],
   alphaCSR[ 52 ][ 379 ],
   alphaCSR[ 52 ][ 380 ],
   alphaCSR[ 52 ][ 381 ],
   alphaCSR[ 52 ][ 382 ],
   alphaCSR[ 52 ][ 383 ],
   alphaCSR[ 53 ][ 0 ],
   alphaCSR[ 53 ][ 1 ],
   alphaCSR[ 53 ][ 2 ],
   alphaCSR[ 53 ][ 3 ],
   alphaCSR[ 53 ][ 4 ],
   alphaCSR[ 53 ][ 5 ],
   alphaCSR[ 53 ][ 6 ],
   alphaCSR[ 53 ][ 7 ],
   alphaCSR[ 53 ][ 8 ],
   alphaCSR[ 53 ][ 9 ],
   alphaCSR[ 53 ][ 10 ],
   alphaCSR[ 53 ][ 11 ],
   alphaCSR[ 53 ][ 12 ],
   alphaCSR[ 53 ][ 13 ],
   alphaCSR[ 53 ][ 14 ],
   alphaCSR[ 53 ][ 15 ],
   alphaCSR[ 53 ][ 16 ],
   alphaCSR[ 53 ][ 17 ],
   alphaCSR[ 53 ][ 18 ],
   alphaCSR[ 53 ][ 19 ],
   alphaCSR[ 53 ][ 20 ],
   alphaCSR[ 53 ][ 21 ],
   alphaCSR[ 53 ][ 22 ],
   alphaCSR[ 53 ][ 23 ],
   alphaCSR[ 53 ][ 24 ],
   alphaCSR[ 53 ][ 25 ],
   alphaCSR[ 53 ][ 26 ],
   alphaCSR[ 53 ][ 27 ],
   alphaCSR[ 53 ][ 28 ],
   alphaCSR[ 53 ][ 29 ],
   alphaCSR[ 53 ][ 30 ],
   alphaCSR[ 53 ][ 31 ],
   alphaCSR[ 53 ][ 32 ],
   alphaCSR[ 53 ][ 33 ],
   alphaCSR[ 53 ][ 34 ],
   alphaCSR[ 53 ][ 35 ],
   alphaCSR[ 53 ][ 36 ],
   alphaCSR[ 53 ][ 37 ],
   alphaCSR[ 53 ][ 38 ],
   alphaCSR[ 53 ][ 39 ],
   alphaCSR[ 53 ][ 40 ],
   alphaCSR[ 53 ][ 41 ],
   alphaCSR[ 53 ][ 42 ],
   alphaCSR[ 53 ][ 43 ],
   alphaCSR[ 53 ][ 44 ],
   alphaCSR[ 53 ][ 45 ],
   alphaCSR[ 53 ][ 46 ],
   alphaCSR[ 53 ][ 47 ],
   alphaCSR[ 53 ][ 48 ],
   alphaCSR[ 53 ][ 49 ],
   alphaCSR[ 53 ][ 50 ],
   alphaCSR[ 53 ][ 51 ],
   alphaCSR[ 53 ][ 52 ],
   alphaCSR[ 53 ][ 53 ],
   alphaCSR[ 53 ][ 54 ],
   alphaCSR[ 53 ][ 55 ],
   alphaCSR[ 53 ][ 56 ],
   alphaCSR[ 53 ][ 57 ],
   alphaCSR[ 53 ][ 58 ],
   alphaCSR[ 53 ][ 59 ],
   alphaCSR[ 53 ][ 60 ],
   alphaCSR[ 53 ][ 61 ],
   alphaCSR[ 53 ][ 62 ],
   alphaCSR[ 53 ][ 63 ],
   alphaCSR[ 53 ][ 64 ],
   alphaCSR[ 53 ][ 65 ],
   alphaCSR[ 53 ][ 66 ],
   alphaCSR[ 53 ][ 67 ],
   alphaCSR[ 53 ][ 68 ],
   alphaCSR[ 53 ][ 69 ],
   alphaCSR[ 53 ][ 70 ],
   alphaCSR[ 53 ][ 71 ],
   alphaCSR[ 53 ][ 72 ],
   alphaCSR[ 53 ][ 73 ],
   alphaCSR[ 53 ][ 74 ],
   alphaCSR[ 53 ][ 75 ],
   alphaCSR[ 53 ][ 76 ],
   alphaCSR[ 53 ][ 77 ],
   alphaCSR[ 53 ][ 78 ],
   alphaCSR[ 53 ][ 79 ],
   alphaCSR[ 53 ][ 80 ],
   alphaCSR[ 53 ][ 81 ],
   alphaCSR[ 53 ][ 82 ],
   alphaCSR[ 53 ][ 83 ],
   alphaCSR[ 53 ][ 84 ],
   alphaCSR[ 53 ][ 85 ],
   alphaCSR[ 53 ][ 86 ],
   alphaCSR[ 53 ][ 87 ],
   alphaCSR[ 53 ][ 88 ],
   alphaCSR[ 53 ][ 89 ],
   alphaCSR[ 53 ][ 90 ],
   alphaCSR[ 53 ][ 91 ],
   alphaCSR[ 53 ][ 92 ],
   alphaCSR[ 53 ][ 93 ],
   alphaCSR[ 53 ][ 94 ],
   alphaCSR[ 53 ][ 95 ],
   alphaCSR[ 53 ][ 96 ],
   alphaCSR[ 53 ][ 97 ],
   alphaCSR[ 53 ][ 98 ],
   alphaCSR[ 53 ][ 99 ],
   alphaCSR[ 53 ][ 100 ],
   alphaCSR[ 53 ][ 101 ],
   alphaCSR[ 53 ][ 102 ],
   alphaCSR[ 53 ][ 103 ],
   alphaCSR[ 53 ][ 104 ],
   alphaCSR[ 53 ][ 105 ],
   alphaCSR[ 53 ][ 106 ],
   alphaCSR[ 53 ][ 107 ],
   alphaCSR[ 53 ][ 108 ],
   alphaCSR[ 53 ][ 109 ],
   alphaCSR[ 53 ][ 110 ],
   alphaCSR[ 53 ][ 111 ],
   alphaCSR[ 53 ][ 112 ],
   alphaCSR[ 53 ][ 113 ],
   alphaCSR[ 53 ][ 114 ],
   alphaCSR[ 53 ][ 115 ],
   alphaCSR[ 53 ][ 116 ],
   alphaCSR[ 53 ][ 117 ],
   alphaCSR[ 53 ][ 118 ],
   alphaCSR[ 53 ][ 119 ],
   alphaCSR[ 53 ][ 120 ],
   alphaCSR[ 53 ][ 121 ],
   alphaCSR[ 53 ][ 122 ],
   alphaCSR[ 53 ][ 123 ],
   alphaCSR[ 53 ][ 124 ],
   alphaCSR[ 53 ][ 125 ],
   alphaCSR[ 53 ][ 126 ],
   alphaCSR[ 53 ][ 127 ],
   alphaCSR[ 53 ][ 128 ],
   alphaCSR[ 53 ][ 129 ],
   alphaCSR[ 53 ][ 130 ],
   alphaCSR[ 53 ][ 131 ],
   alphaCSR[ 53 ][ 132 ],
   alphaCSR[ 53 ][ 133 ],
   alphaCSR[ 53 ][ 134 ],
   alphaCSR[ 53 ][ 135 ],
   alphaCSR[ 53 ][ 136 ],
   alphaCSR[ 53 ][ 137 ],
   alphaCSR[ 53 ][ 138 ],
   alphaCSR[ 53 ][ 139 ],
   alphaCSR[ 53 ][ 140 ],
   alphaCSR[ 53 ][ 141 ],
   alphaCSR[ 53 ][ 142 ],
   alphaCSR[ 53 ][ 143 ],
   alphaCSR[ 53 ][ 144 ],
   alphaCSR[ 53 ][ 145 ],
   alphaCSR[ 53 ][ 146 ],
   alphaCSR[ 53 ][ 147 ],
   alphaCSR[ 53 ][ 148 ],
   alphaCSR[ 53 ][ 149 ],
   alphaCSR[ 53 ][ 150 ],
   alphaCSR[ 53 ][ 151 ],
   alphaCSR[ 53 ][ 152 ],
   alphaCSR[ 53 ][ 153 ],
   alphaCSR[ 53 ][ 154 ],
   alphaCSR[ 53 ][ 155 ],
   alphaCSR[ 53 ][ 156 ],
   alphaCSR[ 53 ][ 157 ],
   alphaCSR[ 53 ][ 158 ],
   alphaCSR[ 53 ][ 159 ],
   alphaCSR[ 53 ][ 160 ],
   alphaCSR[ 53 ][ 161 ],
   alphaCSR[ 53 ][ 162 ],
   alphaCSR[ 53 ][ 163 ],
   alphaCSR[ 53 ][ 164 ],
   alphaCSR[ 53 ][ 165 ],
   alphaCSR[ 53 ][ 166 ],
   alphaCSR[ 53 ][ 167 ],
   alphaCSR[ 53 ][ 168 ],
   alphaCSR[ 53 ][ 169 ],
   alphaCSR[ 53 ][ 170 ],
   alphaCSR[ 53 ][ 171 ],
   alphaCSR[ 53 ][ 172 ],
   alphaCSR[ 53 ][ 173 ],
   alphaCSR[ 53 ][ 174 ],
   alphaCSR[ 53 ][ 175 ],
   alphaCSR[ 53 ][ 176 ],
   alphaCSR[ 53 ][ 177 ],
   alphaCSR[ 53 ][ 178 ],
   alphaCSR[ 53 ][ 179 ],
   alphaCSR[ 53 ][ 180 ],
   alphaCSR[ 53 ][ 181 ],
   alphaCSR[ 53 ][ 182 ],
   alphaCSR[ 53 ][ 183 ],
   alphaCSR[ 53 ][ 184 ],
   alphaCSR[ 53 ][ 185 ],
   alphaCSR[ 53 ][ 186 ],
   alphaCSR[ 53 ][ 187 ],
   alphaCSR[ 53 ][ 188 ],
   alphaCSR[ 53 ][ 189 ],
   alphaCSR[ 53 ][ 190 ],
   alphaCSR[ 53 ][ 191 ],
   alphaCSR[ 53 ][ 192 ],
   alphaCSR[ 53 ][ 193 ],
   alphaCSR[ 53 ][ 194 ],
   alphaCSR[ 53 ][ 195 ],
   alphaCSR[ 53 ][ 196 ],
   alphaCSR[ 53 ][ 197 ],
   alphaCSR[ 53 ][ 198 ],
   alphaCSR[ 53 ][ 199 ],
   alphaCSR[ 53 ][ 200 ],
   alphaCSR[ 53 ][ 201 ],
   alphaCSR[ 53 ][ 202 ],
   alphaCSR[ 53 ][ 203 ],
   alphaCSR[ 53 ][ 204 ],
   alphaCSR[ 53 ][ 205 ],
   alphaCSR[ 53 ][ 206 ],
   alphaCSR[ 53 ][ 207 ],
   alphaCSR[ 53 ][ 208 ],
   alphaCSR[ 53 ][ 209 ],
   alphaCSR[ 53 ][ 210 ],
   alphaCSR[ 53 ][ 211 ],
   alphaCSR[ 53 ][ 212 ],
   alphaCSR[ 53 ][ 213 ],
   alphaCSR[ 53 ][ 214 ],
   alphaCSR[ 53 ][ 215 ],
   alphaCSR[ 53 ][ 216 ],
   alphaCSR[ 53 ][ 217 ],
   alphaCSR[ 53 ][ 218 ],
   alphaCSR[ 53 ][ 219 ],
   alphaCSR[ 53 ][ 220 ],
   alphaCSR[ 53 ][ 221 ],
   alphaCSR[ 53 ][ 222 ],
   alphaCSR[ 53 ][ 223 ],
   alphaCSR[ 53 ][ 224 ],
   alphaCSR[ 53 ][ 225 ],
   alphaCSR[ 53 ][ 226 ],
   alphaCSR[ 53 ][ 227 ],
   alphaCSR[ 53 ][ 228 ],
   alphaCSR[ 53 ][ 229 ],
   alphaCSR[ 53 ][ 230 ],
   alphaCSR[ 53 ][ 231 ],
   alphaCSR[ 53 ][ 232 ],
   alphaCSR[ 53 ][ 233 ],
   alphaCSR[ 53 ][ 234 ],
   alphaCSR[ 53 ][ 235 ],
   alphaCSR[ 53 ][ 236 ],
   alphaCSR[ 53 ][ 237 ],
   alphaCSR[ 53 ][ 238 ],
   alphaCSR[ 53 ][ 239 ],
   alphaCSR[ 53 ][ 240 ],
   alphaCSR[ 53 ][ 241 ],
   alphaCSR[ 53 ][ 242 ],
   alphaCSR[ 53 ][ 243 ],
   alphaCSR[ 53 ][ 244 ],
   alphaCSR[ 53 ][ 245 ],
   alphaCSR[ 53 ][ 246 ],
   alphaCSR[ 53 ][ 247 ],
   alphaCSR[ 53 ][ 248 ],
   alphaCSR[ 53 ][ 249 ],
   alphaCSR[ 53 ][ 250 ],
   alphaCSR[ 53 ][ 251 ],
   alphaCSR[ 53 ][ 252 ],
   alphaCSR[ 53 ][ 253 ],
   alphaCSR[ 53 ][ 254 ],
   alphaCSR[ 53 ][ 255 ],
   alphaCSR[ 53 ][ 256 ],
   alphaCSR[ 53 ][ 257 ],
   alphaCSR[ 53 ][ 258 ],
   alphaCSR[ 53 ][ 259 ],
   alphaCSR[ 53 ][ 260 ],
   alphaCSR[ 53 ][ 261 ],
   alphaCSR[ 53 ][ 262 ],
   alphaCSR[ 53 ][ 263 ],
   alphaCSR[ 53 ][ 264 ],
   alphaCSR[ 53 ][ 265 ],
   alphaCSR[ 53 ][ 266 ],
   alphaCSR[ 53 ][ 267 ],
   alphaCSR[ 53 ][ 268 ],
   alphaCSR[ 53 ][ 269 ],
   alphaCSR[ 53 ][ 270 ],
   alphaCSR[ 53 ][ 271 ],
   alphaCSR[ 53 ][ 272 ],
   alphaCSR[ 53 ][ 273 ],
   alphaCSR[ 53 ][ 274 ],
   alphaCSR[ 53 ][ 275 ],
   alphaCSR[ 53 ][ 276 ],
   alphaCSR[ 53 ][ 277 ],
   alphaCSR[ 53 ][ 278 ],
   alphaCSR[ 53 ][ 279 ],
   alphaCSR[ 53 ][ 280 ],
   alphaCSR[ 53 ][ 281 ],
   alphaCSR[ 53 ][ 282 ],
   alphaCSR[ 53 ][ 283 ],
   alphaCSR[ 53 ][ 284 ],
   alphaCSR[ 53 ][ 285 ],
   alphaCSR[ 53 ][ 286 ],
   alphaCSR[ 53 ][ 287 ],
   alphaCSR[ 53 ][ 288 ],
   alphaCSR[ 53 ][ 289 ],
   alphaCSR[ 53 ][ 290 ],
   alphaCSR[ 53 ][ 291 ],
   alphaCSR[ 53 ][ 292 ],
   alphaCSR[ 53 ][ 293 ],
   alphaCSR[ 53 ][ 294 ],
   alphaCSR[ 53 ][ 295 ],
   alphaCSR[ 53 ][ 296 ],
   alphaCSR[ 53 ][ 297 ],
   alphaCSR[ 53 ][ 298 ],
   alphaCSR[ 53 ][ 299 ],
   alphaCSR[ 53 ][ 300 ],
   alphaCSR[ 53 ][ 301 ],
   alphaCSR[ 53 ][ 302 ],
   alphaCSR[ 53 ][ 303 ],
   alphaCSR[ 53 ][ 304 ],
   alphaCSR[ 53 ][ 305 ],
   alphaCSR[ 53 ][ 306 ],
   alphaCSR[ 53 ][ 307 ],
   alphaCSR[ 53 ][ 308 ],
   alphaCSR[ 53 ][ 309 ],
   alphaCSR[ 53 ][ 310 ],
   alphaCSR[ 53 ][ 311 ],
   alphaCSR[ 53 ][ 312 ],
   alphaCSR[ 53 ][ 313 ],
   alphaCSR[ 53 ][ 314 ],
   alphaCSR[ 53 ][ 315 ],
   alphaCSR[ 53 ][ 316 ],
   alphaCSR[ 53 ][ 317 ],
   alphaCSR[ 53 ][ 318 ],
   alphaCSR[ 53 ][ 319 ],
   alphaCSR[ 53 ][ 320 ],
   alphaCSR[ 53 ][ 321 ],
   alphaCSR[ 53 ][ 322 ],
   alphaCSR[ 53 ][ 323 ],
   alphaCSR[ 53 ][ 324 ],
   alphaCSR[ 53 ][ 325 ],
   alphaCSR[ 53 ][ 326 ],
   alphaCSR[ 53 ][ 327 ],
   alphaCSR[ 53 ][ 328 ],
   alphaCSR[ 53 ][ 329 ],
   alphaCSR[ 53 ][ 330 ],
   alphaCSR[ 53 ][ 331 ],
   alphaCSR[ 53 ][ 332 ],
   alphaCSR[ 53 ][ 333 ],
   alphaCSR[ 53 ][ 334 ],
   alphaCSR[ 53 ][ 335 ],
   alphaCSR[ 53 ][ 336 ],
   alphaCSR[ 53 ][ 337 ],
   alphaCSR[ 53 ][ 338 ],
   alphaCSR[ 53 ][ 339 ],
   alphaCSR[ 53 ][ 340 ],
   alphaCSR[ 53 ][ 341 ],
   alphaCSR[ 53 ][ 342 ],
   alphaCSR[ 53 ][ 343 ],
   alphaCSR[ 53 ][ 344 ],
   alphaCSR[ 53 ][ 345 ],
   alphaCSR[ 53 ][ 346 ],
   alphaCSR[ 53 ][ 347 ],
   alphaCSR[ 53 ][ 348 ],
   alphaCSR[ 53 ][ 349 ],
   alphaCSR[ 53 ][ 350 ],
   alphaCSR[ 53 ][ 351 ],
   alphaCSR[ 53 ][ 352 ],
   alphaCSR[ 53 ][ 353 ],
   alphaCSR[ 53 ][ 354 ],
   alphaCSR[ 53 ][ 355 ],
   alphaCSR[ 53 ][ 356 ],
   alphaCSR[ 53 ][ 357 ],
   alphaCSR[ 53 ][ 358 ],
   alphaCSR[ 53 ][ 359 ],
   alphaCSR[ 53 ][ 360 ],
   alphaCSR[ 53 ][ 361 ],
   alphaCSR[ 53 ][ 362 ],
   alphaCSR[ 53 ][ 363 ],
   alphaCSR[ 53 ][ 364 ],
   alphaCSR[ 53 ][ 365 ],
   alphaCSR[ 53 ][ 366 ],
   alphaCSR[ 53 ][ 367 ],
   alphaCSR[ 53 ][ 368 ],
   alphaCSR[ 53 ][ 369 ],
   alphaCSR[ 53 ][ 370 ],
   alphaCSR[ 53 ][ 371 ],
   alphaCSR[ 53 ][ 372 ],
   alphaCSR[ 53 ][ 373 ],
   alphaCSR[ 53 ][ 374 ],
   alphaCSR[ 53 ][ 375 ],
   alphaCSR[ 53 ][ 376 ],
   alphaCSR[ 53 ][ 377 ],
   alphaCSR[ 53 ][ 378 ],
   alphaCSR[ 53 ][ 379 ],
   alphaCSR[ 53 ][ 380 ],
   alphaCSR[ 53 ][ 381 ],
   alphaCSR[ 53 ][ 382 ],
   alphaCSR[ 53 ][ 383 ],
   alphaCSR[ 54 ][ 0 ],
   alphaCSR[ 54 ][ 1 ],
   alphaCSR[ 54 ][ 2 ],
   alphaCSR[ 54 ][ 3 ],
   alphaCSR[ 54 ][ 4 ],
   alphaCSR[ 54 ][ 5 ],
   alphaCSR[ 54 ][ 6 ],
   alphaCSR[ 54 ][ 7 ],
   alphaCSR[ 54 ][ 8 ],
   alphaCSR[ 54 ][ 9 ],
   alphaCSR[ 54 ][ 10 ],
   alphaCSR[ 54 ][ 11 ],
   alphaCSR[ 54 ][ 12 ],
   alphaCSR[ 54 ][ 13 ],
   alphaCSR[ 54 ][ 14 ],
   alphaCSR[ 54 ][ 15 ],
   alphaCSR[ 54 ][ 16 ],
   alphaCSR[ 54 ][ 17 ],
   alphaCSR[ 54 ][ 18 ],
   alphaCSR[ 54 ][ 19 ],
   alphaCSR[ 54 ][ 20 ],
   alphaCSR[ 54 ][ 21 ],
   alphaCSR[ 54 ][ 22 ],
   alphaCSR[ 54 ][ 23 ],
   alphaCSR[ 54 ][ 24 ],
   alphaCSR[ 54 ][ 25 ],
   alphaCSR[ 54 ][ 26 ],
   alphaCSR[ 54 ][ 27 ],
   alphaCSR[ 54 ][ 28 ],
   alphaCSR[ 54 ][ 29 ],
   alphaCSR[ 54 ][ 30 ],
   alphaCSR[ 54 ][ 31 ],
   alphaCSR[ 54 ][ 32 ],
   alphaCSR[ 54 ][ 33 ],
   alphaCSR[ 54 ][ 34 ],
   alphaCSR[ 54 ][ 35 ],
   alphaCSR[ 54 ][ 36 ],
   alphaCSR[ 54 ][ 37 ],
   alphaCSR[ 54 ][ 38 ],
   alphaCSR[ 54 ][ 39 ],
   alphaCSR[ 54 ][ 40 ],
   alphaCSR[ 54 ][ 41 ],
   alphaCSR[ 54 ][ 42 ],
   alphaCSR[ 54 ][ 43 ],
   alphaCSR[ 54 ][ 44 ],
   alphaCSR[ 54 ][ 45 ],
   alphaCSR[ 54 ][ 46 ],
   alphaCSR[ 54 ][ 47 ],
   alphaCSR[ 54 ][ 48 ],
   alphaCSR[ 54 ][ 49 ],
   alphaCSR[ 54 ][ 50 ],
   alphaCSR[ 54 ][ 51 ],
   alphaCSR[ 54 ][ 52 ],
   alphaCSR[ 54 ][ 53 ],
   alphaCSR[ 54 ][ 54 ],
   alphaCSR[ 54 ][ 55 ],
   alphaCSR[ 54 ][ 56 ],
   alphaCSR[ 54 ][ 57 ],
   alphaCSR[ 54 ][ 58 ],
   alphaCSR[ 54 ][ 59 ],
   alphaCSR[ 54 ][ 60 ],
   alphaCSR[ 54 ][ 61 ],
   alphaCSR[ 54 ][ 62 ],
   alphaCSR[ 54 ][ 63 ],
   alphaCSR[ 54 ][ 64 ],
   alphaCSR[ 54 ][ 65 ],
   alphaCSR[ 54 ][ 66 ],
   alphaCSR[ 54 ][ 67 ],
   alphaCSR[ 54 ][ 68 ],
   alphaCSR[ 54 ][ 69 ],
   alphaCSR[ 54 ][ 70 ],
   alphaCSR[ 54 ][ 71 ],
   alphaCSR[ 54 ][ 72 ],
   alphaCSR[ 54 ][ 73 ],
   alphaCSR[ 54 ][ 74 ],
   alphaCSR[ 54 ][ 75 ],
   alphaCSR[ 54 ][ 76 ],
   alphaCSR[ 54 ][ 77 ],
   alphaCSR[ 54 ][ 78 ],
   alphaCSR[ 54 ][ 79 ],
   alphaCSR[ 54 ][ 80 ],
   alphaCSR[ 54 ][ 81 ],
   alphaCSR[ 54 ][ 82 ],
   alphaCSR[ 54 ][ 83 ],
   alphaCSR[ 54 ][ 84 ],
   alphaCSR[ 54 ][ 85 ],
   alphaCSR[ 54 ][ 86 ],
   alphaCSR[ 54 ][ 87 ],
   alphaCSR[ 54 ][ 88 ],
   alphaCSR[ 54 ][ 89 ],
   alphaCSR[ 54 ][ 90 ],
   alphaCSR[ 54 ][ 91 ],
   alphaCSR[ 54 ][ 92 ],
   alphaCSR[ 54 ][ 93 ],
   alphaCSR[ 54 ][ 94 ],
   alphaCSR[ 54 ][ 95 ],
   alphaCSR[ 54 ][ 96 ],
   alphaCSR[ 54 ][ 97 ],
   alphaCSR[ 54 ][ 98 ],
   alphaCSR[ 54 ][ 99 ],
   alphaCSR[ 54 ][ 100 ],
   alphaCSR[ 54 ][ 101 ],
   alphaCSR[ 54 ][ 102 ],
   alphaCSR[ 54 ][ 103 ],
   alphaCSR[ 54 ][ 104 ],
   alphaCSR[ 54 ][ 105 ],
   alphaCSR[ 54 ][ 106 ],
   alphaCSR[ 54 ][ 107 ],
   alphaCSR[ 54 ][ 108 ],
   alphaCSR[ 54 ][ 109 ],
   alphaCSR[ 54 ][ 110 ],
   alphaCSR[ 54 ][ 111 ],
   alphaCSR[ 54 ][ 112 ],
   alphaCSR[ 54 ][ 113 ],
   alphaCSR[ 54 ][ 114 ],
   alphaCSR[ 54 ][ 115 ],
   alphaCSR[ 54 ][ 116 ],
   alphaCSR[ 54 ][ 117 ],
   alphaCSR[ 54 ][ 118 ],
   alphaCSR[ 54 ][ 119 ],
   alphaCSR[ 54 ][ 120 ],
   alphaCSR[ 54 ][ 121 ],
   alphaCSR[ 54 ][ 122 ],
   alphaCSR[ 54 ][ 123 ],
   alphaCSR[ 54 ][ 124 ],
   alphaCSR[ 54 ][ 125 ],
   alphaCSR[ 54 ][ 126 ],
   alphaCSR[ 54 ][ 127 ],
   alphaCSR[ 54 ][ 128 ],
   alphaCSR[ 54 ][ 129 ],
   alphaCSR[ 54 ][ 130 ],
   alphaCSR[ 54 ][ 131 ],
   alphaCSR[ 54 ][ 132 ],
   alphaCSR[ 54 ][ 133 ],
   alphaCSR[ 54 ][ 134 ],
   alphaCSR[ 54 ][ 135 ],
   alphaCSR[ 54 ][ 136 ],
   alphaCSR[ 54 ][ 137 ],
   alphaCSR[ 54 ][ 138 ],
   alphaCSR[ 54 ][ 139 ],
   alphaCSR[ 54 ][ 140 ],
   alphaCSR[ 54 ][ 141 ],
   alphaCSR[ 54 ][ 142 ],
   alphaCSR[ 54 ][ 143 ],
   alphaCSR[ 54 ][ 144 ],
   alphaCSR[ 54 ][ 145 ],
   alphaCSR[ 54 ][ 146 ],
   alphaCSR[ 54 ][ 147 ],
   alphaCSR[ 54 ][ 148 ],
   alphaCSR[ 54 ][ 149 ],
   alphaCSR[ 54 ][ 150 ],
   alphaCSR[ 54 ][ 151 ],
   alphaCSR[ 54 ][ 152 ],
   alphaCSR[ 54 ][ 153 ],
   alphaCSR[ 54 ][ 154 ],
   alphaCSR[ 54 ][ 155 ],
   alphaCSR[ 54 ][ 156 ],
   alphaCSR[ 54 ][ 157 ],
   alphaCSR[ 54 ][ 158 ],
   alphaCSR[ 54 ][ 159 ],
   alphaCSR[ 54 ][ 160 ],
   alphaCSR[ 54 ][ 161 ],
   alphaCSR[ 54 ][ 162 ],
   alphaCSR[ 54 ][ 163 ],
   alphaCSR[ 54 ][ 164 ],
   alphaCSR[ 54 ][ 165 ],
   alphaCSR[ 54 ][ 166 ],
   alphaCSR[ 54 ][ 167 ],
   alphaCSR[ 54 ][ 168 ],
   alphaCSR[ 54 ][ 169 ],
   alphaCSR[ 54 ][ 170 ],
   alphaCSR[ 54 ][ 171 ],
   alphaCSR[ 54 ][ 172 ],
   alphaCSR[ 54 ][ 173 ],
   alphaCSR[ 54 ][ 174 ],
   alphaCSR[ 54 ][ 175 ],
   alphaCSR[ 54 ][ 176 ],
   alphaCSR[ 54 ][ 177 ],
   alphaCSR[ 54 ][ 178 ],
   alphaCSR[ 54 ][ 179 ],
   alphaCSR[ 54 ][ 180 ],
   alphaCSR[ 54 ][ 181 ],
   alphaCSR[ 54 ][ 182 ],
   alphaCSR[ 54 ][ 183 ],
   alphaCSR[ 54 ][ 184 ],
   alphaCSR[ 54 ][ 185 ],
   alphaCSR[ 54 ][ 186 ],
   alphaCSR[ 54 ][ 187 ],
   alphaCSR[ 54 ][ 188 ],
   alphaCSR[ 54 ][ 189 ],
   alphaCSR[ 54 ][ 190 ],
   alphaCSR[ 54 ][ 191 ],
   alphaCSR[ 54 ][ 192 ],
   alphaCSR[ 54 ][ 193 ],
   alphaCSR[ 54 ][ 194 ],
   alphaCSR[ 54 ][ 195 ],
   alphaCSR[ 54 ][ 196 ],
   alphaCSR[ 54 ][ 197 ],
   alphaCSR[ 54 ][ 198 ],
   alphaCSR[ 54 ][ 199 ],
   alphaCSR[ 54 ][ 200 ],
   alphaCSR[ 54 ][ 201 ],
   alphaCSR[ 54 ][ 202 ],
   alphaCSR[ 54 ][ 203 ],
   alphaCSR[ 54 ][ 204 ],
   alphaCSR[ 54 ][ 205 ],
   alphaCSR[ 54 ][ 206 ],
   alphaCSR[ 54 ][ 207 ],
   alphaCSR[ 54 ][ 208 ],
   alphaCSR[ 54 ][ 209 ],
   alphaCSR[ 54 ][ 210 ],
   alphaCSR[ 54 ][ 211 ],
   alphaCSR[ 54 ][ 212 ],
   alphaCSR[ 54 ][ 213 ],
   alphaCSR[ 54 ][ 214 ],
   alphaCSR[ 54 ][ 215 ],
   alphaCSR[ 54 ][ 216 ],
   alphaCSR[ 54 ][ 217 ],
   alphaCSR[ 54 ][ 218 ],
   alphaCSR[ 54 ][ 219 ],
   alphaCSR[ 54 ][ 220 ],
   alphaCSR[ 54 ][ 221 ],
   alphaCSR[ 54 ][ 222 ],
   alphaCSR[ 54 ][ 223 ],
   alphaCSR[ 54 ][ 224 ],
   alphaCSR[ 54 ][ 225 ],
   alphaCSR[ 54 ][ 226 ],
   alphaCSR[ 54 ][ 227 ],
   alphaCSR[ 54 ][ 228 ],
   alphaCSR[ 54 ][ 229 ],
   alphaCSR[ 54 ][ 230 ],
   alphaCSR[ 54 ][ 231 ],
   alphaCSR[ 54 ][ 232 ],
   alphaCSR[ 54 ][ 233 ],
   alphaCSR[ 54 ][ 234 ],
   alphaCSR[ 54 ][ 235 ],
   alphaCSR[ 54 ][ 236 ],
   alphaCSR[ 54 ][ 237 ],
   alphaCSR[ 54 ][ 238 ],
   alphaCSR[ 54 ][ 239 ],
   alphaCSR[ 54 ][ 240 ],
   alphaCSR[ 54 ][ 241 ],
   alphaCSR[ 54 ][ 242 ],
   alphaCSR[ 54 ][ 243 ],
   alphaCSR[ 54 ][ 244 ],
   alphaCSR[ 54 ][ 245 ],
   alphaCSR[ 54 ][ 246 ],
   alphaCSR[ 54 ][ 247 ],
   alphaCSR[ 54 ][ 248 ],
   alphaCSR[ 54 ][ 249 ],
   alphaCSR[ 54 ][ 250 ],
   alphaCSR[ 54 ][ 251 ],
   alphaCSR[ 54 ][ 252 ],
   alphaCSR[ 54 ][ 253 ],
   alphaCSR[ 54 ][ 254 ],
   alphaCSR[ 54 ][ 255 ],
   alphaCSR[ 54 ][ 256 ],
   alphaCSR[ 54 ][ 257 ],
   alphaCSR[ 54 ][ 258 ],
   alphaCSR[ 54 ][ 259 ],
   alphaCSR[ 54 ][ 260 ],
   alphaCSR[ 54 ][ 261 ],
   alphaCSR[ 54 ][ 262 ],
   alphaCSR[ 54 ][ 263 ],
   alphaCSR[ 54 ][ 264 ],
   alphaCSR[ 54 ][ 265 ],
   alphaCSR[ 54 ][ 266 ],
   alphaCSR[ 54 ][ 267 ],
   alphaCSR[ 54 ][ 268 ],
   alphaCSR[ 54 ][ 269 ],
   alphaCSR[ 54 ][ 270 ],
   alphaCSR[ 54 ][ 271 ],
   alphaCSR[ 54 ][ 272 ],
   alphaCSR[ 54 ][ 273 ],
   alphaCSR[ 54 ][ 274 ],
   alphaCSR[ 54 ][ 275 ],
   alphaCSR[ 54 ][ 276 ],
   alphaCSR[ 54 ][ 277 ],
   alphaCSR[ 54 ][ 278 ],
   alphaCSR[ 54 ][ 279 ],
   alphaCSR[ 54 ][ 280 ],
   alphaCSR[ 54 ][ 281 ],
   alphaCSR[ 54 ][ 282 ],
   alphaCSR[ 54 ][ 283 ],
   alphaCSR[ 54 ][ 284 ],
   alphaCSR[ 54 ][ 285 ],
   alphaCSR[ 54 ][ 286 ],
   alphaCSR[ 54 ][ 287 ],
   alphaCSR[ 54 ][ 288 ],
   alphaCSR[ 54 ][ 289 ],
   alphaCSR[ 54 ][ 290 ],
   alphaCSR[ 54 ][ 291 ],
   alphaCSR[ 54 ][ 292 ],
   alphaCSR[ 54 ][ 293 ],
   alphaCSR[ 54 ][ 294 ],
   alphaCSR[ 54 ][ 295 ],
   alphaCSR[ 54 ][ 296 ],
   alphaCSR[ 54 ][ 297 ],
   alphaCSR[ 54 ][ 298 ],
   alphaCSR[ 54 ][ 299 ],
   alphaCSR[ 54 ][ 300 ],
   alphaCSR[ 54 ][ 301 ],
   alphaCSR[ 54 ][ 302 ],
   alphaCSR[ 54 ][ 303 ],
   alphaCSR[ 54 ][ 304 ],
   alphaCSR[ 54 ][ 305 ],
   alphaCSR[ 54 ][ 306 ],
   alphaCSR[ 54 ][ 307 ],
   alphaCSR[ 54 ][ 308 ],
   alphaCSR[ 54 ][ 309 ],
   alphaCSR[ 54 ][ 310 ],
   alphaCSR[ 54 ][ 311 ],
   alphaCSR[ 54 ][ 312 ],
   alphaCSR[ 54 ][ 313 ],
   alphaCSR[ 54 ][ 314 ],
   alphaCSR[ 54 ][ 315 ],
   alphaCSR[ 54 ][ 316 ],
   alphaCSR[ 54 ][ 317 ],
   alphaCSR[ 54 ][ 318 ],
   alphaCSR[ 54 ][ 319 ],
   alphaCSR[ 54 ][ 320 ],
   alphaCSR[ 54 ][ 321 ],
   alphaCSR[ 54 ][ 322 ],
   alphaCSR[ 54 ][ 323 ],
   alphaCSR[ 54 ][ 324 ],
   alphaCSR[ 54 ][ 325 ],
   alphaCSR[ 54 ][ 326 ],
   alphaCSR[ 54 ][ 327 ],
   alphaCSR[ 54 ][ 328 ],
   alphaCSR[ 54 ][ 329 ],
   alphaCSR[ 54 ][ 330 ],
   alphaCSR[ 54 ][ 331 ],
   alphaCSR[ 54 ][ 332 ],
   alphaCSR[ 54 ][ 333 ],
   alphaCSR[ 54 ][ 334 ],
   alphaCSR[ 54 ][ 335 ],
   alphaCSR[ 54 ][ 336 ],
   alphaCSR[ 54 ][ 337 ],
   alphaCSR[ 54 ][ 338 ],
   alphaCSR[ 54 ][ 339 ],
   alphaCSR[ 54 ][ 340 ],
   alphaCSR[ 54 ][ 341 ],
   alphaCSR[ 54 ][ 342 ],
   alphaCSR[ 54 ][ 343 ],
   alphaCSR[ 54 ][ 344 ],
   alphaCSR[ 54 ][ 345 ],
   alphaCSR[ 54 ][ 346 ],
   alphaCSR[ 54 ][ 347 ],
   alphaCSR[ 54 ][ 348 ],
   alphaCSR[ 54 ][ 349 ],
   alphaCSR[ 54 ][ 350 ],
   alphaCSR[ 54 ][ 351 ],
   alphaCSR[ 54 ][ 352 ],
   alphaCSR[ 54 ][ 353 ],
   alphaCSR[ 54 ][ 354 ],
   alphaCSR[ 54 ][ 355 ],
   alphaCSR[ 54 ][ 356 ],
   alphaCSR[ 54 ][ 357 ],
   alphaCSR[ 54 ][ 358 ],
   alphaCSR[ 54 ][ 359 ],
   alphaCSR[ 54 ][ 360 ],
   alphaCSR[ 54 ][ 361 ],
   alphaCSR[ 54 ][ 362 ],
   alphaCSR[ 54 ][ 363 ],
   alphaCSR[ 54 ][ 364 ],
   alphaCSR[ 54 ][ 365 ],
   alphaCSR[ 54 ][ 366 ],
   alphaCSR[ 54 ][ 367 ],
   alphaCSR[ 54 ][ 368 ],
   alphaCSR[ 54 ][ 369 ],
   alphaCSR[ 54 ][ 370 ],
   alphaCSR[ 54 ][ 371 ],
   alphaCSR[ 54 ][ 372 ],
   alphaCSR[ 54 ][ 373 ],
   alphaCSR[ 54 ][ 374 ],
   alphaCSR[ 54 ][ 375 ],
   alphaCSR[ 54 ][ 376 ],
   alphaCSR[ 54 ][ 377 ],
   alphaCSR[ 54 ][ 378 ],
   alphaCSR[ 54 ][ 379 ],
   alphaCSR[ 54 ][ 380 ],
   alphaCSR[ 54 ][ 381 ],
   alphaCSR[ 54 ][ 382 ],
   alphaCSR[ 54 ][ 383 ],
   alphaCSR[ 55 ][ 0 ],
   alphaCSR[ 55 ][ 1 ],
   alphaCSR[ 55 ][ 2 ],
   alphaCSR[ 55 ][ 3 ],
   alphaCSR[ 55 ][ 4 ],
   alphaCSR[ 55 ][ 5 ],
   alphaCSR[ 55 ][ 6 ],
   alphaCSR[ 55 ][ 7 ],
   alphaCSR[ 55 ][ 8 ],
   alphaCSR[ 55 ][ 9 ],
   alphaCSR[ 55 ][ 10 ],
   alphaCSR[ 55 ][ 11 ],
   alphaCSR[ 55 ][ 12 ],
   alphaCSR[ 55 ][ 13 ],
   alphaCSR[ 55 ][ 14 ],
   alphaCSR[ 55 ][ 15 ],
   alphaCSR[ 55 ][ 16 ],
   alphaCSR[ 55 ][ 17 ],
   alphaCSR[ 55 ][ 18 ],
   alphaCSR[ 55 ][ 19 ],
   alphaCSR[ 55 ][ 20 ],
   alphaCSR[ 55 ][ 21 ],
   alphaCSR[ 55 ][ 22 ],
   alphaCSR[ 55 ][ 23 ],
   alphaCSR[ 55 ][ 24 ],
   alphaCSR[ 55 ][ 25 ],
   alphaCSR[ 55 ][ 26 ],
   alphaCSR[ 55 ][ 27 ],
   alphaCSR[ 55 ][ 28 ],
   alphaCSR[ 55 ][ 29 ],
   alphaCSR[ 55 ][ 30 ],
   alphaCSR[ 55 ][ 31 ],
   alphaCSR[ 55 ][ 32 ],
   alphaCSR[ 55 ][ 33 ],
   alphaCSR[ 55 ][ 34 ],
   alphaCSR[ 55 ][ 35 ],
   alphaCSR[ 55 ][ 36 ],
   alphaCSR[ 55 ][ 37 ],
   alphaCSR[ 55 ][ 38 ],
   alphaCSR[ 55 ][ 39 ],
   alphaCSR[ 55 ][ 40 ],
   alphaCSR[ 55 ][ 41 ],
   alphaCSR[ 55 ][ 42 ],
   alphaCSR[ 55 ][ 43 ],
   alphaCSR[ 55 ][ 44 ],
   alphaCSR[ 55 ][ 45 ],
   alphaCSR[ 55 ][ 46 ],
   alphaCSR[ 55 ][ 47 ],
   alphaCSR[ 55 ][ 48 ],
   alphaCSR[ 55 ][ 49 ],
   alphaCSR[ 55 ][ 50 ],
   alphaCSR[ 55 ][ 51 ],
   alphaCSR[ 55 ][ 52 ],
   alphaCSR[ 55 ][ 53 ],
   alphaCSR[ 55 ][ 54 ],
   alphaCSR[ 55 ][ 55 ],
   alphaCSR[ 55 ][ 56 ],
   alphaCSR[ 55 ][ 57 ],
   alphaCSR[ 55 ][ 58 ],
   alphaCSR[ 55 ][ 59 ],
   alphaCSR[ 55 ][ 60 ],
   alphaCSR[ 55 ][ 61 ],
   alphaCSR[ 55 ][ 62 ],
   alphaCSR[ 55 ][ 63 ],
   alphaCSR[ 55 ][ 64 ],
   alphaCSR[ 55 ][ 65 ],
   alphaCSR[ 55 ][ 66 ],
   alphaCSR[ 55 ][ 67 ],
   alphaCSR[ 55 ][ 68 ],
   alphaCSR[ 55 ][ 69 ],
   alphaCSR[ 55 ][ 70 ],
   alphaCSR[ 55 ][ 71 ],
   alphaCSR[ 55 ][ 72 ],
   alphaCSR[ 55 ][ 73 ],
   alphaCSR[ 55 ][ 74 ],
   alphaCSR[ 55 ][ 75 ],
   alphaCSR[ 55 ][ 76 ],
   alphaCSR[ 55 ][ 77 ],
   alphaCSR[ 55 ][ 78 ],
   alphaCSR[ 55 ][ 79 ],
   alphaCSR[ 55 ][ 80 ],
   alphaCSR[ 55 ][ 81 ],
   alphaCSR[ 55 ][ 82 ],
   alphaCSR[ 55 ][ 83 ],
   alphaCSR[ 55 ][ 84 ],
   alphaCSR[ 55 ][ 85 ],
   alphaCSR[ 55 ][ 86 ],
   alphaCSR[ 55 ][ 87 ],
   alphaCSR[ 55 ][ 88 ],
   alphaCSR[ 55 ][ 89 ],
   alphaCSR[ 55 ][ 90 ],
   alphaCSR[ 55 ][ 91 ],
   alphaCSR[ 55 ][ 92 ],
   alphaCSR[ 55 ][ 93 ],
   alphaCSR[ 55 ][ 94 ],
   alphaCSR[ 55 ][ 95 ],
   alphaCSR[ 55 ][ 96 ],
   alphaCSR[ 55 ][ 97 ],
   alphaCSR[ 55 ][ 98 ],
   alphaCSR[ 55 ][ 99 ],
   alphaCSR[ 55 ][ 100 ],
   alphaCSR[ 55 ][ 101 ],
   alphaCSR[ 55 ][ 102 ],
   alphaCSR[ 55 ][ 103 ],
   alphaCSR[ 55 ][ 104 ],
   alphaCSR[ 55 ][ 105 ],
   alphaCSR[ 55 ][ 106 ],
   alphaCSR[ 55 ][ 107 ],
   alphaCSR[ 55 ][ 108 ],
   alphaCSR[ 55 ][ 109 ],
   alphaCSR[ 55 ][ 110 ],
   alphaCSR[ 55 ][ 111 ],
   alphaCSR[ 55 ][ 112 ],
   alphaCSR[ 55 ][ 113 ],
   alphaCSR[ 55 ][ 114 ],
   alphaCSR[ 55 ][ 115 ],
   alphaCSR[ 55 ][ 116 ],
   alphaCSR[ 55 ][ 117 ],
   alphaCSR[ 55 ][ 118 ],
   alphaCSR[ 55 ][ 119 ],
   alphaCSR[ 55 ][ 120 ],
   alphaCSR[ 55 ][ 121 ],
   alphaCSR[ 55 ][ 122 ],
   alphaCSR[ 55 ][ 123 ],
   alphaCSR[ 55 ][ 124 ],
   alphaCSR[ 55 ][ 125 ],
   alphaCSR[ 55 ][ 126 ],
   alphaCSR[ 55 ][ 127 ],
   alphaCSR[ 55 ][ 128 ],
   alphaCSR[ 55 ][ 129 ],
   alphaCSR[ 55 ][ 130 ],
   alphaCSR[ 55 ][ 131 ],
   alphaCSR[ 55 ][ 132 ],
   alphaCSR[ 55 ][ 133 ],
   alphaCSR[ 55 ][ 134 ],
   alphaCSR[ 55 ][ 135 ],
   alphaCSR[ 55 ][ 136 ],
   alphaCSR[ 55 ][ 137 ],
   alphaCSR[ 55 ][ 138 ],
   alphaCSR[ 55 ][ 139 ],
   alphaCSR[ 55 ][ 140 ],
   alphaCSR[ 55 ][ 141 ],
   alphaCSR[ 55 ][ 142 ],
   alphaCSR[ 55 ][ 143 ],
   alphaCSR[ 55 ][ 144 ],
   alphaCSR[ 55 ][ 145 ],
   alphaCSR[ 55 ][ 146 ],
   alphaCSR[ 55 ][ 147 ],
   alphaCSR[ 55 ][ 148 ],
   alphaCSR[ 55 ][ 149 ],
   alphaCSR[ 55 ][ 150 ],
   alphaCSR[ 55 ][ 151 ],
   alphaCSR[ 55 ][ 152 ],
   alphaCSR[ 55 ][ 153 ],
   alphaCSR[ 55 ][ 154 ],
   alphaCSR[ 55 ][ 155 ],
   alphaCSR[ 55 ][ 156 ],
   alphaCSR[ 55 ][ 157 ],
   alphaCSR[ 55 ][ 158 ],
   alphaCSR[ 55 ][ 159 ],
   alphaCSR[ 55 ][ 160 ],
   alphaCSR[ 55 ][ 161 ],
   alphaCSR[ 55 ][ 162 ],
   alphaCSR[ 55 ][ 163 ],
   alphaCSR[ 55 ][ 164 ],
   alphaCSR[ 55 ][ 165 ],
   alphaCSR[ 55 ][ 166 ],
   alphaCSR[ 55 ][ 167 ],
   alphaCSR[ 55 ][ 168 ],
   alphaCSR[ 55 ][ 169 ],
   alphaCSR[ 55 ][ 170 ],
   alphaCSR[ 55 ][ 171 ],
   alphaCSR[ 55 ][ 172 ],
   alphaCSR[ 55 ][ 173 ],
   alphaCSR[ 55 ][ 174 ],
   alphaCSR[ 55 ][ 175 ],
   alphaCSR[ 55 ][ 176 ],
   alphaCSR[ 55 ][ 177 ],
   alphaCSR[ 55 ][ 178 ],
   alphaCSR[ 55 ][ 179 ],
   alphaCSR[ 55 ][ 180 ],
   alphaCSR[ 55 ][ 181 ],
   alphaCSR[ 55 ][ 182 ],
   alphaCSR[ 55 ][ 183 ],
   alphaCSR[ 55 ][ 184 ],
   alphaCSR[ 55 ][ 185 ],
   alphaCSR[ 55 ][ 186 ],
   alphaCSR[ 55 ][ 187 ],
   alphaCSR[ 55 ][ 188 ],
   alphaCSR[ 55 ][ 189 ],
   alphaCSR[ 55 ][ 190 ],
   alphaCSR[ 55 ][ 191 ],
   alphaCSR[ 55 ][ 192 ],
   alphaCSR[ 55 ][ 193 ],
   alphaCSR[ 55 ][ 194 ],
   alphaCSR[ 55 ][ 195 ],
   alphaCSR[ 55 ][ 196 ],
   alphaCSR[ 55 ][ 197 ],
   alphaCSR[ 55 ][ 198 ],
   alphaCSR[ 55 ][ 199 ],
   alphaCSR[ 55 ][ 200 ],
   alphaCSR[ 55 ][ 201 ],
   alphaCSR[ 55 ][ 202 ],
   alphaCSR[ 55 ][ 203 ],
   alphaCSR[ 55 ][ 204 ],
   alphaCSR[ 55 ][ 205 ],
   alphaCSR[ 55 ][ 206 ],
   alphaCSR[ 55 ][ 207 ],
   alphaCSR[ 55 ][ 208 ],
   alphaCSR[ 55 ][ 209 ],
   alphaCSR[ 55 ][ 210 ],
   alphaCSR[ 55 ][ 211 ],
   alphaCSR[ 55 ][ 212 ],
   alphaCSR[ 55 ][ 213 ],
   alphaCSR[ 55 ][ 214 ],
   alphaCSR[ 55 ][ 215 ],
   alphaCSR[ 55 ][ 216 ],
   alphaCSR[ 55 ][ 217 ],
   alphaCSR[ 55 ][ 218 ],
   alphaCSR[ 55 ][ 219 ],
   alphaCSR[ 55 ][ 220 ],
   alphaCSR[ 55 ][ 221 ],
   alphaCSR[ 55 ][ 222 ],
   alphaCSR[ 55 ][ 223 ],
   alphaCSR[ 55 ][ 224 ],
   alphaCSR[ 55 ][ 225 ],
   alphaCSR[ 55 ][ 226 ],
   alphaCSR[ 55 ][ 227 ],
   alphaCSR[ 55 ][ 228 ],
   alphaCSR[ 55 ][ 229 ],
   alphaCSR[ 55 ][ 230 ],
   alphaCSR[ 55 ][ 231 ],
   alphaCSR[ 55 ][ 232 ],
   alphaCSR[ 55 ][ 233 ],
   alphaCSR[ 55 ][ 234 ],
   alphaCSR[ 55 ][ 235 ],
   alphaCSR[ 55 ][ 236 ],
   alphaCSR[ 55 ][ 237 ],
   alphaCSR[ 55 ][ 238 ],
   alphaCSR[ 55 ][ 239 ],
   alphaCSR[ 55 ][ 240 ],
   alphaCSR[ 55 ][ 241 ],
   alphaCSR[ 55 ][ 242 ],
   alphaCSR[ 55 ][ 243 ],
   alphaCSR[ 55 ][ 244 ],
   alphaCSR[ 55 ][ 245 ],
   alphaCSR[ 55 ][ 246 ],
   alphaCSR[ 55 ][ 247 ],
   alphaCSR[ 55 ][ 248 ],
   alphaCSR[ 55 ][ 249 ],
   alphaCSR[ 55 ][ 250 ],
   alphaCSR[ 55 ][ 251 ],
   alphaCSR[ 55 ][ 252 ],
   alphaCSR[ 55 ][ 253 ],
   alphaCSR[ 55 ][ 254 ],
   alphaCSR[ 55 ][ 255 ],
   alphaCSR[ 55 ][ 256 ],
   alphaCSR[ 55 ][ 257 ],
   alphaCSR[ 55 ][ 258 ],
   alphaCSR[ 55 ][ 259 ],
   alphaCSR[ 55 ][ 260 ],
   alphaCSR[ 55 ][ 261 ],
   alphaCSR[ 55 ][ 262 ],
   alphaCSR[ 55 ][ 263 ],
   alphaCSR[ 55 ][ 264 ],
   alphaCSR[ 55 ][ 265 ],
   alphaCSR[ 55 ][ 266 ],
   alphaCSR[ 55 ][ 267 ],
   alphaCSR[ 55 ][ 268 ],
   alphaCSR[ 55 ][ 269 ],
   alphaCSR[ 55 ][ 270 ],
   alphaCSR[ 55 ][ 271 ],
   alphaCSR[ 55 ][ 272 ],
   alphaCSR[ 55 ][ 273 ],
   alphaCSR[ 55 ][ 274 ],
   alphaCSR[ 55 ][ 275 ],
   alphaCSR[ 55 ][ 276 ],
   alphaCSR[ 55 ][ 277 ],
   alphaCSR[ 55 ][ 278 ],
   alphaCSR[ 55 ][ 279 ],
   alphaCSR[ 55 ][ 280 ],
   alphaCSR[ 55 ][ 281 ],
   alphaCSR[ 55 ][ 282 ],
   alphaCSR[ 55 ][ 283 ],
   alphaCSR[ 55 ][ 284 ],
   alphaCSR[ 55 ][ 285 ],
   alphaCSR[ 55 ][ 286 ],
   alphaCSR[ 55 ][ 287 ],
   alphaCSR[ 55 ][ 288 ],
   alphaCSR[ 55 ][ 289 ],
   alphaCSR[ 55 ][ 290 ],
   alphaCSR[ 55 ][ 291 ],
   alphaCSR[ 55 ][ 292 ],
   alphaCSR[ 55 ][ 293 ],
   alphaCSR[ 55 ][ 294 ],
   alphaCSR[ 55 ][ 295 ],
   alphaCSR[ 55 ][ 296 ],
   alphaCSR[ 55 ][ 297 ],
   alphaCSR[ 55 ][ 298 ],
   alphaCSR[ 55 ][ 299 ],
   alphaCSR[ 55 ][ 300 ],
   alphaCSR[ 55 ][ 301 ],
   alphaCSR[ 55 ][ 302 ],
   alphaCSR[ 55 ][ 303 ],
   alphaCSR[ 55 ][ 304 ],
   alphaCSR[ 55 ][ 305 ],
   alphaCSR[ 55 ][ 306 ],
   alphaCSR[ 55 ][ 307 ],
   alphaCSR[ 55 ][ 308 ],
   alphaCSR[ 55 ][ 309 ],
   alphaCSR[ 55 ][ 310 ],
   alphaCSR[ 55 ][ 311 ],
   alphaCSR[ 55 ][ 312 ],
   alphaCSR[ 55 ][ 313 ],
   alphaCSR[ 55 ][ 314 ],
   alphaCSR[ 55 ][ 315 ],
   alphaCSR[ 55 ][ 316 ],
   alphaCSR[ 55 ][ 317 ],
   alphaCSR[ 55 ][ 318 ],
   alphaCSR[ 55 ][ 319 ],
   alphaCSR[ 55 ][ 320 ],
   alphaCSR[ 55 ][ 321 ],
   alphaCSR[ 55 ][ 322 ],
   alphaCSR[ 55 ][ 323 ],
   alphaCSR[ 55 ][ 324 ],
   alphaCSR[ 55 ][ 325 ],
   alphaCSR[ 55 ][ 326 ],
   alphaCSR[ 55 ][ 327 ],
   alphaCSR[ 55 ][ 328 ],
   alphaCSR[ 55 ][ 329 ],
   alphaCSR[ 55 ][ 330 ],
   alphaCSR[ 55 ][ 331 ],
   alphaCSR[ 55 ][ 332 ],
   alphaCSR[ 55 ][ 333 ],
   alphaCSR[ 55 ][ 334 ],
   alphaCSR[ 55 ][ 335 ],
   alphaCSR[ 55 ][ 336 ],
   alphaCSR[ 55 ][ 337 ],
   alphaCSR[ 55 ][ 338 ],
   alphaCSR[ 55 ][ 339 ],
   alphaCSR[ 55 ][ 340 ],
   alphaCSR[ 55 ][ 341 ],
   alphaCSR[ 55 ][ 342 ],
   alphaCSR[ 55 ][ 343 ],
   alphaCSR[ 55 ][ 344 ],
   alphaCSR[ 55 ][ 345 ],
   alphaCSR[ 55 ][ 346 ],
   alphaCSR[ 55 ][ 347 ],
   alphaCSR[ 55 ][ 348 ],
   alphaCSR[ 55 ][ 349 ],
   alphaCSR[ 55 ][ 350 ],
   alphaCSR[ 55 ][ 351 ],
   alphaCSR[ 55 ][ 352 ],
   alphaCSR[ 55 ][ 353 ],
   alphaCSR[ 55 ][ 354 ],
   alphaCSR[ 55 ][ 355 ],
   alphaCSR[ 55 ][ 356 ],
   alphaCSR[ 55 ][ 357 ],
   alphaCSR[ 55 ][ 358 ],
   alphaCSR[ 55 ][ 359 ],
   alphaCSR[ 55 ][ 360 ],
   alphaCSR[ 55 ][ 361 ],
   alphaCSR[ 55 ][ 362 ],
   alphaCSR[ 55 ][ 363 ],
   alphaCSR[ 55 ][ 364 ],
   alphaCSR[ 55 ][ 365 ],
   alphaCSR[ 55 ][ 366 ],
   alphaCSR[ 55 ][ 367 ],
   alphaCSR[ 55 ][ 368 ],
   alphaCSR[ 55 ][ 369 ],
   alphaCSR[ 55 ][ 370 ],
   alphaCSR[ 55 ][ 371 ],
   alphaCSR[ 55 ][ 372 ],
   alphaCSR[ 55 ][ 373 ],
   alphaCSR[ 55 ][ 374 ],
   alphaCSR[ 55 ][ 375 ],
   alphaCSR[ 55 ][ 376 ],
   alphaCSR[ 55 ][ 377 ],
   alphaCSR[ 55 ][ 378 ],
   alphaCSR[ 55 ][ 379 ],
   alphaCSR[ 55 ][ 380 ],
   alphaCSR[ 55 ][ 381 ],
   alphaCSR[ 55 ][ 382 ],
   alphaCSR[ 55 ][ 383 ],
   alphaCSR[ 56 ][ 0 ],
   alphaCSR[ 56 ][ 1 ],
   alphaCSR[ 56 ][ 2 ],
   alphaCSR[ 56 ][ 3 ],
   alphaCSR[ 56 ][ 4 ],
   alphaCSR[ 56 ][ 5 ],
   alphaCSR[ 56 ][ 6 ],
   alphaCSR[ 56 ][ 7 ],
   alphaCSR[ 56 ][ 8 ],
   alphaCSR[ 56 ][ 9 ],
   alphaCSR[ 56 ][ 10 ],
   alphaCSR[ 56 ][ 11 ],
   alphaCSR[ 56 ][ 12 ],
   alphaCSR[ 56 ][ 13 ],
   alphaCSR[ 56 ][ 14 ],
   alphaCSR[ 56 ][ 15 ],
   alphaCSR[ 56 ][ 16 ],
   alphaCSR[ 56 ][ 17 ],
   alphaCSR[ 56 ][ 18 ],
   alphaCSR[ 56 ][ 19 ],
   alphaCSR[ 56 ][ 20 ],
   alphaCSR[ 56 ][ 21 ],
   alphaCSR[ 56 ][ 22 ],
   alphaCSR[ 56 ][ 23 ],
   alphaCSR[ 56 ][ 24 ],
   alphaCSR[ 56 ][ 25 ],
   alphaCSR[ 56 ][ 26 ],
   alphaCSR[ 56 ][ 27 ],
   alphaCSR[ 56 ][ 28 ],
   alphaCSR[ 56 ][ 29 ],
   alphaCSR[ 56 ][ 30 ],
   alphaCSR[ 56 ][ 31 ],
   alphaCSR[ 56 ][ 32 ],
   alphaCSR[ 56 ][ 33 ],
   alphaCSR[ 56 ][ 34 ],
   alphaCSR[ 56 ][ 35 ],
   alphaCSR[ 56 ][ 36 ],
   alphaCSR[ 56 ][ 37 ],
   alphaCSR[ 56 ][ 38 ],
   alphaCSR[ 56 ][ 39 ],
   alphaCSR[ 56 ][ 40 ],
   alphaCSR[ 56 ][ 41 ],
   alphaCSR[ 56 ][ 42 ],
   alphaCSR[ 56 ][ 43 ],
   alphaCSR[ 56 ][ 44 ],
   alphaCSR[ 56 ][ 45 ],
   alphaCSR[ 56 ][ 46 ],
   alphaCSR[ 56 ][ 47 ],
   alphaCSR[ 56 ][ 48 ],
   alphaCSR[ 56 ][ 49 ],
   alphaCSR[ 56 ][ 50 ],
   alphaCSR[ 56 ][ 51 ],
   alphaCSR[ 56 ][ 52 ],
   alphaCSR[ 56 ][ 53 ],
   alphaCSR[ 56 ][ 54 ],
   alphaCSR[ 56 ][ 55 ],
   alphaCSR[ 56 ][ 56 ],
   alphaCSR[ 56 ][ 57 ],
   alphaCSR[ 56 ][ 58 ],
   alphaCSR[ 56 ][ 59 ],
   alphaCSR[ 56 ][ 60 ],
   alphaCSR[ 56 ][ 61 ],
   alphaCSR[ 56 ][ 62 ],
   alphaCSR[ 56 ][ 63 ],
   alphaCSR[ 56 ][ 64 ],
   alphaCSR[ 56 ][ 65 ],
   alphaCSR[ 56 ][ 66 ],
   alphaCSR[ 56 ][ 67 ],
   alphaCSR[ 56 ][ 68 ],
   alphaCSR[ 56 ][ 69 ],
   alphaCSR[ 56 ][ 70 ],
   alphaCSR[ 56 ][ 71 ],
   alphaCSR[ 56 ][ 72 ],
   alphaCSR[ 56 ][ 73 ],
   alphaCSR[ 56 ][ 74 ],
   alphaCSR[ 56 ][ 75 ],
   alphaCSR[ 56 ][ 76 ],
   alphaCSR[ 56 ][ 77 ],
   alphaCSR[ 56 ][ 78 ],
   alphaCSR[ 56 ][ 79 ],
   alphaCSR[ 56 ][ 80 ],
   alphaCSR[ 56 ][ 81 ],
   alphaCSR[ 56 ][ 82 ],
   alphaCSR[ 56 ][ 83 ],
   alphaCSR[ 56 ][ 84 ],
   alphaCSR[ 56 ][ 85 ],
   alphaCSR[ 56 ][ 86 ],
   alphaCSR[ 56 ][ 87 ],
   alphaCSR[ 56 ][ 88 ],
   alphaCSR[ 56 ][ 89 ],
   alphaCSR[ 56 ][ 90 ],
   alphaCSR[ 56 ][ 91 ],
   alphaCSR[ 56 ][ 92 ],
   alphaCSR[ 56 ][ 93 ],
   alphaCSR[ 56 ][ 94 ],
   alphaCSR[ 56 ][ 95 ],
   alphaCSR[ 56 ][ 96 ],
   alphaCSR[ 56 ][ 97 ],
   alphaCSR[ 56 ][ 98 ],
   alphaCSR[ 56 ][ 99 ],
   alphaCSR[ 56 ][ 100 ],
   alphaCSR[ 56 ][ 101 ],
   alphaCSR[ 56 ][ 102 ],
   alphaCSR[ 56 ][ 103 ],
   alphaCSR[ 56 ][ 104 ],
   alphaCSR[ 56 ][ 105 ],
   alphaCSR[ 56 ][ 106 ],
   alphaCSR[ 56 ][ 107 ],
   alphaCSR[ 56 ][ 108 ],
   alphaCSR[ 56 ][ 109 ],
   alphaCSR[ 56 ][ 110 ],
   alphaCSR[ 56 ][ 111 ],
   alphaCSR[ 56 ][ 112 ],
   alphaCSR[ 56 ][ 113 ],
   alphaCSR[ 56 ][ 114 ],
   alphaCSR[ 56 ][ 115 ],
   alphaCSR[ 56 ][ 116 ],
   alphaCSR[ 56 ][ 117 ],
   alphaCSR[ 56 ][ 118 ],
   alphaCSR[ 56 ][ 119 ],
   alphaCSR[ 56 ][ 120 ],
   alphaCSR[ 56 ][ 121 ],
   alphaCSR[ 56 ][ 122 ],
   alphaCSR[ 56 ][ 123 ],
   alphaCSR[ 56 ][ 124 ],
   alphaCSR[ 56 ][ 125 ],
   alphaCSR[ 56 ][ 126 ],
   alphaCSR[ 56 ][ 127 ],
   alphaCSR[ 56 ][ 128 ],
   alphaCSR[ 56 ][ 129 ],
   alphaCSR[ 56 ][ 130 ],
   alphaCSR[ 56 ][ 131 ],
   alphaCSR[ 56 ][ 132 ],
   alphaCSR[ 56 ][ 133 ],
   alphaCSR[ 56 ][ 134 ],
   alphaCSR[ 56 ][ 135 ],
   alphaCSR[ 56 ][ 136 ],
   alphaCSR[ 56 ][ 137 ],
   alphaCSR[ 56 ][ 138 ],
   alphaCSR[ 56 ][ 139 ],
   alphaCSR[ 56 ][ 140 ],
   alphaCSR[ 56 ][ 141 ],
   alphaCSR[ 56 ][ 142 ],
   alphaCSR[ 56 ][ 143 ],
   alphaCSR[ 56 ][ 144 ],
   alphaCSR[ 56 ][ 145 ],
   alphaCSR[ 56 ][ 146 ],
   alphaCSR[ 56 ][ 147 ],
   alphaCSR[ 56 ][ 148 ],
   alphaCSR[ 56 ][ 149 ],
   alphaCSR[ 56 ][ 150 ],
   alphaCSR[ 56 ][ 151 ],
   alphaCSR[ 56 ][ 152 ],
   alphaCSR[ 56 ][ 153 ],
   alphaCSR[ 56 ][ 154 ],
   alphaCSR[ 56 ][ 155 ],
   alphaCSR[ 56 ][ 156 ],
   alphaCSR[ 56 ][ 157 ],
   alphaCSR[ 56 ][ 158 ],
   alphaCSR[ 56 ][ 159 ],
   alphaCSR[ 56 ][ 160 ],
   alphaCSR[ 56 ][ 161 ],
   alphaCSR[ 56 ][ 162 ],
   alphaCSR[ 56 ][ 163 ],
   alphaCSR[ 56 ][ 164 ],
   alphaCSR[ 56 ][ 165 ],
   alphaCSR[ 56 ][ 166 ],
   alphaCSR[ 56 ][ 167 ],
   alphaCSR[ 56 ][ 168 ],
   alphaCSR[ 56 ][ 169 ],
   alphaCSR[ 56 ][ 170 ],
   alphaCSR[ 56 ][ 171 ],
   alphaCSR[ 56 ][ 172 ],
   alphaCSR[ 56 ][ 173 ],
   alphaCSR[ 56 ][ 174 ],
   alphaCSR[ 56 ][ 175 ],
   alphaCSR[ 56 ][ 176 ],
   alphaCSR[ 56 ][ 177 ],
   alphaCSR[ 56 ][ 178 ],
   alphaCSR[ 56 ][ 179 ],
   alphaCSR[ 56 ][ 180 ],
   alphaCSR[ 56 ][ 181 ],
   alphaCSR[ 56 ][ 182 ],
   alphaCSR[ 56 ][ 183 ],
   alphaCSR[ 56 ][ 184 ],
   alphaCSR[ 56 ][ 185 ],
   alphaCSR[ 56 ][ 186 ],
   alphaCSR[ 56 ][ 187 ],
   alphaCSR[ 56 ][ 188 ],
   alphaCSR[ 56 ][ 189 ],
   alphaCSR[ 56 ][ 190 ],
   alphaCSR[ 56 ][ 191 ],
   alphaCSR[ 56 ][ 192 ],
   alphaCSR[ 56 ][ 193 ],
   alphaCSR[ 56 ][ 194 ],
   alphaCSR[ 56 ][ 195 ],
   alphaCSR[ 56 ][ 196 ],
   alphaCSR[ 56 ][ 197 ],
   alphaCSR[ 56 ][ 198 ],
   alphaCSR[ 56 ][ 199 ],
   alphaCSR[ 56 ][ 200 ],
   alphaCSR[ 56 ][ 201 ],
   alphaCSR[ 56 ][ 202 ],
   alphaCSR[ 56 ][ 203 ],
   alphaCSR[ 56 ][ 204 ],
   alphaCSR[ 56 ][ 205 ],
   alphaCSR[ 56 ][ 206 ],
   alphaCSR[ 56 ][ 207 ],
   alphaCSR[ 56 ][ 208 ],
   alphaCSR[ 56 ][ 209 ],
   alphaCSR[ 56 ][ 210 ],
   alphaCSR[ 56 ][ 211 ],
   alphaCSR[ 56 ][ 212 ],
   alphaCSR[ 56 ][ 213 ],
   alphaCSR[ 56 ][ 214 ],
   alphaCSR[ 56 ][ 215 ],
   alphaCSR[ 56 ][ 216 ],
   alphaCSR[ 56 ][ 217 ],
   alphaCSR[ 56 ][ 218 ],
   alphaCSR[ 56 ][ 219 ],
   alphaCSR[ 56 ][ 220 ],
   alphaCSR[ 56 ][ 221 ],
   alphaCSR[ 56 ][ 222 ],
   alphaCSR[ 56 ][ 223 ],
   alphaCSR[ 56 ][ 224 ],
   alphaCSR[ 56 ][ 225 ],
   alphaCSR[ 56 ][ 226 ],
   alphaCSR[ 56 ][ 227 ],
   alphaCSR[ 56 ][ 228 ],
   alphaCSR[ 56 ][ 229 ],
   alphaCSR[ 56 ][ 230 ],
   alphaCSR[ 56 ][ 231 ],
   alphaCSR[ 56 ][ 232 ],
   alphaCSR[ 56 ][ 233 ],
   alphaCSR[ 56 ][ 234 ],
   alphaCSR[ 56 ][ 235 ],
   alphaCSR[ 56 ][ 236 ],
   alphaCSR[ 56 ][ 237 ],
   alphaCSR[ 56 ][ 238 ],
   alphaCSR[ 56 ][ 239 ],
   alphaCSR[ 56 ][ 240 ],
   alphaCSR[ 56 ][ 241 ],
   alphaCSR[ 56 ][ 242 ],
   alphaCSR[ 56 ][ 243 ],
   alphaCSR[ 56 ][ 244 ],
   alphaCSR[ 56 ][ 245 ],
   alphaCSR[ 56 ][ 246 ],
   alphaCSR[ 56 ][ 247 ],
   alphaCSR[ 56 ][ 248 ],
   alphaCSR[ 56 ][ 249 ],
   alphaCSR[ 56 ][ 250 ],
   alphaCSR[ 56 ][ 251 ],
   alphaCSR[ 56 ][ 252 ],
   alphaCSR[ 56 ][ 253 ],
   alphaCSR[ 56 ][ 254 ],
   alphaCSR[ 56 ][ 255 ],
   alphaCSR[ 56 ][ 256 ],
   alphaCSR[ 56 ][ 257 ],
   alphaCSR[ 56 ][ 258 ],
   alphaCSR[ 56 ][ 259 ],
   alphaCSR[ 56 ][ 260 ],
   alphaCSR[ 56 ][ 261 ],
   alphaCSR[ 56 ][ 262 ],
   alphaCSR[ 56 ][ 263 ],
   alphaCSR[ 56 ][ 264 ],
   alphaCSR[ 56 ][ 265 ],
   alphaCSR[ 56 ][ 266 ],
   alphaCSR[ 56 ][ 267 ],
   alphaCSR[ 56 ][ 268 ],
   alphaCSR[ 56 ][ 269 ],
   alphaCSR[ 56 ][ 270 ],
   alphaCSR[ 56 ][ 271 ],
   alphaCSR[ 56 ][ 272 ],
   alphaCSR[ 56 ][ 273 ],
   alphaCSR[ 56 ][ 274 ],
   alphaCSR[ 56 ][ 275 ],
   alphaCSR[ 56 ][ 276 ],
   alphaCSR[ 56 ][ 277 ],
   alphaCSR[ 56 ][ 278 ],
   alphaCSR[ 56 ][ 279 ],
   alphaCSR[ 56 ][ 280 ],
   alphaCSR[ 56 ][ 281 ],
   alphaCSR[ 56 ][ 282 ],
   alphaCSR[ 56 ][ 283 ],
   alphaCSR[ 56 ][ 284 ],
   alphaCSR[ 56 ][ 285 ],
   alphaCSR[ 56 ][ 286 ],
   alphaCSR[ 56 ][ 287 ],
   alphaCSR[ 56 ][ 288 ],
   alphaCSR[ 56 ][ 289 ],
   alphaCSR[ 56 ][ 290 ],
   alphaCSR[ 56 ][ 291 ],
   alphaCSR[ 56 ][ 292 ],
   alphaCSR[ 56 ][ 293 ],
   alphaCSR[ 56 ][ 294 ],
   alphaCSR[ 56 ][ 295 ],
   alphaCSR[ 56 ][ 296 ],
   alphaCSR[ 56 ][ 297 ],
   alphaCSR[ 56 ][ 298 ],
   alphaCSR[ 56 ][ 299 ],
   alphaCSR[ 56 ][ 300 ],
   alphaCSR[ 56 ][ 301 ],
   alphaCSR[ 56 ][ 302 ],
   alphaCSR[ 56 ][ 303 ],
   alphaCSR[ 56 ][ 304 ],
   alphaCSR[ 56 ][ 305 ],
   alphaCSR[ 56 ][ 306 ],
   alphaCSR[ 56 ][ 307 ],
   alphaCSR[ 56 ][ 308 ],
   alphaCSR[ 56 ][ 309 ],
   alphaCSR[ 56 ][ 310 ],
   alphaCSR[ 56 ][ 311 ],
   alphaCSR[ 56 ][ 312 ],
   alphaCSR[ 56 ][ 313 ],
   alphaCSR[ 56 ][ 314 ],
   alphaCSR[ 56 ][ 315 ],
   alphaCSR[ 56 ][ 316 ],
   alphaCSR[ 56 ][ 317 ],
   alphaCSR[ 56 ][ 318 ],
   alphaCSR[ 56 ][ 319 ],
   alphaCSR[ 56 ][ 320 ],
   alphaCSR[ 56 ][ 321 ],
   alphaCSR[ 56 ][ 322 ],
   alphaCSR[ 56 ][ 323 ],
   alphaCSR[ 56 ][ 324 ],
   alphaCSR[ 56 ][ 325 ],
   alphaCSR[ 56 ][ 326 ],
   alphaCSR[ 56 ][ 327 ],
   alphaCSR[ 56 ][ 328 ],
   alphaCSR[ 56 ][ 329 ],
   alphaCSR[ 56 ][ 330 ],
   alphaCSR[ 56 ][ 331 ],
   alphaCSR[ 56 ][ 332 ],
   alphaCSR[ 56 ][ 333 ],
   alphaCSR[ 56 ][ 334 ],
   alphaCSR[ 56 ][ 335 ],
   alphaCSR[ 56 ][ 336 ],
   alphaCSR[ 56 ][ 337 ],
   alphaCSR[ 56 ][ 338 ],
   alphaCSR[ 56 ][ 339 ],
   alphaCSR[ 56 ][ 340 ],
   alphaCSR[ 56 ][ 341 ],
   alphaCSR[ 56 ][ 342 ],
   alphaCSR[ 56 ][ 343 ],
   alphaCSR[ 56 ][ 344 ],
   alphaCSR[ 56 ][ 345 ],
   alphaCSR[ 56 ][ 346 ],
   alphaCSR[ 56 ][ 347 ],
   alphaCSR[ 56 ][ 348 ],
   alphaCSR[ 56 ][ 349 ],
   alphaCSR[ 56 ][ 350 ],
   alphaCSR[ 56 ][ 351 ],
   alphaCSR[ 56 ][ 352 ],
   alphaCSR[ 56 ][ 353 ],
   alphaCSR[ 56 ][ 354 ],
   alphaCSR[ 56 ][ 355 ],
   alphaCSR[ 56 ][ 356 ],
   alphaCSR[ 56 ][ 357 ],
   alphaCSR[ 56 ][ 358 ],
   alphaCSR[ 56 ][ 359 ],
   alphaCSR[ 56 ][ 360 ],
   alphaCSR[ 56 ][ 361 ],
   alphaCSR[ 56 ][ 362 ],
   alphaCSR[ 56 ][ 363 ],
   alphaCSR[ 56 ][ 364 ],
   alphaCSR[ 56 ][ 365 ],
   alphaCSR[ 56 ][ 366 ],
   alphaCSR[ 56 ][ 367 ],
   alphaCSR[ 56 ][ 368 ],
   alphaCSR[ 56 ][ 369 ],
   alphaCSR[ 56 ][ 370 ],
   alphaCSR[ 56 ][ 371 ],
   alphaCSR[ 56 ][ 372 ],
   alphaCSR[ 56 ][ 373 ],
   alphaCSR[ 56 ][ 374 ],
   alphaCSR[ 56 ][ 375 ],
   alphaCSR[ 56 ][ 376 ],
   alphaCSR[ 56 ][ 377 ],
   alphaCSR[ 56 ][ 378 ],
   alphaCSR[ 56 ][ 379 ],
   alphaCSR[ 56 ][ 380 ],
   alphaCSR[ 56 ][ 381 ],
   alphaCSR[ 56 ][ 382 ],
   alphaCSR[ 56 ][ 383 ],
   alphaCSR[ 57 ][ 0 ],
   alphaCSR[ 57 ][ 1 ],
   alphaCSR[ 57 ][ 2 ],
   alphaCSR[ 57 ][ 3 ],
   alphaCSR[ 57 ][ 4 ],
   alphaCSR[ 57 ][ 5 ],
   alphaCSR[ 57 ][ 6 ],
   alphaCSR[ 57 ][ 7 ],
   alphaCSR[ 57 ][ 8 ],
   alphaCSR[ 57 ][ 9 ],
   alphaCSR[ 57 ][ 10 ],
   alphaCSR[ 57 ][ 11 ],
   alphaCSR[ 57 ][ 12 ],
   alphaCSR[ 57 ][ 13 ],
   alphaCSR[ 57 ][ 14 ],
   alphaCSR[ 57 ][ 15 ],
   alphaCSR[ 57 ][ 16 ],
   alphaCSR[ 57 ][ 17 ],
   alphaCSR[ 57 ][ 18 ],
   alphaCSR[ 57 ][ 19 ],
   alphaCSR[ 57 ][ 20 ],
   alphaCSR[ 57 ][ 21 ],
   alphaCSR[ 57 ][ 22 ],
   alphaCSR[ 57 ][ 23 ],
   alphaCSR[ 57 ][ 24 ],
   alphaCSR[ 57 ][ 25 ],
   alphaCSR[ 57 ][ 26 ],
   alphaCSR[ 57 ][ 27 ],
   alphaCSR[ 57 ][ 28 ],
   alphaCSR[ 57 ][ 29 ],
   alphaCSR[ 57 ][ 30 ],
   alphaCSR[ 57 ][ 31 ],
   alphaCSR[ 57 ][ 32 ],
   alphaCSR[ 57 ][ 33 ],
   alphaCSR[ 57 ][ 34 ],
   alphaCSR[ 57 ][ 35 ],
   alphaCSR[ 57 ][ 36 ],
   alphaCSR[ 57 ][ 37 ],
   alphaCSR[ 57 ][ 38 ],
   alphaCSR[ 57 ][ 39 ],
   alphaCSR[ 57 ][ 40 ],
   alphaCSR[ 57 ][ 41 ],
   alphaCSR[ 57 ][ 42 ],
   alphaCSR[ 57 ][ 43 ],
   alphaCSR[ 57 ][ 44 ],
   alphaCSR[ 57 ][ 45 ],
   alphaCSR[ 57 ][ 46 ],
   alphaCSR[ 57 ][ 47 ],
   alphaCSR[ 57 ][ 48 ],
   alphaCSR[ 57 ][ 49 ],
   alphaCSR[ 57 ][ 50 ],
   alphaCSR[ 57 ][ 51 ],
   alphaCSR[ 57 ][ 52 ],
   alphaCSR[ 57 ][ 53 ],
   alphaCSR[ 57 ][ 54 ],
   alphaCSR[ 57 ][ 55 ],
   alphaCSR[ 57 ][ 56 ],
   alphaCSR[ 57 ][ 57 ],
   alphaCSR[ 57 ][ 58 ],
   alphaCSR[ 57 ][ 59 ],
   alphaCSR[ 57 ][ 60 ],
   alphaCSR[ 57 ][ 61 ],
   alphaCSR[ 57 ][ 62 ],
   alphaCSR[ 57 ][ 63 ],
   alphaCSR[ 57 ][ 64 ],
   alphaCSR[ 57 ][ 65 ],
   alphaCSR[ 57 ][ 66 ],
   alphaCSR[ 57 ][ 67 ],
   alphaCSR[ 57 ][ 68 ],
   alphaCSR[ 57 ][ 69 ],
   alphaCSR[ 57 ][ 70 ],
   alphaCSR[ 57 ][ 71 ],
   alphaCSR[ 57 ][ 72 ],
   alphaCSR[ 57 ][ 73 ],
   alphaCSR[ 57 ][ 74 ],
   alphaCSR[ 57 ][ 75 ],
   alphaCSR[ 57 ][ 76 ],
   alphaCSR[ 57 ][ 77 ],
   alphaCSR[ 57 ][ 78 ],
   alphaCSR[ 57 ][ 79 ],
   alphaCSR[ 57 ][ 80 ],
   alphaCSR[ 57 ][ 81 ],
   alphaCSR[ 57 ][ 82 ],
   alphaCSR[ 57 ][ 83 ],
   alphaCSR[ 57 ][ 84 ],
   alphaCSR[ 57 ][ 85 ],
   alphaCSR[ 57 ][ 86 ],
   alphaCSR[ 57 ][ 87 ],
   alphaCSR[ 57 ][ 88 ],
   alphaCSR[ 57 ][ 89 ],
   alphaCSR[ 57 ][ 90 ],
   alphaCSR[ 57 ][ 91 ],
   alphaCSR[ 57 ][ 92 ],
   alphaCSR[ 57 ][ 93 ],
   alphaCSR[ 57 ][ 94 ],
   alphaCSR[ 57 ][ 95 ],
   alphaCSR[ 57 ][ 96 ],
   alphaCSR[ 57 ][ 97 ],
   alphaCSR[ 57 ][ 98 ],
   alphaCSR[ 57 ][ 99 ],
   alphaCSR[ 57 ][ 100 ],
   alphaCSR[ 57 ][ 101 ],
   alphaCSR[ 57 ][ 102 ],
   alphaCSR[ 57 ][ 103 ],
   alphaCSR[ 57 ][ 104 ],
   alphaCSR[ 57 ][ 105 ],
   alphaCSR[ 57 ][ 106 ],
   alphaCSR[ 57 ][ 107 ],
   alphaCSR[ 57 ][ 108 ],
   alphaCSR[ 57 ][ 109 ],
   alphaCSR[ 57 ][ 110 ],
   alphaCSR[ 57 ][ 111 ],
   alphaCSR[ 57 ][ 112 ],
   alphaCSR[ 57 ][ 113 ],
   alphaCSR[ 57 ][ 114 ],
   alphaCSR[ 57 ][ 115 ],
   alphaCSR[ 57 ][ 116 ],
   alphaCSR[ 57 ][ 117 ],
   alphaCSR[ 57 ][ 118 ],
   alphaCSR[ 57 ][ 119 ],
   alphaCSR[ 57 ][ 120 ],
   alphaCSR[ 57 ][ 121 ],
   alphaCSR[ 57 ][ 122 ],
   alphaCSR[ 57 ][ 123 ],
   alphaCSR[ 57 ][ 124 ],
   alphaCSR[ 57 ][ 125 ],
   alphaCSR[ 57 ][ 126 ],
   alphaCSR[ 57 ][ 127 ],
   alphaCSR[ 57 ][ 128 ],
   alphaCSR[ 57 ][ 129 ],
   alphaCSR[ 57 ][ 130 ],
   alphaCSR[ 57 ][ 131 ],
   alphaCSR[ 57 ][ 132 ],
   alphaCSR[ 57 ][ 133 ],
   alphaCSR[ 57 ][ 134 ],
   alphaCSR[ 57 ][ 135 ],
   alphaCSR[ 57 ][ 136 ],
   alphaCSR[ 57 ][ 137 ],
   alphaCSR[ 57 ][ 138 ],
   alphaCSR[ 57 ][ 139 ],
   alphaCSR[ 57 ][ 140 ],
   alphaCSR[ 57 ][ 141 ],
   alphaCSR[ 57 ][ 142 ],
   alphaCSR[ 57 ][ 143 ],
   alphaCSR[ 57 ][ 144 ],
   alphaCSR[ 57 ][ 145 ],
   alphaCSR[ 57 ][ 146 ],
   alphaCSR[ 57 ][ 147 ],
   alphaCSR[ 57 ][ 148 ],
   alphaCSR[ 57 ][ 149 ],
   alphaCSR[ 57 ][ 150 ],
   alphaCSR[ 57 ][ 151 ],
   alphaCSR[ 57 ][ 152 ],
   alphaCSR[ 57 ][ 153 ],
   alphaCSR[ 57 ][ 154 ],
   alphaCSR[ 57 ][ 155 ],
   alphaCSR[ 57 ][ 156 ],
   alphaCSR[ 57 ][ 157 ],
   alphaCSR[ 57 ][ 158 ],
   alphaCSR[ 57 ][ 159 ],
   alphaCSR[ 57 ][ 160 ],
   alphaCSR[ 57 ][ 161 ],
   alphaCSR[ 57 ][ 162 ],
   alphaCSR[ 57 ][ 163 ],
   alphaCSR[ 57 ][ 164 ],
   alphaCSR[ 57 ][ 165 ],
   alphaCSR[ 57 ][ 166 ],
   alphaCSR[ 57 ][ 167 ],
   alphaCSR[ 57 ][ 168 ],
   alphaCSR[ 57 ][ 169 ],
   alphaCSR[ 57 ][ 170 ],
   alphaCSR[ 57 ][ 171 ],
   alphaCSR[ 57 ][ 172 ],
   alphaCSR[ 57 ][ 173 ],
   alphaCSR[ 57 ][ 174 ],
   alphaCSR[ 57 ][ 175 ],
   alphaCSR[ 57 ][ 176 ],
   alphaCSR[ 57 ][ 177 ],
   alphaCSR[ 57 ][ 178 ],
   alphaCSR[ 57 ][ 179 ],
   alphaCSR[ 57 ][ 180 ],
   alphaCSR[ 57 ][ 181 ],
   alphaCSR[ 57 ][ 182 ],
   alphaCSR[ 57 ][ 183 ],
   alphaCSR[ 57 ][ 184 ],
   alphaCSR[ 57 ][ 185 ],
   alphaCSR[ 57 ][ 186 ],
   alphaCSR[ 57 ][ 187 ],
   alphaCSR[ 57 ][ 188 ],
   alphaCSR[ 57 ][ 189 ],
   alphaCSR[ 57 ][ 190 ],
   alphaCSR[ 57 ][ 191 ],
   alphaCSR[ 57 ][ 192 ],
   alphaCSR[ 57 ][ 193 ],
   alphaCSR[ 57 ][ 194 ],
   alphaCSR[ 57 ][ 195 ],
   alphaCSR[ 57 ][ 196 ],
   alphaCSR[ 57 ][ 197 ],
   alphaCSR[ 57 ][ 198 ],
   alphaCSR[ 57 ][ 199 ],
   alphaCSR[ 57 ][ 200 ],
   alphaCSR[ 57 ][ 201 ],
   alphaCSR[ 57 ][ 202 ],
   alphaCSR[ 57 ][ 203 ],
   alphaCSR[ 57 ][ 204 ],
   alphaCSR[ 57 ][ 205 ],
   alphaCSR[ 57 ][ 206 ],
   alphaCSR[ 57 ][ 207 ],
   alphaCSR[ 57 ][ 208 ],
   alphaCSR[ 57 ][ 209 ],
   alphaCSR[ 57 ][ 210 ],
   alphaCSR[ 57 ][ 211 ],
   alphaCSR[ 57 ][ 212 ],
   alphaCSR[ 57 ][ 213 ],
   alphaCSR[ 57 ][ 214 ],
   alphaCSR[ 57 ][ 215 ],
   alphaCSR[ 57 ][ 216 ],
   alphaCSR[ 57 ][ 217 ],
   alphaCSR[ 57 ][ 218 ],
   alphaCSR[ 57 ][ 219 ],
   alphaCSR[ 57 ][ 220 ],
   alphaCSR[ 57 ][ 221 ],
   alphaCSR[ 57 ][ 222 ],
   alphaCSR[ 57 ][ 223 ],
   alphaCSR[ 57 ][ 224 ],
   alphaCSR[ 57 ][ 225 ],
   alphaCSR[ 57 ][ 226 ],
   alphaCSR[ 57 ][ 227 ],
   alphaCSR[ 57 ][ 228 ],
   alphaCSR[ 57 ][ 229 ],
   alphaCSR[ 57 ][ 230 ],
   alphaCSR[ 57 ][ 231 ],
   alphaCSR[ 57 ][ 232 ],
   alphaCSR[ 57 ][ 233 ],
   alphaCSR[ 57 ][ 234 ],
   alphaCSR[ 57 ][ 235 ],
   alphaCSR[ 57 ][ 236 ],
   alphaCSR[ 57 ][ 237 ],
   alphaCSR[ 57 ][ 238 ],
   alphaCSR[ 57 ][ 239 ],
   alphaCSR[ 57 ][ 240 ],
   alphaCSR[ 57 ][ 241 ],
   alphaCSR[ 57 ][ 242 ],
   alphaCSR[ 57 ][ 243 ],
   alphaCSR[ 57 ][ 244 ],
   alphaCSR[ 57 ][ 245 ],
   alphaCSR[ 57 ][ 246 ],
   alphaCSR[ 57 ][ 247 ],
   alphaCSR[ 57 ][ 248 ],
   alphaCSR[ 57 ][ 249 ],
   alphaCSR[ 57 ][ 250 ],
   alphaCSR[ 57 ][ 251 ],
   alphaCSR[ 57 ][ 252 ],
   alphaCSR[ 57 ][ 253 ],
   alphaCSR[ 57 ][ 254 ],
   alphaCSR[ 57 ][ 255 ],
   alphaCSR[ 57 ][ 256 ],
   alphaCSR[ 57 ][ 257 ],
   alphaCSR[ 57 ][ 258 ],
   alphaCSR[ 57 ][ 259 ],
   alphaCSR[ 57 ][ 260 ],
   alphaCSR[ 57 ][ 261 ],
   alphaCSR[ 57 ][ 262 ],
   alphaCSR[ 57 ][ 263 ],
   alphaCSR[ 57 ][ 264 ],
   alphaCSR[ 57 ][ 265 ],
   alphaCSR[ 57 ][ 266 ],
   alphaCSR[ 57 ][ 267 ],
   alphaCSR[ 57 ][ 268 ],
   alphaCSR[ 57 ][ 269 ],
   alphaCSR[ 57 ][ 270 ],
   alphaCSR[ 57 ][ 271 ],
   alphaCSR[ 57 ][ 272 ],
   alphaCSR[ 57 ][ 273 ],
   alphaCSR[ 57 ][ 274 ],
   alphaCSR[ 57 ][ 275 ],
   alphaCSR[ 57 ][ 276 ],
   alphaCSR[ 57 ][ 277 ],
   alphaCSR[ 57 ][ 278 ],
   alphaCSR[ 57 ][ 279 ],
   alphaCSR[ 57 ][ 280 ],
   alphaCSR[ 57 ][ 281 ],
   alphaCSR[ 57 ][ 282 ],
   alphaCSR[ 57 ][ 283 ],
   alphaCSR[ 57 ][ 284 ],
   alphaCSR[ 57 ][ 285 ],
   alphaCSR[ 57 ][ 286 ],
   alphaCSR[ 57 ][ 287 ],
   alphaCSR[ 57 ][ 288 ],
   alphaCSR[ 57 ][ 289 ],
   alphaCSR[ 57 ][ 290 ],
   alphaCSR[ 57 ][ 291 ],
   alphaCSR[ 57 ][ 292 ],
   alphaCSR[ 57 ][ 293 ],
   alphaCSR[ 57 ][ 294 ],
   alphaCSR[ 57 ][ 295 ],
   alphaCSR[ 57 ][ 296 ],
   alphaCSR[ 57 ][ 297 ],
   alphaCSR[ 57 ][ 298 ],
   alphaCSR[ 57 ][ 299 ],
   alphaCSR[ 57 ][ 300 ],
   alphaCSR[ 57 ][ 301 ],
   alphaCSR[ 57 ][ 302 ],
   alphaCSR[ 57 ][ 303 ],
   alphaCSR[ 57 ][ 304 ],
   alphaCSR[ 57 ][ 305 ],
   alphaCSR[ 57 ][ 306 ],
   alphaCSR[ 57 ][ 307 ],
   alphaCSR[ 57 ][ 308 ],
   alphaCSR[ 57 ][ 309 ],
   alphaCSR[ 57 ][ 310 ],
   alphaCSR[ 57 ][ 311 ],
   alphaCSR[ 57 ][ 312 ],
   alphaCSR[ 57 ][ 313 ],
   alphaCSR[ 57 ][ 314 ],
   alphaCSR[ 57 ][ 315 ],
   alphaCSR[ 57 ][ 316 ],
   alphaCSR[ 57 ][ 317 ],
   alphaCSR[ 57 ][ 318 ],
   alphaCSR[ 57 ][ 319 ],
   alphaCSR[ 57 ][ 320 ],
   alphaCSR[ 57 ][ 321 ],
   alphaCSR[ 57 ][ 322 ],
   alphaCSR[ 57 ][ 323 ],
   alphaCSR[ 57 ][ 324 ],
   alphaCSR[ 57 ][ 325 ],
   alphaCSR[ 57 ][ 326 ],
   alphaCSR[ 57 ][ 327 ],
   alphaCSR[ 57 ][ 328 ],
   alphaCSR[ 57 ][ 329 ],
   alphaCSR[ 57 ][ 330 ],
   alphaCSR[ 57 ][ 331 ],
   alphaCSR[ 57 ][ 332 ],
   alphaCSR[ 57 ][ 333 ],
   alphaCSR[ 57 ][ 334 ],
   alphaCSR[ 57 ][ 335 ],
   alphaCSR[ 57 ][ 336 ],
   alphaCSR[ 57 ][ 337 ],
   alphaCSR[ 57 ][ 338 ],
   alphaCSR[ 57 ][ 339 ],
   alphaCSR[ 57 ][ 340 ],
   alphaCSR[ 57 ][ 341 ],
   alphaCSR[ 57 ][ 342 ],
   alphaCSR[ 57 ][ 343 ],
   alphaCSR[ 57 ][ 344 ],
   alphaCSR[ 57 ][ 345 ],
   alphaCSR[ 57 ][ 346 ],
   alphaCSR[ 57 ][ 347 ],
   alphaCSR[ 57 ][ 348 ],
   alphaCSR[ 57 ][ 349 ],
   alphaCSR[ 57 ][ 350 ],
   alphaCSR[ 57 ][ 351 ],
   alphaCSR[ 57 ][ 352 ],
   alphaCSR[ 57 ][ 353 ],
   alphaCSR[ 57 ][ 354 ],
   alphaCSR[ 57 ][ 355 ],
   alphaCSR[ 57 ][ 356 ],
   alphaCSR[ 57 ][ 357 ],
   alphaCSR[ 57 ][ 358 ],
   alphaCSR[ 57 ][ 359 ],
   alphaCSR[ 57 ][ 360 ],
   alphaCSR[ 57 ][ 361 ],
   alphaCSR[ 57 ][ 362 ],
   alphaCSR[ 57 ][ 363 ],
   alphaCSR[ 57 ][ 364 ],
   alphaCSR[ 57 ][ 365 ],
   alphaCSR[ 57 ][ 366 ],
   alphaCSR[ 57 ][ 367 ],
   alphaCSR[ 57 ][ 368 ],
   alphaCSR[ 57 ][ 369 ],
   alphaCSR[ 57 ][ 370 ],
   alphaCSR[ 57 ][ 371 ],
   alphaCSR[ 57 ][ 372 ],
   alphaCSR[ 57 ][ 373 ],
   alphaCSR[ 57 ][ 374 ],
   alphaCSR[ 57 ][ 375 ],
   alphaCSR[ 57 ][ 376 ],
   alphaCSR[ 57 ][ 377 ],
   alphaCSR[ 57 ][ 378 ],
   alphaCSR[ 57 ][ 379 ],
   alphaCSR[ 57 ][ 380 ],
   alphaCSR[ 57 ][ 381 ],
   alphaCSR[ 57 ][ 382 ],
   alphaCSR[ 57 ][ 383 ],
   alphaCSR[ 58 ][ 0 ],
   alphaCSR[ 58 ][ 1 ],
   alphaCSR[ 58 ][ 2 ],
   alphaCSR[ 58 ][ 3 ],
   alphaCSR[ 58 ][ 4 ],
   alphaCSR[ 58 ][ 5 ],
   alphaCSR[ 58 ][ 6 ],
   alphaCSR[ 58 ][ 7 ],
   alphaCSR[ 58 ][ 8 ],
   alphaCSR[ 58 ][ 9 ],
   alphaCSR[ 58 ][ 10 ],
   alphaCSR[ 58 ][ 11 ],
   alphaCSR[ 58 ][ 12 ],
   alphaCSR[ 58 ][ 13 ],
   alphaCSR[ 58 ][ 14 ],
   alphaCSR[ 58 ][ 15 ],
   alphaCSR[ 58 ][ 16 ],
   alphaCSR[ 58 ][ 17 ],
   alphaCSR[ 58 ][ 18 ],
   alphaCSR[ 58 ][ 19 ],
   alphaCSR[ 58 ][ 20 ],
   alphaCSR[ 58 ][ 21 ],
   alphaCSR[ 58 ][ 22 ],
   alphaCSR[ 58 ][ 23 ],
   alphaCSR[ 58 ][ 24 ],
   alphaCSR[ 58 ][ 25 ],
   alphaCSR[ 58 ][ 26 ],
   alphaCSR[ 58 ][ 27 ],
   alphaCSR[ 58 ][ 28 ],
   alphaCSR[ 58 ][ 29 ],
   alphaCSR[ 58 ][ 30 ],
   alphaCSR[ 58 ][ 31 ],
   alphaCSR[ 58 ][ 32 ],
   alphaCSR[ 58 ][ 33 ],
   alphaCSR[ 58 ][ 34 ],
   alphaCSR[ 58 ][ 35 ],
   alphaCSR[ 58 ][ 36 ],
   alphaCSR[ 58 ][ 37 ],
   alphaCSR[ 58 ][ 38 ],
   alphaCSR[ 58 ][ 39 ],
   alphaCSR[ 58 ][ 40 ],
   alphaCSR[ 58 ][ 41 ],
   alphaCSR[ 58 ][ 42 ],
   alphaCSR[ 58 ][ 43 ],
   alphaCSR[ 58 ][ 44 ],
   alphaCSR[ 58 ][ 45 ],
   alphaCSR[ 58 ][ 46 ],
   alphaCSR[ 58 ][ 47 ],
   alphaCSR[ 58 ][ 48 ],
   alphaCSR[ 58 ][ 49 ],
   alphaCSR[ 58 ][ 50 ],
   alphaCSR[ 58 ][ 51 ],
   alphaCSR[ 58 ][ 52 ],
   alphaCSR[ 58 ][ 53 ],
   alphaCSR[ 58 ][ 54 ],
   alphaCSR[ 58 ][ 55 ],
   alphaCSR[ 58 ][ 56 ],
   alphaCSR[ 58 ][ 57 ],
   alphaCSR[ 58 ][ 58 ],
   alphaCSR[ 58 ][ 59 ],
   alphaCSR[ 58 ][ 60 ],
   alphaCSR[ 58 ][ 61 ],
   alphaCSR[ 58 ][ 62 ],
   alphaCSR[ 58 ][ 63 ],
   alphaCSR[ 58 ][ 64 ],
   alphaCSR[ 58 ][ 65 ],
   alphaCSR[ 58 ][ 66 ],
   alphaCSR[ 58 ][ 67 ],
   alphaCSR[ 58 ][ 68 ],
   alphaCSR[ 58 ][ 69 ],
   alphaCSR[ 58 ][ 70 ],
   alphaCSR[ 58 ][ 71 ],
   alphaCSR[ 58 ][ 72 ],
   alphaCSR[ 58 ][ 73 ],
   alphaCSR[ 58 ][ 74 ],
   alphaCSR[ 58 ][ 75 ],
   alphaCSR[ 58 ][ 76 ],
   alphaCSR[ 58 ][ 77 ],
   alphaCSR[ 58 ][ 78 ],
   alphaCSR[ 58 ][ 79 ],
   alphaCSR[ 58 ][ 80 ],
   alphaCSR[ 58 ][ 81 ],
   alphaCSR[ 58 ][ 82 ],
   alphaCSR[ 58 ][ 83 ],
   alphaCSR[ 58 ][ 84 ],
   alphaCSR[ 58 ][ 85 ],
   alphaCSR[ 58 ][ 86 ],
   alphaCSR[ 58 ][ 87 ],
   alphaCSR[ 58 ][ 88 ],
   alphaCSR[ 58 ][ 89 ],
   alphaCSR[ 58 ][ 90 ],
   alphaCSR[ 58 ][ 91 ],
   alphaCSR[ 58 ][ 92 ],
   alphaCSR[ 58 ][ 93 ],
   alphaCSR[ 58 ][ 94 ],
   alphaCSR[ 58 ][ 95 ],
   alphaCSR[ 58 ][ 96 ],
   alphaCSR[ 58 ][ 97 ],
   alphaCSR[ 58 ][ 98 ],
   alphaCSR[ 58 ][ 99 ],
   alphaCSR[ 58 ][ 100 ],
   alphaCSR[ 58 ][ 101 ],
   alphaCSR[ 58 ][ 102 ],
   alphaCSR[ 58 ][ 103 ],
   alphaCSR[ 58 ][ 104 ],
   alphaCSR[ 58 ][ 105 ],
   alphaCSR[ 58 ][ 106 ],
   alphaCSR[ 58 ][ 107 ],
   alphaCSR[ 58 ][ 108 ],
   alphaCSR[ 58 ][ 109 ],
   alphaCSR[ 58 ][ 110 ],
   alphaCSR[ 58 ][ 111 ],
   alphaCSR[ 58 ][ 112 ],
   alphaCSR[ 58 ][ 113 ],
   alphaCSR[ 58 ][ 114 ],
   alphaCSR[ 58 ][ 115 ],
   alphaCSR[ 58 ][ 116 ],
   alphaCSR[ 58 ][ 117 ],
   alphaCSR[ 58 ][ 118 ],
   alphaCSR[ 58 ][ 119 ],
   alphaCSR[ 58 ][ 120 ],
   alphaCSR[ 58 ][ 121 ],
   alphaCSR[ 58 ][ 122 ],
   alphaCSR[ 58 ][ 123 ],
   alphaCSR[ 58 ][ 124 ],
   alphaCSR[ 58 ][ 125 ],
   alphaCSR[ 58 ][ 126 ],
   alphaCSR[ 58 ][ 127 ],
   alphaCSR[ 58 ][ 128 ],
   alphaCSR[ 58 ][ 129 ],
   alphaCSR[ 58 ][ 130 ],
   alphaCSR[ 58 ][ 131 ],
   alphaCSR[ 58 ][ 132 ],
   alphaCSR[ 58 ][ 133 ],
   alphaCSR[ 58 ][ 134 ],
   alphaCSR[ 58 ][ 135 ],
   alphaCSR[ 58 ][ 136 ],
   alphaCSR[ 58 ][ 137 ],
   alphaCSR[ 58 ][ 138 ],
   alphaCSR[ 58 ][ 139 ],
   alphaCSR[ 58 ][ 140 ],
   alphaCSR[ 58 ][ 141 ],
   alphaCSR[ 58 ][ 142 ],
   alphaCSR[ 58 ][ 143 ],
   alphaCSR[ 58 ][ 144 ],
   alphaCSR[ 58 ][ 145 ],
   alphaCSR[ 58 ][ 146 ],
   alphaCSR[ 58 ][ 147 ],
   alphaCSR[ 58 ][ 148 ],
   alphaCSR[ 58 ][ 149 ],
   alphaCSR[ 58 ][ 150 ],
   alphaCSR[ 58 ][ 151 ],
   alphaCSR[ 58 ][ 152 ],
   alphaCSR[ 58 ][ 153 ],
   alphaCSR[ 58 ][ 154 ],
   alphaCSR[ 58 ][ 155 ],
   alphaCSR[ 58 ][ 156 ],
   alphaCSR[ 58 ][ 157 ],
   alphaCSR[ 58 ][ 158 ],
   alphaCSR[ 58 ][ 159 ],
   alphaCSR[ 58 ][ 160 ],
   alphaCSR[ 58 ][ 161 ],
   alphaCSR[ 58 ][ 162 ],
   alphaCSR[ 58 ][ 163 ],
   alphaCSR[ 58 ][ 164 ],
   alphaCSR[ 58 ][ 165 ],
   alphaCSR[ 58 ][ 166 ],
   alphaCSR[ 58 ][ 167 ],
   alphaCSR[ 58 ][ 168 ],
   alphaCSR[ 58 ][ 169 ],
   alphaCSR[ 58 ][ 170 ],
   alphaCSR[ 58 ][ 171 ],
   alphaCSR[ 58 ][ 172 ],
   alphaCSR[ 58 ][ 173 ],
   alphaCSR[ 58 ][ 174 ],
   alphaCSR[ 58 ][ 175 ],
   alphaCSR[ 58 ][ 176 ],
   alphaCSR[ 58 ][ 177 ],
   alphaCSR[ 58 ][ 178 ],
   alphaCSR[ 58 ][ 179 ],
   alphaCSR[ 58 ][ 180 ],
   alphaCSR[ 58 ][ 181 ],
   alphaCSR[ 58 ][ 182 ],
   alphaCSR[ 58 ][ 183 ],
   alphaCSR[ 58 ][ 184 ],
   alphaCSR[ 58 ][ 185 ],
   alphaCSR[ 58 ][ 186 ],
   alphaCSR[ 58 ][ 187 ],
   alphaCSR[ 58 ][ 188 ],
   alphaCSR[ 58 ][ 189 ],
   alphaCSR[ 58 ][ 190 ],
   alphaCSR[ 58 ][ 191 ],
   alphaCSR[ 58 ][ 192 ],
   alphaCSR[ 58 ][ 193 ],
   alphaCSR[ 58 ][ 194 ],
   alphaCSR[ 58 ][ 195 ],
   alphaCSR[ 58 ][ 196 ],
   alphaCSR[ 58 ][ 197 ],
   alphaCSR[ 58 ][ 198 ],
   alphaCSR[ 58 ][ 199 ],
   alphaCSR[ 58 ][ 200 ],
   alphaCSR[ 58 ][ 201 ],
   alphaCSR[ 58 ][ 202 ],
   alphaCSR[ 58 ][ 203 ],
   alphaCSR[ 58 ][ 204 ],
   alphaCSR[ 58 ][ 205 ],
   alphaCSR[ 58 ][ 206 ],
   alphaCSR[ 58 ][ 207 ],
   alphaCSR[ 58 ][ 208 ],
   alphaCSR[ 58 ][ 209 ],
   alphaCSR[ 58 ][ 210 ],
   alphaCSR[ 58 ][ 211 ],
   alphaCSR[ 58 ][ 212 ],
   alphaCSR[ 58 ][ 213 ],
   alphaCSR[ 58 ][ 214 ],
   alphaCSR[ 58 ][ 215 ],
   alphaCSR[ 58 ][ 216 ],
   alphaCSR[ 58 ][ 217 ],
   alphaCSR[ 58 ][ 218 ],
   alphaCSR[ 58 ][ 219 ],
   alphaCSR[ 58 ][ 220 ],
   alphaCSR[ 58 ][ 221 ],
   alphaCSR[ 58 ][ 222 ],
   alphaCSR[ 58 ][ 223 ],
   alphaCSR[ 58 ][ 224 ],
   alphaCSR[ 58 ][ 225 ],
   alphaCSR[ 58 ][ 226 ],
   alphaCSR[ 58 ][ 227 ],
   alphaCSR[ 58 ][ 228 ],
   alphaCSR[ 58 ][ 229 ],
   alphaCSR[ 58 ][ 230 ],
   alphaCSR[ 58 ][ 231 ],
   alphaCSR[ 58 ][ 232 ],
   alphaCSR[ 58 ][ 233 ],
   alphaCSR[ 58 ][ 234 ],
   alphaCSR[ 58 ][ 235 ],
   alphaCSR[ 58 ][ 236 ],
   alphaCSR[ 58 ][ 237 ],
   alphaCSR[ 58 ][ 238 ],
   alphaCSR[ 58 ][ 239 ],
   alphaCSR[ 58 ][ 240 ],
   alphaCSR[ 58 ][ 241 ],
   alphaCSR[ 58 ][ 242 ],
   alphaCSR[ 58 ][ 243 ],
   alphaCSR[ 58 ][ 244 ],
   alphaCSR[ 58 ][ 245 ],
   alphaCSR[ 58 ][ 246 ],
   alphaCSR[ 58 ][ 247 ],
   alphaCSR[ 58 ][ 248 ],
   alphaCSR[ 58 ][ 249 ],
   alphaCSR[ 58 ][ 250 ],
   alphaCSR[ 58 ][ 251 ],
   alphaCSR[ 58 ][ 252 ],
   alphaCSR[ 58 ][ 253 ],
   alphaCSR[ 58 ][ 254 ],
   alphaCSR[ 58 ][ 255 ],
   alphaCSR[ 58 ][ 256 ],
   alphaCSR[ 58 ][ 257 ],
   alphaCSR[ 58 ][ 258 ],
   alphaCSR[ 58 ][ 259 ],
   alphaCSR[ 58 ][ 260 ],
   alphaCSR[ 58 ][ 261 ],
   alphaCSR[ 58 ][ 262 ],
   alphaCSR[ 58 ][ 263 ],
   alphaCSR[ 58 ][ 264 ],
   alphaCSR[ 58 ][ 265 ],
   alphaCSR[ 58 ][ 266 ],
   alphaCSR[ 58 ][ 267 ],
   alphaCSR[ 58 ][ 268 ],
   alphaCSR[ 58 ][ 269 ],
   alphaCSR[ 58 ][ 270 ],
   alphaCSR[ 58 ][ 271 ],
   alphaCSR[ 58 ][ 272 ],
   alphaCSR[ 58 ][ 273 ],
   alphaCSR[ 58 ][ 274 ],
   alphaCSR[ 58 ][ 275 ],
   alphaCSR[ 58 ][ 276 ],
   alphaCSR[ 58 ][ 277 ],
   alphaCSR[ 58 ][ 278 ],
   alphaCSR[ 58 ][ 279 ],
   alphaCSR[ 58 ][ 280 ],
   alphaCSR[ 58 ][ 281 ],
   alphaCSR[ 58 ][ 282 ],
   alphaCSR[ 58 ][ 283 ],
   alphaCSR[ 58 ][ 284 ],
   alphaCSR[ 58 ][ 285 ],
   alphaCSR[ 58 ][ 286 ],
   alphaCSR[ 58 ][ 287 ],
   alphaCSR[ 58 ][ 288 ],
   alphaCSR[ 58 ][ 289 ],
   alphaCSR[ 58 ][ 290 ],
   alphaCSR[ 58 ][ 291 ],
   alphaCSR[ 58 ][ 292 ],
   alphaCSR[ 58 ][ 293 ],
   alphaCSR[ 58 ][ 294 ],
   alphaCSR[ 58 ][ 295 ],
   alphaCSR[ 58 ][ 296 ],
   alphaCSR[ 58 ][ 297 ],
   alphaCSR[ 58 ][ 298 ],
   alphaCSR[ 58 ][ 299 ],
   alphaCSR[ 58 ][ 300 ],
   alphaCSR[ 58 ][ 301 ],
   alphaCSR[ 58 ][ 302 ],
   alphaCSR[ 58 ][ 303 ],
   alphaCSR[ 58 ][ 304 ],
   alphaCSR[ 58 ][ 305 ],
   alphaCSR[ 58 ][ 306 ],
   alphaCSR[ 58 ][ 307 ],
   alphaCSR[ 58 ][ 308 ],
   alphaCSR[ 58 ][ 309 ],
   alphaCSR[ 58 ][ 310 ],
   alphaCSR[ 58 ][ 311 ],
   alphaCSR[ 58 ][ 312 ],
   alphaCSR[ 58 ][ 313 ],
   alphaCSR[ 58 ][ 314 ],
   alphaCSR[ 58 ][ 315 ],
   alphaCSR[ 58 ][ 316 ],
   alphaCSR[ 58 ][ 317 ],
   alphaCSR[ 58 ][ 318 ],
   alphaCSR[ 58 ][ 319 ],
   alphaCSR[ 58 ][ 320 ],
   alphaCSR[ 58 ][ 321 ],
   alphaCSR[ 58 ][ 322 ],
   alphaCSR[ 58 ][ 323 ],
   alphaCSR[ 58 ][ 324 ],
   alphaCSR[ 58 ][ 325 ],
   alphaCSR[ 58 ][ 326 ],
   alphaCSR[ 58 ][ 327 ],
   alphaCSR[ 58 ][ 328 ],
   alphaCSR[ 58 ][ 329 ],
   alphaCSR[ 58 ][ 330 ],
   alphaCSR[ 58 ][ 331 ],
   alphaCSR[ 58 ][ 332 ],
   alphaCSR[ 58 ][ 333 ],
   alphaCSR[ 58 ][ 334 ],
   alphaCSR[ 58 ][ 335 ],
   alphaCSR[ 58 ][ 336 ],
   alphaCSR[ 58 ][ 337 ],
   alphaCSR[ 58 ][ 338 ],
   alphaCSR[ 58 ][ 339 ],
   alphaCSR[ 58 ][ 340 ],
   alphaCSR[ 58 ][ 341 ],
   alphaCSR[ 58 ][ 342 ],
   alphaCSR[ 58 ][ 343 ],
   alphaCSR[ 58 ][ 344 ],
   alphaCSR[ 58 ][ 345 ],
   alphaCSR[ 58 ][ 346 ],
   alphaCSR[ 58 ][ 347 ],
   alphaCSR[ 58 ][ 348 ],
   alphaCSR[ 58 ][ 349 ],
   alphaCSR[ 58 ][ 350 ],
   alphaCSR[ 58 ][ 351 ],
   alphaCSR[ 58 ][ 352 ],
   alphaCSR[ 58 ][ 353 ],
   alphaCSR[ 58 ][ 354 ],
   alphaCSR[ 58 ][ 355 ],
   alphaCSR[ 58 ][ 356 ],
   alphaCSR[ 58 ][ 357 ],
   alphaCSR[ 58 ][ 358 ],
   alphaCSR[ 58 ][ 359 ],
   alphaCSR[ 58 ][ 360 ],
   alphaCSR[ 58 ][ 361 ],
   alphaCSR[ 58 ][ 362 ],
   alphaCSR[ 58 ][ 363 ],
   alphaCSR[ 58 ][ 364 ],
   alphaCSR[ 58 ][ 365 ],
   alphaCSR[ 58 ][ 366 ],
   alphaCSR[ 58 ][ 367 ],
   alphaCSR[ 58 ][ 368 ],
   alphaCSR[ 58 ][ 369 ],
   alphaCSR[ 58 ][ 370 ],
   alphaCSR[ 58 ][ 371 ],
   alphaCSR[ 58 ][ 372 ],
   alphaCSR[ 58 ][ 373 ],
   alphaCSR[ 58 ][ 374 ],
   alphaCSR[ 58 ][ 375 ],
   alphaCSR[ 58 ][ 376 ],
   alphaCSR[ 58 ][ 377 ],
   alphaCSR[ 58 ][ 378 ],
   alphaCSR[ 58 ][ 379 ],
   alphaCSR[ 58 ][ 380 ],
   alphaCSR[ 58 ][ 381 ],
   alphaCSR[ 58 ][ 382 ],
   alphaCSR[ 58 ][ 383 ],
   alphaCSR[ 59 ][ 0 ],
   alphaCSR[ 59 ][ 1 ],
   alphaCSR[ 59 ][ 2 ],
   alphaCSR[ 59 ][ 3 ],
   alphaCSR[ 59 ][ 4 ],
   alphaCSR[ 59 ][ 5 ],
   alphaCSR[ 59 ][ 6 ],
   alphaCSR[ 59 ][ 7 ],
   alphaCSR[ 59 ][ 8 ],
   alphaCSR[ 59 ][ 9 ],
   alphaCSR[ 59 ][ 10 ],
   alphaCSR[ 59 ][ 11 ],
   alphaCSR[ 59 ][ 12 ],
   alphaCSR[ 59 ][ 13 ],
   alphaCSR[ 59 ][ 14 ],
   alphaCSR[ 59 ][ 15 ],
   alphaCSR[ 59 ][ 16 ],
   alphaCSR[ 59 ][ 17 ],
   alphaCSR[ 59 ][ 18 ],
   alphaCSR[ 59 ][ 19 ],
   alphaCSR[ 59 ][ 20 ],
   alphaCSR[ 59 ][ 21 ],
   alphaCSR[ 59 ][ 22 ],
   alphaCSR[ 59 ][ 23 ],
   alphaCSR[ 59 ][ 24 ],
   alphaCSR[ 59 ][ 25 ],
   alphaCSR[ 59 ][ 26 ],
   alphaCSR[ 59 ][ 27 ],
   alphaCSR[ 59 ][ 28 ],
   alphaCSR[ 59 ][ 29 ],
   alphaCSR[ 59 ][ 30 ],
   alphaCSR[ 59 ][ 31 ],
   alphaCSR[ 59 ][ 32 ],
   alphaCSR[ 59 ][ 33 ],
   alphaCSR[ 59 ][ 34 ],
   alphaCSR[ 59 ][ 35 ],
   alphaCSR[ 59 ][ 36 ],
   alphaCSR[ 59 ][ 37 ],
   alphaCSR[ 59 ][ 38 ],
   alphaCSR[ 59 ][ 39 ],
   alphaCSR[ 59 ][ 40 ],
   alphaCSR[ 59 ][ 41 ],
   alphaCSR[ 59 ][ 42 ],
   alphaCSR[ 59 ][ 43 ],
   alphaCSR[ 59 ][ 44 ],
   alphaCSR[ 59 ][ 45 ],
   alphaCSR[ 59 ][ 46 ],
   alphaCSR[ 59 ][ 47 ],
   alphaCSR[ 59 ][ 48 ],
   alphaCSR[ 59 ][ 49 ],
   alphaCSR[ 59 ][ 50 ],
   alphaCSR[ 59 ][ 51 ],
   alphaCSR[ 59 ][ 52 ],
   alphaCSR[ 59 ][ 53 ],
   alphaCSR[ 59 ][ 54 ],
   alphaCSR[ 59 ][ 55 ],
   alphaCSR[ 59 ][ 56 ],
   alphaCSR[ 59 ][ 57 ],
   alphaCSR[ 59 ][ 58 ],
   alphaCSR[ 59 ][ 59 ],
   alphaCSR[ 59 ][ 60 ],
   alphaCSR[ 59 ][ 61 ],
   alphaCSR[ 59 ][ 62 ],
   alphaCSR[ 59 ][ 63 ],
   alphaCSR[ 59 ][ 64 ],
   alphaCSR[ 59 ][ 65 ],
   alphaCSR[ 59 ][ 66 ],
   alphaCSR[ 59 ][ 67 ],
   alphaCSR[ 59 ][ 68 ],
   alphaCSR[ 59 ][ 69 ],
   alphaCSR[ 59 ][ 70 ],
   alphaCSR[ 59 ][ 71 ],
   alphaCSR[ 59 ][ 72 ],
   alphaCSR[ 59 ][ 73 ],
   alphaCSR[ 59 ][ 74 ],
   alphaCSR[ 59 ][ 75 ],
   alphaCSR[ 59 ][ 76 ],
   alphaCSR[ 59 ][ 77 ],
   alphaCSR[ 59 ][ 78 ],
   alphaCSR[ 59 ][ 79 ],
   alphaCSR[ 59 ][ 80 ],
   alphaCSR[ 59 ][ 81 ],
   alphaCSR[ 59 ][ 82 ],
   alphaCSR[ 59 ][ 83 ],
   alphaCSR[ 59 ][ 84 ],
   alphaCSR[ 59 ][ 85 ],
   alphaCSR[ 59 ][ 86 ],
   alphaCSR[ 59 ][ 87 ],
   alphaCSR[ 59 ][ 88 ],
   alphaCSR[ 59 ][ 89 ],
   alphaCSR[ 59 ][ 90 ],
   alphaCSR[ 59 ][ 91 ],
   alphaCSR[ 59 ][ 92 ],
   alphaCSR[ 59 ][ 93 ],
   alphaCSR[ 59 ][ 94 ],
   alphaCSR[ 59 ][ 95 ],
   alphaCSR[ 59 ][ 96 ],
   alphaCSR[ 59 ][ 97 ],
   alphaCSR[ 59 ][ 98 ],
   alphaCSR[ 59 ][ 99 ],
   alphaCSR[ 59 ][ 100 ],
   alphaCSR[ 59 ][ 101 ],
   alphaCSR[ 59 ][ 102 ],
   alphaCSR[ 59 ][ 103 ],
   alphaCSR[ 59 ][ 104 ],
   alphaCSR[ 59 ][ 105 ],
   alphaCSR[ 59 ][ 106 ],
   alphaCSR[ 59 ][ 107 ],
   alphaCSR[ 59 ][ 108 ],
   alphaCSR[ 59 ][ 109 ],
   alphaCSR[ 59 ][ 110 ],
   alphaCSR[ 59 ][ 111 ],
   alphaCSR[ 59 ][ 112 ],
   alphaCSR[ 59 ][ 113 ],
   alphaCSR[ 59 ][ 114 ],
   alphaCSR[ 59 ][ 115 ],
   alphaCSR[ 59 ][ 116 ],
   alphaCSR[ 59 ][ 117 ],
   alphaCSR[ 59 ][ 118 ],
   alphaCSR[ 59 ][ 119 ],
   alphaCSR[ 59 ][ 120 ],
   alphaCSR[ 59 ][ 121 ],
   alphaCSR[ 59 ][ 122 ],
   alphaCSR[ 59 ][ 123 ],
   alphaCSR[ 59 ][ 124 ],
   alphaCSR[ 59 ][ 125 ],
   alphaCSR[ 59 ][ 126 ],
   alphaCSR[ 59 ][ 127 ],
   alphaCSR[ 59 ][ 128 ],
   alphaCSR[ 59 ][ 129 ],
   alphaCSR[ 59 ][ 130 ],
   alphaCSR[ 59 ][ 131 ],
   alphaCSR[ 59 ][ 132 ],
   alphaCSR[ 59 ][ 133 ],
   alphaCSR[ 59 ][ 134 ],
   alphaCSR[ 59 ][ 135 ],
   alphaCSR[ 59 ][ 136 ],
   alphaCSR[ 59 ][ 137 ],
   alphaCSR[ 59 ][ 138 ],
   alphaCSR[ 59 ][ 139 ],
   alphaCSR[ 59 ][ 140 ],
   alphaCSR[ 59 ][ 141 ],
   alphaCSR[ 59 ][ 142 ],
   alphaCSR[ 59 ][ 143 ],
   alphaCSR[ 59 ][ 144 ],
   alphaCSR[ 59 ][ 145 ],
   alphaCSR[ 59 ][ 146 ],
   alphaCSR[ 59 ][ 147 ],
   alphaCSR[ 59 ][ 148 ],
   alphaCSR[ 59 ][ 149 ],
   alphaCSR[ 59 ][ 150 ],
   alphaCSR[ 59 ][ 151 ],
   alphaCSR[ 59 ][ 152 ],
   alphaCSR[ 59 ][ 153 ],
   alphaCSR[ 59 ][ 154 ],
   alphaCSR[ 59 ][ 155 ],
   alphaCSR[ 59 ][ 156 ],
   alphaCSR[ 59 ][ 157 ],
   alphaCSR[ 59 ][ 158 ],
   alphaCSR[ 59 ][ 159 ],
   alphaCSR[ 59 ][ 160 ],
   alphaCSR[ 59 ][ 161 ],
   alphaCSR[ 59 ][ 162 ],
   alphaCSR[ 59 ][ 163 ],
   alphaCSR[ 59 ][ 164 ],
   alphaCSR[ 59 ][ 165 ],
   alphaCSR[ 59 ][ 166 ],
   alphaCSR[ 59 ][ 167 ],
   alphaCSR[ 59 ][ 168 ],
   alphaCSR[ 59 ][ 169 ],
   alphaCSR[ 59 ][ 170 ],
   alphaCSR[ 59 ][ 171 ],
   alphaCSR[ 59 ][ 172 ],
   alphaCSR[ 59 ][ 173 ],
   alphaCSR[ 59 ][ 174 ],
   alphaCSR[ 59 ][ 175 ],
   alphaCSR[ 59 ][ 176 ],
   alphaCSR[ 59 ][ 177 ],
   alphaCSR[ 59 ][ 178 ],
   alphaCSR[ 59 ][ 179 ],
   alphaCSR[ 59 ][ 180 ],
   alphaCSR[ 59 ][ 181 ],
   alphaCSR[ 59 ][ 182 ],
   alphaCSR[ 59 ][ 183 ],
   alphaCSR[ 59 ][ 184 ],
   alphaCSR[ 59 ][ 185 ],
   alphaCSR[ 59 ][ 186 ],
   alphaCSR[ 59 ][ 187 ],
   alphaCSR[ 59 ][ 188 ],
   alphaCSR[ 59 ][ 189 ],
   alphaCSR[ 59 ][ 190 ],
   alphaCSR[ 59 ][ 191 ],
   alphaCSR[ 59 ][ 192 ],
   alphaCSR[ 59 ][ 193 ],
   alphaCSR[ 59 ][ 194 ],
   alphaCSR[ 59 ][ 195 ],
   alphaCSR[ 59 ][ 196 ],
   alphaCSR[ 59 ][ 197 ],
   alphaCSR[ 59 ][ 198 ],
   alphaCSR[ 59 ][ 199 ],
   alphaCSR[ 59 ][ 200 ],
   alphaCSR[ 59 ][ 201 ],
   alphaCSR[ 59 ][ 202 ],
   alphaCSR[ 59 ][ 203 ],
   alphaCSR[ 59 ][ 204 ],
   alphaCSR[ 59 ][ 205 ],
   alphaCSR[ 59 ][ 206 ],
   alphaCSR[ 59 ][ 207 ],
   alphaCSR[ 59 ][ 208 ],
   alphaCSR[ 59 ][ 209 ],
   alphaCSR[ 59 ][ 210 ],
   alphaCSR[ 59 ][ 211 ],
   alphaCSR[ 59 ][ 212 ],
   alphaCSR[ 59 ][ 213 ],
   alphaCSR[ 59 ][ 214 ],
   alphaCSR[ 59 ][ 215 ],
   alphaCSR[ 59 ][ 216 ],
   alphaCSR[ 59 ][ 217 ],
   alphaCSR[ 59 ][ 218 ],
   alphaCSR[ 59 ][ 219 ],
   alphaCSR[ 59 ][ 220 ],
   alphaCSR[ 59 ][ 221 ],
   alphaCSR[ 59 ][ 222 ],
   alphaCSR[ 59 ][ 223 ],
   alphaCSR[ 59 ][ 224 ],
   alphaCSR[ 59 ][ 225 ],
   alphaCSR[ 59 ][ 226 ],
   alphaCSR[ 59 ][ 227 ],
   alphaCSR[ 59 ][ 228 ],
   alphaCSR[ 59 ][ 229 ],
   alphaCSR[ 59 ][ 230 ],
   alphaCSR[ 59 ][ 231 ],
   alphaCSR[ 59 ][ 232 ],
   alphaCSR[ 59 ][ 233 ],
   alphaCSR[ 59 ][ 234 ],
   alphaCSR[ 59 ][ 235 ],
   alphaCSR[ 59 ][ 236 ],
   alphaCSR[ 59 ][ 237 ],
   alphaCSR[ 59 ][ 238 ],
   alphaCSR[ 59 ][ 239 ],
   alphaCSR[ 59 ][ 240 ],
   alphaCSR[ 59 ][ 241 ],
   alphaCSR[ 59 ][ 242 ],
   alphaCSR[ 59 ][ 243 ],
   alphaCSR[ 59 ][ 244 ],
   alphaCSR[ 59 ][ 245 ],
   alphaCSR[ 59 ][ 246 ],
   alphaCSR[ 59 ][ 247 ],
   alphaCSR[ 59 ][ 248 ],
   alphaCSR[ 59 ][ 249 ],
   alphaCSR[ 59 ][ 250 ],
   alphaCSR[ 59 ][ 251 ],
   alphaCSR[ 59 ][ 252 ],
   alphaCSR[ 59 ][ 253 ],
   alphaCSR[ 59 ][ 254 ],
   alphaCSR[ 59 ][ 255 ],
   alphaCSR[ 59 ][ 256 ],
   alphaCSR[ 59 ][ 257 ],
   alphaCSR[ 59 ][ 258 ],
   alphaCSR[ 59 ][ 259 ],
   alphaCSR[ 59 ][ 260 ],
   alphaCSR[ 59 ][ 261 ],
   alphaCSR[ 59 ][ 262 ],
   alphaCSR[ 59 ][ 263 ],
   alphaCSR[ 59 ][ 264 ],
   alphaCSR[ 59 ][ 265 ],
   alphaCSR[ 59 ][ 266 ],
   alphaCSR[ 59 ][ 267 ],
   alphaCSR[ 59 ][ 268 ],
   alphaCSR[ 59 ][ 269 ],
   alphaCSR[ 59 ][ 270 ],
   alphaCSR[ 59 ][ 271 ],
   alphaCSR[ 59 ][ 272 ],
   alphaCSR[ 59 ][ 273 ],
   alphaCSR[ 59 ][ 274 ],
   alphaCSR[ 59 ][ 275 ],
   alphaCSR[ 59 ][ 276 ],
   alphaCSR[ 59 ][ 277 ],
   alphaCSR[ 59 ][ 278 ],
   alphaCSR[ 59 ][ 279 ],
   alphaCSR[ 59 ][ 280 ],
   alphaCSR[ 59 ][ 281 ],
   alphaCSR[ 59 ][ 282 ],
   alphaCSR[ 59 ][ 283 ],
   alphaCSR[ 59 ][ 284 ],
   alphaCSR[ 59 ][ 285 ],
   alphaCSR[ 59 ][ 286 ],
   alphaCSR[ 59 ][ 287 ],
   alphaCSR[ 59 ][ 288 ],
   alphaCSR[ 59 ][ 289 ],
   alphaCSR[ 59 ][ 290 ],
   alphaCSR[ 59 ][ 291 ],
   alphaCSR[ 59 ][ 292 ],
   alphaCSR[ 59 ][ 293 ],
   alphaCSR[ 59 ][ 294 ],
   alphaCSR[ 59 ][ 295 ],
   alphaCSR[ 59 ][ 296 ],
   alphaCSR[ 59 ][ 297 ],
   alphaCSR[ 59 ][ 298 ],
   alphaCSR[ 59 ][ 299 ],
   alphaCSR[ 59 ][ 300 ],
   alphaCSR[ 59 ][ 301 ],
   alphaCSR[ 59 ][ 302 ],
   alphaCSR[ 59 ][ 303 ],
   alphaCSR[ 59 ][ 304 ],
   alphaCSR[ 59 ][ 305 ],
   alphaCSR[ 59 ][ 306 ],
   alphaCSR[ 59 ][ 307 ],
   alphaCSR[ 59 ][ 308 ],
   alphaCSR[ 59 ][ 309 ],
   alphaCSR[ 59 ][ 310 ],
   alphaCSR[ 59 ][ 311 ],
   alphaCSR[ 59 ][ 312 ],
   alphaCSR[ 59 ][ 313 ],
   alphaCSR[ 59 ][ 314 ],
   alphaCSR[ 59 ][ 315 ],
   alphaCSR[ 59 ][ 316 ],
   alphaCSR[ 59 ][ 317 ],
   alphaCSR[ 59 ][ 318 ],
   alphaCSR[ 59 ][ 319 ],
   alphaCSR[ 59 ][ 320 ],
   alphaCSR[ 59 ][ 321 ],
   alphaCSR[ 59 ][ 322 ],
   alphaCSR[ 59 ][ 323 ],
   alphaCSR[ 59 ][ 324 ],
   alphaCSR[ 59 ][ 325 ],
   alphaCSR[ 59 ][ 326 ],
   alphaCSR[ 59 ][ 327 ],
   alphaCSR[ 59 ][ 328 ],
   alphaCSR[ 59 ][ 329 ],
   alphaCSR[ 59 ][ 330 ],
   alphaCSR[ 59 ][ 331 ],
   alphaCSR[ 59 ][ 332 ],
   alphaCSR[ 59 ][ 333 ],
   alphaCSR[ 59 ][ 334 ],
   alphaCSR[ 59 ][ 335 ],
   alphaCSR[ 59 ][ 336 ],
   alphaCSR[ 59 ][ 337 ],
   alphaCSR[ 59 ][ 338 ],
   alphaCSR[ 59 ][ 339 ],
   alphaCSR[ 59 ][ 340 ],
   alphaCSR[ 59 ][ 341 ],
   alphaCSR[ 59 ][ 342 ],
   alphaCSR[ 59 ][ 343 ],
   alphaCSR[ 59 ][ 344 ],
   alphaCSR[ 59 ][ 345 ],
   alphaCSR[ 59 ][ 346 ],
   alphaCSR[ 59 ][ 347 ],
   alphaCSR[ 59 ][ 348 ],
   alphaCSR[ 59 ][ 349 ],
   alphaCSR[ 59 ][ 350 ],
   alphaCSR[ 59 ][ 351 ],
   alphaCSR[ 59 ][ 352 ],
   alphaCSR[ 59 ][ 353 ],
   alphaCSR[ 59 ][ 354 ],
   alphaCSR[ 59 ][ 355 ],
   alphaCSR[ 59 ][ 356 ],
   alphaCSR[ 59 ][ 357 ],
   alphaCSR[ 59 ][ 358 ],
   alphaCSR[ 59 ][ 359 ],
   alphaCSR[ 59 ][ 360 ],
   alphaCSR[ 59 ][ 361 ],
   alphaCSR[ 59 ][ 362 ],
   alphaCSR[ 59 ][ 363 ],
   alphaCSR[ 59 ][ 364 ],
   alphaCSR[ 59 ][ 365 ],
   alphaCSR[ 59 ][ 366 ],
   alphaCSR[ 59 ][ 367 ],
   alphaCSR[ 59 ][ 368 ],
   alphaCSR[ 59 ][ 369 ],
   alphaCSR[ 59 ][ 370 ],
   alphaCSR[ 59 ][ 371 ],
   alphaCSR[ 59 ][ 372 ],
   alphaCSR[ 59 ][ 373 ],
   alphaCSR[ 59 ][ 374 ],
   alphaCSR[ 59 ][ 375 ],
   alphaCSR[ 59 ][ 376 ],
   alphaCSR[ 59 ][ 377 ],
   alphaCSR[ 59 ][ 378 ],
   alphaCSR[ 59 ][ 379 ],
   alphaCSR[ 59 ][ 380 ],
   alphaCSR[ 59 ][ 381 ],
   alphaCSR[ 59 ][ 382 ],
   alphaCSR[ 59 ][ 383 ],
   alphaCSR[ 60 ][ 0 ],
   alphaCSR[ 60 ][ 1 ],
   alphaCSR[ 60 ][ 2 ],
   alphaCSR[ 60 ][ 3 ],
   alphaCSR[ 60 ][ 4 ],
   alphaCSR[ 60 ][ 5 ],
   alphaCSR[ 60 ][ 6 ],
   alphaCSR[ 60 ][ 7 ],
   alphaCSR[ 60 ][ 8 ],
   alphaCSR[ 60 ][ 9 ],
   alphaCSR[ 60 ][ 10 ],
   alphaCSR[ 60 ][ 11 ],
   alphaCSR[ 60 ][ 12 ],
   alphaCSR[ 60 ][ 13 ],
   alphaCSR[ 60 ][ 14 ],
   alphaCSR[ 60 ][ 15 ],
   alphaCSR[ 60 ][ 16 ],
   alphaCSR[ 60 ][ 17 ],
   alphaCSR[ 60 ][ 18 ],
   alphaCSR[ 60 ][ 19 ],
   alphaCSR[ 60 ][ 20 ],
   alphaCSR[ 60 ][ 21 ],
   alphaCSR[ 60 ][ 22 ],
   alphaCSR[ 60 ][ 23 ],
   alphaCSR[ 60 ][ 24 ],
   alphaCSR[ 60 ][ 25 ],
   alphaCSR[ 60 ][ 26 ],
   alphaCSR[ 60 ][ 27 ],
   alphaCSR[ 60 ][ 28 ],
   alphaCSR[ 60 ][ 29 ],
   alphaCSR[ 60 ][ 30 ],
   alphaCSR[ 60 ][ 31 ],
   alphaCSR[ 60 ][ 32 ],
   alphaCSR[ 60 ][ 33 ],
   alphaCSR[ 60 ][ 34 ],
   alphaCSR[ 60 ][ 35 ],
   alphaCSR[ 60 ][ 36 ],
   alphaCSR[ 60 ][ 37 ],
   alphaCSR[ 60 ][ 38 ],
   alphaCSR[ 60 ][ 39 ],
   alphaCSR[ 60 ][ 40 ],
   alphaCSR[ 60 ][ 41 ],
   alphaCSR[ 60 ][ 42 ],
   alphaCSR[ 60 ][ 43 ],
   alphaCSR[ 60 ][ 44 ],
   alphaCSR[ 60 ][ 45 ],
   alphaCSR[ 60 ][ 46 ],
   alphaCSR[ 60 ][ 47 ],
   alphaCSR[ 60 ][ 48 ],
   alphaCSR[ 60 ][ 49 ],
   alphaCSR[ 60 ][ 50 ],
   alphaCSR[ 60 ][ 51 ],
   alphaCSR[ 60 ][ 52 ],
   alphaCSR[ 60 ][ 53 ],
   alphaCSR[ 60 ][ 54 ],
   alphaCSR[ 60 ][ 55 ],
   alphaCSR[ 60 ][ 56 ],
   alphaCSR[ 60 ][ 57 ],
   alphaCSR[ 60 ][ 58 ],
   alphaCSR[ 60 ][ 59 ],
   alphaCSR[ 60 ][ 60 ],
   alphaCSR[ 60 ][ 61 ],
   alphaCSR[ 60 ][ 62 ],
   alphaCSR[ 60 ][ 63 ],
   alphaCSR[ 60 ][ 64 ],
   alphaCSR[ 60 ][ 65 ],
   alphaCSR[ 60 ][ 66 ],
   alphaCSR[ 60 ][ 67 ],
   alphaCSR[ 60 ][ 68 ],
   alphaCSR[ 60 ][ 69 ],
   alphaCSR[ 60 ][ 70 ],
   alphaCSR[ 60 ][ 71 ],
   alphaCSR[ 60 ][ 72 ],
   alphaCSR[ 60 ][ 73 ],
   alphaCSR[ 60 ][ 74 ],
   alphaCSR[ 60 ][ 75 ],
   alphaCSR[ 60 ][ 76 ],
   alphaCSR[ 60 ][ 77 ],
   alphaCSR[ 60 ][ 78 ],
   alphaCSR[ 60 ][ 79 ],
   alphaCSR[ 60 ][ 80 ],
   alphaCSR[ 60 ][ 81 ],
   alphaCSR[ 60 ][ 82 ],
   alphaCSR[ 60 ][ 83 ],
   alphaCSR[ 60 ][ 84 ],
   alphaCSR[ 60 ][ 85 ],
   alphaCSR[ 60 ][ 86 ],
   alphaCSR[ 60 ][ 87 ],
   alphaCSR[ 60 ][ 88 ],
   alphaCSR[ 60 ][ 89 ],
   alphaCSR[ 60 ][ 90 ],
   alphaCSR[ 60 ][ 91 ],
   alphaCSR[ 60 ][ 92 ],
   alphaCSR[ 60 ][ 93 ],
   alphaCSR[ 60 ][ 94 ],
   alphaCSR[ 60 ][ 95 ],
   alphaCSR[ 60 ][ 96 ],
   alphaCSR[ 60 ][ 97 ],
   alphaCSR[ 60 ][ 98 ],
   alphaCSR[ 60 ][ 99 ],
   alphaCSR[ 60 ][ 100 ],
   alphaCSR[ 60 ][ 101 ],
   alphaCSR[ 60 ][ 102 ],
   alphaCSR[ 60 ][ 103 ],
   alphaCSR[ 60 ][ 104 ],
   alphaCSR[ 60 ][ 105 ],
   alphaCSR[ 60 ][ 106 ],
   alphaCSR[ 60 ][ 107 ],
   alphaCSR[ 60 ][ 108 ],
   alphaCSR[ 60 ][ 109 ],
   alphaCSR[ 60 ][ 110 ],
   alphaCSR[ 60 ][ 111 ],
   alphaCSR[ 60 ][ 112 ],
   alphaCSR[ 60 ][ 113 ],
   alphaCSR[ 60 ][ 114 ],
   alphaCSR[ 60 ][ 115 ],
   alphaCSR[ 60 ][ 116 ],
   alphaCSR[ 60 ][ 117 ],
   alphaCSR[ 60 ][ 118 ],
   alphaCSR[ 60 ][ 119 ],
   alphaCSR[ 60 ][ 120 ],
   alphaCSR[ 60 ][ 121 ],
   alphaCSR[ 60 ][ 122 ],
   alphaCSR[ 60 ][ 123 ],
   alphaCSR[ 60 ][ 124 ],
   alphaCSR[ 60 ][ 125 ],
   alphaCSR[ 60 ][ 126 ],
   alphaCSR[ 60 ][ 127 ],
   alphaCSR[ 60 ][ 128 ],
   alphaCSR[ 60 ][ 129 ],
   alphaCSR[ 60 ][ 130 ],
   alphaCSR[ 60 ][ 131 ],
   alphaCSR[ 60 ][ 132 ],
   alphaCSR[ 60 ][ 133 ],
   alphaCSR[ 60 ][ 134 ],
   alphaCSR[ 60 ][ 135 ],
   alphaCSR[ 60 ][ 136 ],
   alphaCSR[ 60 ][ 137 ],
   alphaCSR[ 60 ][ 138 ],
   alphaCSR[ 60 ][ 139 ],
   alphaCSR[ 60 ][ 140 ],
   alphaCSR[ 60 ][ 141 ],
   alphaCSR[ 60 ][ 142 ],
   alphaCSR[ 60 ][ 143 ],
   alphaCSR[ 60 ][ 144 ],
   alphaCSR[ 60 ][ 145 ],
   alphaCSR[ 60 ][ 146 ],
   alphaCSR[ 60 ][ 147 ],
   alphaCSR[ 60 ][ 148 ],
   alphaCSR[ 60 ][ 149 ],
   alphaCSR[ 60 ][ 150 ],
   alphaCSR[ 60 ][ 151 ],
   alphaCSR[ 60 ][ 152 ],
   alphaCSR[ 60 ][ 153 ],
   alphaCSR[ 60 ][ 154 ],
   alphaCSR[ 60 ][ 155 ],
   alphaCSR[ 60 ][ 156 ],
   alphaCSR[ 60 ][ 157 ],
   alphaCSR[ 60 ][ 158 ],
   alphaCSR[ 60 ][ 159 ],
   alphaCSR[ 60 ][ 160 ],
   alphaCSR[ 60 ][ 161 ],
   alphaCSR[ 60 ][ 162 ],
   alphaCSR[ 60 ][ 163 ],
   alphaCSR[ 60 ][ 164 ],
   alphaCSR[ 60 ][ 165 ],
   alphaCSR[ 60 ][ 166 ],
   alphaCSR[ 60 ][ 167 ],
   alphaCSR[ 60 ][ 168 ],
   alphaCSR[ 60 ][ 169 ],
   alphaCSR[ 60 ][ 170 ],
   alphaCSR[ 60 ][ 171 ],
   alphaCSR[ 60 ][ 172 ],
   alphaCSR[ 60 ][ 173 ],
   alphaCSR[ 60 ][ 174 ],
   alphaCSR[ 60 ][ 175 ],
   alphaCSR[ 60 ][ 176 ],
   alphaCSR[ 60 ][ 177 ],
   alphaCSR[ 60 ][ 178 ],
   alphaCSR[ 60 ][ 179 ],
   alphaCSR[ 60 ][ 180 ],
   alphaCSR[ 60 ][ 181 ],
   alphaCSR[ 60 ][ 182 ],
   alphaCSR[ 60 ][ 183 ],
   alphaCSR[ 60 ][ 184 ],
   alphaCSR[ 60 ][ 185 ],
   alphaCSR[ 60 ][ 186 ],
   alphaCSR[ 60 ][ 187 ],
   alphaCSR[ 60 ][ 188 ],
   alphaCSR[ 60 ][ 189 ],
   alphaCSR[ 60 ][ 190 ],
   alphaCSR[ 60 ][ 191 ],
   alphaCSR[ 60 ][ 192 ],
   alphaCSR[ 60 ][ 193 ],
   alphaCSR[ 60 ][ 194 ],
   alphaCSR[ 60 ][ 195 ],
   alphaCSR[ 60 ][ 196 ],
   alphaCSR[ 60 ][ 197 ],
   alphaCSR[ 60 ][ 198 ],
   alphaCSR[ 60 ][ 199 ],
   alphaCSR[ 60 ][ 200 ],
   alphaCSR[ 60 ][ 201 ],
   alphaCSR[ 60 ][ 202 ],
   alphaCSR[ 60 ][ 203 ],
   alphaCSR[ 60 ][ 204 ],
   alphaCSR[ 60 ][ 205 ],
   alphaCSR[ 60 ][ 206 ],
   alphaCSR[ 60 ][ 207 ],
   alphaCSR[ 60 ][ 208 ],
   alphaCSR[ 60 ][ 209 ],
   alphaCSR[ 60 ][ 210 ],
   alphaCSR[ 60 ][ 211 ],
   alphaCSR[ 60 ][ 212 ],
   alphaCSR[ 60 ][ 213 ],
   alphaCSR[ 60 ][ 214 ],
   alphaCSR[ 60 ][ 215 ],
   alphaCSR[ 60 ][ 216 ],
   alphaCSR[ 60 ][ 217 ],
   alphaCSR[ 60 ][ 218 ],
   alphaCSR[ 60 ][ 219 ],
   alphaCSR[ 60 ][ 220 ],
   alphaCSR[ 60 ][ 221 ],
   alphaCSR[ 60 ][ 222 ],
   alphaCSR[ 60 ][ 223 ],
   alphaCSR[ 60 ][ 224 ],
   alphaCSR[ 60 ][ 225 ],
   alphaCSR[ 60 ][ 226 ],
   alphaCSR[ 60 ][ 227 ],
   alphaCSR[ 60 ][ 228 ],
   alphaCSR[ 60 ][ 229 ],
   alphaCSR[ 60 ][ 230 ],
   alphaCSR[ 60 ][ 231 ],
   alphaCSR[ 60 ][ 232 ],
   alphaCSR[ 60 ][ 233 ],
   alphaCSR[ 60 ][ 234 ],
   alphaCSR[ 60 ][ 235 ],
   alphaCSR[ 60 ][ 236 ],
   alphaCSR[ 60 ][ 237 ],
   alphaCSR[ 60 ][ 238 ],
   alphaCSR[ 60 ][ 239 ],
   alphaCSR[ 60 ][ 240 ],
   alphaCSR[ 60 ][ 241 ],
   alphaCSR[ 60 ][ 242 ],
   alphaCSR[ 60 ][ 243 ],
   alphaCSR[ 60 ][ 244 ],
   alphaCSR[ 60 ][ 245 ],
   alphaCSR[ 60 ][ 246 ],
   alphaCSR[ 60 ][ 247 ],
   alphaCSR[ 60 ][ 248 ],
   alphaCSR[ 60 ][ 249 ],
   alphaCSR[ 60 ][ 250 ],
   alphaCSR[ 60 ][ 251 ],
   alphaCSR[ 60 ][ 252 ],
   alphaCSR[ 60 ][ 253 ],
   alphaCSR[ 60 ][ 254 ],
   alphaCSR[ 60 ][ 255 ],
   alphaCSR[ 60 ][ 256 ],
   alphaCSR[ 60 ][ 257 ],
   alphaCSR[ 60 ][ 258 ],
   alphaCSR[ 60 ][ 259 ],
   alphaCSR[ 60 ][ 260 ],
   alphaCSR[ 60 ][ 261 ],
   alphaCSR[ 60 ][ 262 ],
   alphaCSR[ 60 ][ 263 ],
   alphaCSR[ 60 ][ 264 ],
   alphaCSR[ 60 ][ 265 ],
   alphaCSR[ 60 ][ 266 ],
   alphaCSR[ 60 ][ 267 ],
   alphaCSR[ 60 ][ 268 ],
   alphaCSR[ 60 ][ 269 ],
   alphaCSR[ 60 ][ 270 ],
   alphaCSR[ 60 ][ 271 ],
   alphaCSR[ 60 ][ 272 ],
   alphaCSR[ 60 ][ 273 ],
   alphaCSR[ 60 ][ 274 ],
   alphaCSR[ 60 ][ 275 ],
   alphaCSR[ 60 ][ 276 ],
   alphaCSR[ 60 ][ 277 ],
   alphaCSR[ 60 ][ 278 ],
   alphaCSR[ 60 ][ 279 ],
   alphaCSR[ 60 ][ 280 ],
   alphaCSR[ 60 ][ 281 ],
   alphaCSR[ 60 ][ 282 ],
   alphaCSR[ 60 ][ 283 ],
   alphaCSR[ 60 ][ 284 ],
   alphaCSR[ 60 ][ 285 ],
   alphaCSR[ 60 ][ 286 ],
   alphaCSR[ 60 ][ 287 ],
   alphaCSR[ 60 ][ 288 ],
   alphaCSR[ 60 ][ 289 ],
   alphaCSR[ 60 ][ 290 ],
   alphaCSR[ 60 ][ 291 ],
   alphaCSR[ 60 ][ 292 ],
   alphaCSR[ 60 ][ 293 ],
   alphaCSR[ 60 ][ 294 ],
   alphaCSR[ 60 ][ 295 ],
   alphaCSR[ 60 ][ 296 ],
   alphaCSR[ 60 ][ 297 ],
   alphaCSR[ 60 ][ 298 ],
   alphaCSR[ 60 ][ 299 ],
   alphaCSR[ 60 ][ 300 ],
   alphaCSR[ 60 ][ 301 ],
   alphaCSR[ 60 ][ 302 ],
   alphaCSR[ 60 ][ 303 ],
   alphaCSR[ 60 ][ 304 ],
   alphaCSR[ 60 ][ 305 ],
   alphaCSR[ 60 ][ 306 ],
   alphaCSR[ 60 ][ 307 ],
   alphaCSR[ 60 ][ 308 ],
   alphaCSR[ 60 ][ 309 ],
   alphaCSR[ 60 ][ 310 ],
   alphaCSR[ 60 ][ 311 ],
   alphaCSR[ 60 ][ 312 ],
   alphaCSR[ 60 ][ 313 ],
   alphaCSR[ 60 ][ 314 ],
   alphaCSR[ 60 ][ 315 ],
   alphaCSR[ 60 ][ 316 ],
   alphaCSR[ 60 ][ 317 ],
   alphaCSR[ 60 ][ 318 ],
   alphaCSR[ 60 ][ 319 ],
   alphaCSR[ 60 ][ 320 ],
   alphaCSR[ 60 ][ 321 ],
   alphaCSR[ 60 ][ 322 ],
   alphaCSR[ 60 ][ 323 ],
   alphaCSR[ 60 ][ 324 ],
   alphaCSR[ 60 ][ 325 ],
   alphaCSR[ 60 ][ 326 ],
   alphaCSR[ 60 ][ 327 ],
   alphaCSR[ 60 ][ 328 ],
   alphaCSR[ 60 ][ 329 ],
   alphaCSR[ 60 ][ 330 ],
   alphaCSR[ 60 ][ 331 ],
   alphaCSR[ 60 ][ 332 ],
   alphaCSR[ 60 ][ 333 ],
   alphaCSR[ 60 ][ 334 ],
   alphaCSR[ 60 ][ 335 ],
   alphaCSR[ 60 ][ 336 ],
   alphaCSR[ 60 ][ 337 ],
   alphaCSR[ 60 ][ 338 ],
   alphaCSR[ 60 ][ 339 ],
   alphaCSR[ 60 ][ 340 ],
   alphaCSR[ 60 ][ 341 ],
   alphaCSR[ 60 ][ 342 ],
   alphaCSR[ 60 ][ 343 ],
   alphaCSR[ 60 ][ 344 ],
   alphaCSR[ 60 ][ 345 ],
   alphaCSR[ 60 ][ 346 ],
   alphaCSR[ 60 ][ 347 ],
   alphaCSR[ 60 ][ 348 ],
   alphaCSR[ 60 ][ 349 ],
   alphaCSR[ 60 ][ 350 ],
   alphaCSR[ 60 ][ 351 ],
   alphaCSR[ 60 ][ 352 ],
   alphaCSR[ 60 ][ 353 ],
   alphaCSR[ 60 ][ 354 ],
   alphaCSR[ 60 ][ 355 ],
   alphaCSR[ 60 ][ 356 ],
   alphaCSR[ 60 ][ 357 ],
   alphaCSR[ 60 ][ 358 ],
   alphaCSR[ 60 ][ 359 ],
   alphaCSR[ 60 ][ 360 ],
   alphaCSR[ 60 ][ 361 ],
   alphaCSR[ 60 ][ 362 ],
   alphaCSR[ 60 ][ 363 ],
   alphaCSR[ 60 ][ 364 ],
   alphaCSR[ 60 ][ 365 ],
   alphaCSR[ 60 ][ 366 ],
   alphaCSR[ 60 ][ 367 ],
   alphaCSR[ 60 ][ 368 ],
   alphaCSR[ 60 ][ 369 ],
   alphaCSR[ 60 ][ 370 ],
   alphaCSR[ 60 ][ 371 ],
   alphaCSR[ 60 ][ 372 ],
   alphaCSR[ 60 ][ 373 ],
   alphaCSR[ 60 ][ 374 ],
   alphaCSR[ 60 ][ 375 ],
   alphaCSR[ 60 ][ 376 ],
   alphaCSR[ 60 ][ 377 ],
   alphaCSR[ 60 ][ 378 ],
   alphaCSR[ 60 ][ 379 ],
   alphaCSR[ 60 ][ 380 ],
   alphaCSR[ 60 ][ 381 ],
   alphaCSR[ 60 ][ 382 ],
   alphaCSR[ 60 ][ 383 ],
   alphaCSR[ 61 ][ 0 ],
   alphaCSR[ 61 ][ 1 ],
   alphaCSR[ 61 ][ 2 ],
   alphaCSR[ 61 ][ 3 ],
   alphaCSR[ 61 ][ 4 ],
   alphaCSR[ 61 ][ 5 ],
   alphaCSR[ 61 ][ 6 ],
   alphaCSR[ 61 ][ 7 ],
   alphaCSR[ 61 ][ 8 ],
   alphaCSR[ 61 ][ 9 ],
   alphaCSR[ 61 ][ 10 ],
   alphaCSR[ 61 ][ 11 ],
   alphaCSR[ 61 ][ 12 ],
   alphaCSR[ 61 ][ 13 ],
   alphaCSR[ 61 ][ 14 ],
   alphaCSR[ 61 ][ 15 ],
   alphaCSR[ 61 ][ 16 ],
   alphaCSR[ 61 ][ 17 ],
   alphaCSR[ 61 ][ 18 ],
   alphaCSR[ 61 ][ 19 ],
   alphaCSR[ 61 ][ 20 ],
   alphaCSR[ 61 ][ 21 ],
   alphaCSR[ 61 ][ 22 ],
   alphaCSR[ 61 ][ 23 ],
   alphaCSR[ 61 ][ 24 ],
   alphaCSR[ 61 ][ 25 ],
   alphaCSR[ 61 ][ 26 ],
   alphaCSR[ 61 ][ 27 ],
   alphaCSR[ 61 ][ 28 ],
   alphaCSR[ 61 ][ 29 ],
   alphaCSR[ 61 ][ 30 ],
   alphaCSR[ 61 ][ 31 ],
   alphaCSR[ 61 ][ 32 ],
   alphaCSR[ 61 ][ 33 ],
   alphaCSR[ 61 ][ 34 ],
   alphaCSR[ 61 ][ 35 ],
   alphaCSR[ 61 ][ 36 ],
   alphaCSR[ 61 ][ 37 ],
   alphaCSR[ 61 ][ 38 ],
   alphaCSR[ 61 ][ 39 ],
   alphaCSR[ 61 ][ 40 ],
   alphaCSR[ 61 ][ 41 ],
   alphaCSR[ 61 ][ 42 ],
   alphaCSR[ 61 ][ 43 ],
   alphaCSR[ 61 ][ 44 ],
   alphaCSR[ 61 ][ 45 ],
   alphaCSR[ 61 ][ 46 ],
   alphaCSR[ 61 ][ 47 ],
   alphaCSR[ 61 ][ 48 ],
   alphaCSR[ 61 ][ 49 ],
   alphaCSR[ 61 ][ 50 ],
   alphaCSR[ 61 ][ 51 ],
   alphaCSR[ 61 ][ 52 ],
   alphaCSR[ 61 ][ 53 ],
   alphaCSR[ 61 ][ 54 ],
   alphaCSR[ 61 ][ 55 ],
   alphaCSR[ 61 ][ 56 ],
   alphaCSR[ 61 ][ 57 ],
   alphaCSR[ 61 ][ 58 ],
   alphaCSR[ 61 ][ 59 ],
   alphaCSR[ 61 ][ 60 ],
   alphaCSR[ 61 ][ 61 ],
   alphaCSR[ 61 ][ 62 ],
   alphaCSR[ 61 ][ 63 ],
   alphaCSR[ 61 ][ 64 ],
   alphaCSR[ 61 ][ 65 ],
   alphaCSR[ 61 ][ 66 ],
   alphaCSR[ 61 ][ 67 ],
   alphaCSR[ 61 ][ 68 ],
   alphaCSR[ 61 ][ 69 ],
   alphaCSR[ 61 ][ 70 ],
   alphaCSR[ 61 ][ 71 ],
   alphaCSR[ 61 ][ 72 ],
   alphaCSR[ 61 ][ 73 ],
   alphaCSR[ 61 ][ 74 ],
   alphaCSR[ 61 ][ 75 ],
   alphaCSR[ 61 ][ 76 ],
   alphaCSR[ 61 ][ 77 ],
   alphaCSR[ 61 ][ 78 ],
   alphaCSR[ 61 ][ 79 ],
   alphaCSR[ 61 ][ 80 ],
   alphaCSR[ 61 ][ 81 ],
   alphaCSR[ 61 ][ 82 ],
   alphaCSR[ 61 ][ 83 ],
   alphaCSR[ 61 ][ 84 ],
   alphaCSR[ 61 ][ 85 ],
   alphaCSR[ 61 ][ 86 ],
   alphaCSR[ 61 ][ 87 ],
   alphaCSR[ 61 ][ 88 ],
   alphaCSR[ 61 ][ 89 ],
   alphaCSR[ 61 ][ 90 ],
   alphaCSR[ 61 ][ 91 ],
   alphaCSR[ 61 ][ 92 ],
   alphaCSR[ 61 ][ 93 ],
   alphaCSR[ 61 ][ 94 ],
   alphaCSR[ 61 ][ 95 ],
   alphaCSR[ 61 ][ 96 ],
   alphaCSR[ 61 ][ 97 ],
   alphaCSR[ 61 ][ 98 ],
   alphaCSR[ 61 ][ 99 ],
   alphaCSR[ 61 ][ 100 ],
   alphaCSR[ 61 ][ 101 ],
   alphaCSR[ 61 ][ 102 ],
   alphaCSR[ 61 ][ 103 ],
   alphaCSR[ 61 ][ 104 ],
   alphaCSR[ 61 ][ 105 ],
   alphaCSR[ 61 ][ 106 ],
   alphaCSR[ 61 ][ 107 ],
   alphaCSR[ 61 ][ 108 ],
   alphaCSR[ 61 ][ 109 ],
   alphaCSR[ 61 ][ 110 ],
   alphaCSR[ 61 ][ 111 ],
   alphaCSR[ 61 ][ 112 ],
   alphaCSR[ 61 ][ 113 ],
   alphaCSR[ 61 ][ 114 ],
   alphaCSR[ 61 ][ 115 ],
   alphaCSR[ 61 ][ 116 ],
   alphaCSR[ 61 ][ 117 ],
   alphaCSR[ 61 ][ 118 ],
   alphaCSR[ 61 ][ 119 ],
   alphaCSR[ 61 ][ 120 ],
   alphaCSR[ 61 ][ 121 ],
   alphaCSR[ 61 ][ 122 ],
   alphaCSR[ 61 ][ 123 ],
   alphaCSR[ 61 ][ 124 ],
   alphaCSR[ 61 ][ 125 ],
   alphaCSR[ 61 ][ 126 ],
   alphaCSR[ 61 ][ 127 ],
   alphaCSR[ 61 ][ 128 ],
   alphaCSR[ 61 ][ 129 ],
   alphaCSR[ 61 ][ 130 ],
   alphaCSR[ 61 ][ 131 ],
   alphaCSR[ 61 ][ 132 ],
   alphaCSR[ 61 ][ 133 ],
   alphaCSR[ 61 ][ 134 ],
   alphaCSR[ 61 ][ 135 ],
   alphaCSR[ 61 ][ 136 ],
   alphaCSR[ 61 ][ 137 ],
   alphaCSR[ 61 ][ 138 ],
   alphaCSR[ 61 ][ 139 ],
   alphaCSR[ 61 ][ 140 ],
   alphaCSR[ 61 ][ 141 ],
   alphaCSR[ 61 ][ 142 ],
   alphaCSR[ 61 ][ 143 ],
   alphaCSR[ 61 ][ 144 ],
   alphaCSR[ 61 ][ 145 ],
   alphaCSR[ 61 ][ 146 ],
   alphaCSR[ 61 ][ 147 ],
   alphaCSR[ 61 ][ 148 ],
   alphaCSR[ 61 ][ 149 ],
   alphaCSR[ 61 ][ 150 ],
   alphaCSR[ 61 ][ 151 ],
   alphaCSR[ 61 ][ 152 ],
   alphaCSR[ 61 ][ 153 ],
   alphaCSR[ 61 ][ 154 ],
   alphaCSR[ 61 ][ 155 ],
   alphaCSR[ 61 ][ 156 ],
   alphaCSR[ 61 ][ 157 ],
   alphaCSR[ 61 ][ 158 ],
   alphaCSR[ 61 ][ 159 ],
   alphaCSR[ 61 ][ 160 ],
   alphaCSR[ 61 ][ 161 ],
   alphaCSR[ 61 ][ 162 ],
   alphaCSR[ 61 ][ 163 ],
   alphaCSR[ 61 ][ 164 ],
   alphaCSR[ 61 ][ 165 ],
   alphaCSR[ 61 ][ 166 ],
   alphaCSR[ 61 ][ 167 ],
   alphaCSR[ 61 ][ 168 ],
   alphaCSR[ 61 ][ 169 ],
   alphaCSR[ 61 ][ 170 ],
   alphaCSR[ 61 ][ 171 ],
   alphaCSR[ 61 ][ 172 ],
   alphaCSR[ 61 ][ 173 ],
   alphaCSR[ 61 ][ 174 ],
   alphaCSR[ 61 ][ 175 ],
   alphaCSR[ 61 ][ 176 ],
   alphaCSR[ 61 ][ 177 ],
   alphaCSR[ 61 ][ 178 ],
   alphaCSR[ 61 ][ 179 ],
   alphaCSR[ 61 ][ 180 ],
   alphaCSR[ 61 ][ 181 ],
   alphaCSR[ 61 ][ 182 ],
   alphaCSR[ 61 ][ 183 ],
   alphaCSR[ 61 ][ 184 ],
   alphaCSR[ 61 ][ 185 ],
   alphaCSR[ 61 ][ 186 ],
   alphaCSR[ 61 ][ 187 ],
   alphaCSR[ 61 ][ 188 ],
   alphaCSR[ 61 ][ 189 ],
   alphaCSR[ 61 ][ 190 ],
   alphaCSR[ 61 ][ 191 ],
   alphaCSR[ 61 ][ 192 ],
   alphaCSR[ 61 ][ 193 ],
   alphaCSR[ 61 ][ 194 ],
   alphaCSR[ 61 ][ 195 ],
   alphaCSR[ 61 ][ 196 ],
   alphaCSR[ 61 ][ 197 ],
   alphaCSR[ 61 ][ 198 ],
   alphaCSR[ 61 ][ 199 ],
   alphaCSR[ 61 ][ 200 ],
   alphaCSR[ 61 ][ 201 ],
   alphaCSR[ 61 ][ 202 ],
   alphaCSR[ 61 ][ 203 ],
   alphaCSR[ 61 ][ 204 ],
   alphaCSR[ 61 ][ 205 ],
   alphaCSR[ 61 ][ 206 ],
   alphaCSR[ 61 ][ 207 ],
   alphaCSR[ 61 ][ 208 ],
   alphaCSR[ 61 ][ 209 ],
   alphaCSR[ 61 ][ 210 ],
   alphaCSR[ 61 ][ 211 ],
   alphaCSR[ 61 ][ 212 ],
   alphaCSR[ 61 ][ 213 ],
   alphaCSR[ 61 ][ 214 ],
   alphaCSR[ 61 ][ 215 ],
   alphaCSR[ 61 ][ 216 ],
   alphaCSR[ 61 ][ 217 ],
   alphaCSR[ 61 ][ 218 ],
   alphaCSR[ 61 ][ 219 ],
   alphaCSR[ 61 ][ 220 ],
   alphaCSR[ 61 ][ 221 ],
   alphaCSR[ 61 ][ 222 ],
   alphaCSR[ 61 ][ 223 ],
   alphaCSR[ 61 ][ 224 ],
   alphaCSR[ 61 ][ 225 ],
   alphaCSR[ 61 ][ 226 ],
   alphaCSR[ 61 ][ 227 ],
   alphaCSR[ 61 ][ 228 ],
   alphaCSR[ 61 ][ 229 ],
   alphaCSR[ 61 ][ 230 ],
   alphaCSR[ 61 ][ 231 ],
   alphaCSR[ 61 ][ 232 ],
   alphaCSR[ 61 ][ 233 ],
   alphaCSR[ 61 ][ 234 ],
   alphaCSR[ 61 ][ 235 ],
   alphaCSR[ 61 ][ 236 ],
   alphaCSR[ 61 ][ 237 ],
   alphaCSR[ 61 ][ 238 ],
   alphaCSR[ 61 ][ 239 ],
   alphaCSR[ 61 ][ 240 ],
   alphaCSR[ 61 ][ 241 ],
   alphaCSR[ 61 ][ 242 ],
   alphaCSR[ 61 ][ 243 ],
   alphaCSR[ 61 ][ 244 ],
   alphaCSR[ 61 ][ 245 ],
   alphaCSR[ 61 ][ 246 ],
   alphaCSR[ 61 ][ 247 ],
   alphaCSR[ 61 ][ 248 ],
   alphaCSR[ 61 ][ 249 ],
   alphaCSR[ 61 ][ 250 ],
   alphaCSR[ 61 ][ 251 ],
   alphaCSR[ 61 ][ 252 ],
   alphaCSR[ 61 ][ 253 ],
   alphaCSR[ 61 ][ 254 ],
   alphaCSR[ 61 ][ 255 ],
   alphaCSR[ 61 ][ 256 ],
   alphaCSR[ 61 ][ 257 ],
   alphaCSR[ 61 ][ 258 ],
   alphaCSR[ 61 ][ 259 ],
   alphaCSR[ 61 ][ 260 ],
   alphaCSR[ 61 ][ 261 ],
   alphaCSR[ 61 ][ 262 ],
   alphaCSR[ 61 ][ 263 ],
   alphaCSR[ 61 ][ 264 ],
   alphaCSR[ 61 ][ 265 ],
   alphaCSR[ 61 ][ 266 ],
   alphaCSR[ 61 ][ 267 ],
   alphaCSR[ 61 ][ 268 ],
   alphaCSR[ 61 ][ 269 ],
   alphaCSR[ 61 ][ 270 ],
   alphaCSR[ 61 ][ 271 ],
   alphaCSR[ 61 ][ 272 ],
   alphaCSR[ 61 ][ 273 ],
   alphaCSR[ 61 ][ 274 ],
   alphaCSR[ 61 ][ 275 ],
   alphaCSR[ 61 ][ 276 ],
   alphaCSR[ 61 ][ 277 ],
   alphaCSR[ 61 ][ 278 ],
   alphaCSR[ 61 ][ 279 ],
   alphaCSR[ 61 ][ 280 ],
   alphaCSR[ 61 ][ 281 ],
   alphaCSR[ 61 ][ 282 ],
   alphaCSR[ 61 ][ 283 ],
   alphaCSR[ 61 ][ 284 ],
   alphaCSR[ 61 ][ 285 ],
   alphaCSR[ 61 ][ 286 ],
   alphaCSR[ 61 ][ 287 ],
   alphaCSR[ 61 ][ 288 ],
   alphaCSR[ 61 ][ 289 ],
   alphaCSR[ 61 ][ 290 ],
   alphaCSR[ 61 ][ 291 ],
   alphaCSR[ 61 ][ 292 ],
   alphaCSR[ 61 ][ 293 ],
   alphaCSR[ 61 ][ 294 ],
   alphaCSR[ 61 ][ 295 ],
   alphaCSR[ 61 ][ 296 ],
   alphaCSR[ 61 ][ 297 ],
   alphaCSR[ 61 ][ 298 ],
   alphaCSR[ 61 ][ 299 ],
   alphaCSR[ 61 ][ 300 ],
   alphaCSR[ 61 ][ 301 ],
   alphaCSR[ 61 ][ 302 ],
   alphaCSR[ 61 ][ 303 ],
   alphaCSR[ 61 ][ 304 ],
   alphaCSR[ 61 ][ 305 ],
   alphaCSR[ 61 ][ 306 ],
   alphaCSR[ 61 ][ 307 ],
   alphaCSR[ 61 ][ 308 ],
   alphaCSR[ 61 ][ 309 ],
   alphaCSR[ 61 ][ 310 ],
   alphaCSR[ 61 ][ 311 ],
   alphaCSR[ 61 ][ 312 ],
   alphaCSR[ 61 ][ 313 ],
   alphaCSR[ 61 ][ 314 ],
   alphaCSR[ 61 ][ 315 ],
   alphaCSR[ 61 ][ 316 ],
   alphaCSR[ 61 ][ 317 ],
   alphaCSR[ 61 ][ 318 ],
   alphaCSR[ 61 ][ 319 ],
   alphaCSR[ 61 ][ 320 ],
   alphaCSR[ 61 ][ 321 ],
   alphaCSR[ 61 ][ 322 ],
   alphaCSR[ 61 ][ 323 ],
   alphaCSR[ 61 ][ 324 ],
   alphaCSR[ 61 ][ 325 ],
   alphaCSR[ 61 ][ 326 ],
   alphaCSR[ 61 ][ 327 ],
   alphaCSR[ 61 ][ 328 ],
   alphaCSR[ 61 ][ 329 ],
   alphaCSR[ 61 ][ 330 ],
   alphaCSR[ 61 ][ 331 ],
   alphaCSR[ 61 ][ 332 ],
   alphaCSR[ 61 ][ 333 ],
   alphaCSR[ 61 ][ 334 ],
   alphaCSR[ 61 ][ 335 ],
   alphaCSR[ 61 ][ 336 ],
   alphaCSR[ 61 ][ 337 ],
   alphaCSR[ 61 ][ 338 ],
   alphaCSR[ 61 ][ 339 ],
   alphaCSR[ 61 ][ 340 ],
   alphaCSR[ 61 ][ 341 ],
   alphaCSR[ 61 ][ 342 ],
   alphaCSR[ 61 ][ 343 ],
   alphaCSR[ 61 ][ 344 ],
   alphaCSR[ 61 ][ 345 ],
   alphaCSR[ 61 ][ 346 ],
   alphaCSR[ 61 ][ 347 ],
   alphaCSR[ 61 ][ 348 ],
   alphaCSR[ 61 ][ 349 ],
   alphaCSR[ 61 ][ 350 ],
   alphaCSR[ 61 ][ 351 ],
   alphaCSR[ 61 ][ 352 ],
   alphaCSR[ 61 ][ 353 ],
   alphaCSR[ 61 ][ 354 ],
   alphaCSR[ 61 ][ 355 ],
   alphaCSR[ 61 ][ 356 ],
   alphaCSR[ 61 ][ 357 ],
   alphaCSR[ 61 ][ 358 ],
   alphaCSR[ 61 ][ 359 ],
   alphaCSR[ 61 ][ 360 ],
   alphaCSR[ 61 ][ 361 ],
   alphaCSR[ 61 ][ 362 ],
   alphaCSR[ 61 ][ 363 ],
   alphaCSR[ 61 ][ 364 ],
   alphaCSR[ 61 ][ 365 ],
   alphaCSR[ 61 ][ 366 ],
   alphaCSR[ 61 ][ 367 ],
   alphaCSR[ 61 ][ 368 ],
   alphaCSR[ 61 ][ 369 ],
   alphaCSR[ 61 ][ 370 ],
   alphaCSR[ 61 ][ 371 ],
   alphaCSR[ 61 ][ 372 ],
   alphaCSR[ 61 ][ 373 ],
   alphaCSR[ 61 ][ 374 ],
   alphaCSR[ 61 ][ 375 ],
   alphaCSR[ 61 ][ 376 ],
   alphaCSR[ 61 ][ 377 ],
   alphaCSR[ 61 ][ 378 ],
   alphaCSR[ 61 ][ 379 ],
   alphaCSR[ 61 ][ 380 ],
   alphaCSR[ 61 ][ 381 ],
   alphaCSR[ 61 ][ 382 ],
   alphaCSR[ 61 ][ 383 ],
   alphaCSR[ 62 ][ 0 ],
   alphaCSR[ 62 ][ 1 ],
   alphaCSR[ 62 ][ 2 ],
   alphaCSR[ 62 ][ 3 ],
   alphaCSR[ 62 ][ 4 ],
   alphaCSR[ 62 ][ 5 ],
   alphaCSR[ 62 ][ 6 ],
   alphaCSR[ 62 ][ 7 ],
   alphaCSR[ 62 ][ 8 ],
   alphaCSR[ 62 ][ 9 ],
   alphaCSR[ 62 ][ 10 ],
   alphaCSR[ 62 ][ 11 ],
   alphaCSR[ 62 ][ 12 ],
   alphaCSR[ 62 ][ 13 ],
   alphaCSR[ 62 ][ 14 ],
   alphaCSR[ 62 ][ 15 ],
   alphaCSR[ 62 ][ 16 ],
   alphaCSR[ 62 ][ 17 ],
   alphaCSR[ 62 ][ 18 ],
   alphaCSR[ 62 ][ 19 ],
   alphaCSR[ 62 ][ 20 ],
   alphaCSR[ 62 ][ 21 ],
   alphaCSR[ 62 ][ 22 ],
   alphaCSR[ 62 ][ 23 ],
   alphaCSR[ 62 ][ 24 ],
   alphaCSR[ 62 ][ 25 ],
   alphaCSR[ 62 ][ 26 ],
   alphaCSR[ 62 ][ 27 ],
   alphaCSR[ 62 ][ 28 ],
   alphaCSR[ 62 ][ 29 ],
   alphaCSR[ 62 ][ 30 ],
   alphaCSR[ 62 ][ 31 ],
   alphaCSR[ 62 ][ 32 ],
   alphaCSR[ 62 ][ 33 ],
   alphaCSR[ 62 ][ 34 ],
   alphaCSR[ 62 ][ 35 ],
   alphaCSR[ 62 ][ 36 ],
   alphaCSR[ 62 ][ 37 ],
   alphaCSR[ 62 ][ 38 ],
   alphaCSR[ 62 ][ 39 ],
   alphaCSR[ 62 ][ 40 ],
   alphaCSR[ 62 ][ 41 ],
   alphaCSR[ 62 ][ 42 ],
   alphaCSR[ 62 ][ 43 ],
   alphaCSR[ 62 ][ 44 ],
   alphaCSR[ 62 ][ 45 ],
   alphaCSR[ 62 ][ 46 ],
   alphaCSR[ 62 ][ 47 ],
   alphaCSR[ 62 ][ 48 ],
   alphaCSR[ 62 ][ 49 ],
   alphaCSR[ 62 ][ 50 ],
   alphaCSR[ 62 ][ 51 ],
   alphaCSR[ 62 ][ 52 ],
   alphaCSR[ 62 ][ 53 ],
   alphaCSR[ 62 ][ 54 ],
   alphaCSR[ 62 ][ 55 ],
   alphaCSR[ 62 ][ 56 ],
   alphaCSR[ 62 ][ 57 ],
   alphaCSR[ 62 ][ 58 ],
   alphaCSR[ 62 ][ 59 ],
   alphaCSR[ 62 ][ 60 ],
   alphaCSR[ 62 ][ 61 ],
   alphaCSR[ 62 ][ 62 ],
   alphaCSR[ 62 ][ 63 ],
   alphaCSR[ 62 ][ 64 ],
   alphaCSR[ 62 ][ 65 ],
   alphaCSR[ 62 ][ 66 ],
   alphaCSR[ 62 ][ 67 ],
   alphaCSR[ 62 ][ 68 ],
   alphaCSR[ 62 ][ 69 ],
   alphaCSR[ 62 ][ 70 ],
   alphaCSR[ 62 ][ 71 ],
   alphaCSR[ 62 ][ 72 ],
   alphaCSR[ 62 ][ 73 ],
   alphaCSR[ 62 ][ 74 ],
   alphaCSR[ 62 ][ 75 ],
   alphaCSR[ 62 ][ 76 ],
   alphaCSR[ 62 ][ 77 ],
   alphaCSR[ 62 ][ 78 ],
   alphaCSR[ 62 ][ 79 ],
   alphaCSR[ 62 ][ 80 ],
   alphaCSR[ 62 ][ 81 ],
   alphaCSR[ 62 ][ 82 ],
   alphaCSR[ 62 ][ 83 ],
   alphaCSR[ 62 ][ 84 ],
   alphaCSR[ 62 ][ 85 ],
   alphaCSR[ 62 ][ 86 ],
   alphaCSR[ 62 ][ 87 ],
   alphaCSR[ 62 ][ 88 ],
   alphaCSR[ 62 ][ 89 ],
   alphaCSR[ 62 ][ 90 ],
   alphaCSR[ 62 ][ 91 ],
   alphaCSR[ 62 ][ 92 ],
   alphaCSR[ 62 ][ 93 ],
   alphaCSR[ 62 ][ 94 ],
   alphaCSR[ 62 ][ 95 ],
   alphaCSR[ 62 ][ 96 ],
   alphaCSR[ 62 ][ 97 ],
   alphaCSR[ 62 ][ 98 ],
   alphaCSR[ 62 ][ 99 ],
   alphaCSR[ 62 ][ 100 ],
   alphaCSR[ 62 ][ 101 ],
   alphaCSR[ 62 ][ 102 ],
   alphaCSR[ 62 ][ 103 ],
   alphaCSR[ 62 ][ 104 ],
   alphaCSR[ 62 ][ 105 ],
   alphaCSR[ 62 ][ 106 ],
   alphaCSR[ 62 ][ 107 ],
   alphaCSR[ 62 ][ 108 ],
   alphaCSR[ 62 ][ 109 ],
   alphaCSR[ 62 ][ 110 ],
   alphaCSR[ 62 ][ 111 ],
   alphaCSR[ 62 ][ 112 ],
   alphaCSR[ 62 ][ 113 ],
   alphaCSR[ 62 ][ 114 ],
   alphaCSR[ 62 ][ 115 ],
   alphaCSR[ 62 ][ 116 ],
   alphaCSR[ 62 ][ 117 ],
   alphaCSR[ 62 ][ 118 ],
   alphaCSR[ 62 ][ 119 ],
   alphaCSR[ 62 ][ 120 ],
   alphaCSR[ 62 ][ 121 ],
   alphaCSR[ 62 ][ 122 ],
   alphaCSR[ 62 ][ 123 ],
   alphaCSR[ 62 ][ 124 ],
   alphaCSR[ 62 ][ 125 ],
   alphaCSR[ 62 ][ 126 ],
   alphaCSR[ 62 ][ 127 ],
   alphaCSR[ 62 ][ 128 ],
   alphaCSR[ 62 ][ 129 ],
   alphaCSR[ 62 ][ 130 ],
   alphaCSR[ 62 ][ 131 ],
   alphaCSR[ 62 ][ 132 ],
   alphaCSR[ 62 ][ 133 ],
   alphaCSR[ 62 ][ 134 ],
   alphaCSR[ 62 ][ 135 ],
   alphaCSR[ 62 ][ 136 ],
   alphaCSR[ 62 ][ 137 ],
   alphaCSR[ 62 ][ 138 ],
   alphaCSR[ 62 ][ 139 ],
   alphaCSR[ 62 ][ 140 ],
   alphaCSR[ 62 ][ 141 ],
   alphaCSR[ 62 ][ 142 ],
   alphaCSR[ 62 ][ 143 ],
   alphaCSR[ 62 ][ 144 ],
   alphaCSR[ 62 ][ 145 ],
   alphaCSR[ 62 ][ 146 ],
   alphaCSR[ 62 ][ 147 ],
   alphaCSR[ 62 ][ 148 ],
   alphaCSR[ 62 ][ 149 ],
   alphaCSR[ 62 ][ 150 ],
   alphaCSR[ 62 ][ 151 ],
   alphaCSR[ 62 ][ 152 ],
   alphaCSR[ 62 ][ 153 ],
   alphaCSR[ 62 ][ 154 ],
   alphaCSR[ 62 ][ 155 ],
   alphaCSR[ 62 ][ 156 ],
   alphaCSR[ 62 ][ 157 ],
   alphaCSR[ 62 ][ 158 ],
   alphaCSR[ 62 ][ 159 ],
   alphaCSR[ 62 ][ 160 ],
   alphaCSR[ 62 ][ 161 ],
   alphaCSR[ 62 ][ 162 ],
   alphaCSR[ 62 ][ 163 ],
   alphaCSR[ 62 ][ 164 ],
   alphaCSR[ 62 ][ 165 ],
   alphaCSR[ 62 ][ 166 ],
   alphaCSR[ 62 ][ 167 ],
   alphaCSR[ 62 ][ 168 ],
   alphaCSR[ 62 ][ 169 ],
   alphaCSR[ 62 ][ 170 ],
   alphaCSR[ 62 ][ 171 ],
   alphaCSR[ 62 ][ 172 ],
   alphaCSR[ 62 ][ 173 ],
   alphaCSR[ 62 ][ 174 ],
   alphaCSR[ 62 ][ 175 ],
   alphaCSR[ 62 ][ 176 ],
   alphaCSR[ 62 ][ 177 ],
   alphaCSR[ 62 ][ 178 ],
   alphaCSR[ 62 ][ 179 ],
   alphaCSR[ 62 ][ 180 ],
   alphaCSR[ 62 ][ 181 ],
   alphaCSR[ 62 ][ 182 ],
   alphaCSR[ 62 ][ 183 ],
   alphaCSR[ 62 ][ 184 ],
   alphaCSR[ 62 ][ 185 ],
   alphaCSR[ 62 ][ 186 ],
   alphaCSR[ 62 ][ 187 ],
   alphaCSR[ 62 ][ 188 ],
   alphaCSR[ 62 ][ 189 ],
   alphaCSR[ 62 ][ 190 ],
   alphaCSR[ 62 ][ 191 ],
   alphaCSR[ 62 ][ 192 ],
   alphaCSR[ 62 ][ 193 ],
   alphaCSR[ 62 ][ 194 ],
   alphaCSR[ 62 ][ 195 ],
   alphaCSR[ 62 ][ 196 ],
   alphaCSR[ 62 ][ 197 ],
   alphaCSR[ 62 ][ 198 ],
   alphaCSR[ 62 ][ 199 ],
   alphaCSR[ 62 ][ 200 ],
   alphaCSR[ 62 ][ 201 ],
   alphaCSR[ 62 ][ 202 ],
   alphaCSR[ 62 ][ 203 ],
   alphaCSR[ 62 ][ 204 ],
   alphaCSR[ 62 ][ 205 ],
   alphaCSR[ 62 ][ 206 ],
   alphaCSR[ 62 ][ 207 ],
   alphaCSR[ 62 ][ 208 ],
   alphaCSR[ 62 ][ 209 ],
   alphaCSR[ 62 ][ 210 ],
   alphaCSR[ 62 ][ 211 ],
   alphaCSR[ 62 ][ 212 ],
   alphaCSR[ 62 ][ 213 ],
   alphaCSR[ 62 ][ 214 ],
   alphaCSR[ 62 ][ 215 ],
   alphaCSR[ 62 ][ 216 ],
   alphaCSR[ 62 ][ 217 ],
   alphaCSR[ 62 ][ 218 ],
   alphaCSR[ 62 ][ 219 ],
   alphaCSR[ 62 ][ 220 ],
   alphaCSR[ 62 ][ 221 ],
   alphaCSR[ 62 ][ 222 ],
   alphaCSR[ 62 ][ 223 ],
   alphaCSR[ 62 ][ 224 ],
   alphaCSR[ 62 ][ 225 ],
   alphaCSR[ 62 ][ 226 ],
   alphaCSR[ 62 ][ 227 ],
   alphaCSR[ 62 ][ 228 ],
   alphaCSR[ 62 ][ 229 ],
   alphaCSR[ 62 ][ 230 ],
   alphaCSR[ 62 ][ 231 ],
   alphaCSR[ 62 ][ 232 ],
   alphaCSR[ 62 ][ 233 ],
   alphaCSR[ 62 ][ 234 ],
   alphaCSR[ 62 ][ 235 ],
   alphaCSR[ 62 ][ 236 ],
   alphaCSR[ 62 ][ 237 ],
   alphaCSR[ 62 ][ 238 ],
   alphaCSR[ 62 ][ 239 ],
   alphaCSR[ 62 ][ 240 ],
   alphaCSR[ 62 ][ 241 ],
   alphaCSR[ 62 ][ 242 ],
   alphaCSR[ 62 ][ 243 ],
   alphaCSR[ 62 ][ 244 ],
   alphaCSR[ 62 ][ 245 ],
   alphaCSR[ 62 ][ 246 ],
   alphaCSR[ 62 ][ 247 ],
   alphaCSR[ 62 ][ 248 ],
   alphaCSR[ 62 ][ 249 ],
   alphaCSR[ 62 ][ 250 ],
   alphaCSR[ 62 ][ 251 ],
   alphaCSR[ 62 ][ 252 ],
   alphaCSR[ 62 ][ 253 ],
   alphaCSR[ 62 ][ 254 ],
   alphaCSR[ 62 ][ 255 ],
   alphaCSR[ 62 ][ 256 ],
   alphaCSR[ 62 ][ 257 ],
   alphaCSR[ 62 ][ 258 ],
   alphaCSR[ 62 ][ 259 ],
   alphaCSR[ 62 ][ 260 ],
   alphaCSR[ 62 ][ 261 ],
   alphaCSR[ 62 ][ 262 ],
   alphaCSR[ 62 ][ 263 ],
   alphaCSR[ 62 ][ 264 ],
   alphaCSR[ 62 ][ 265 ],
   alphaCSR[ 62 ][ 266 ],
   alphaCSR[ 62 ][ 267 ],
   alphaCSR[ 62 ][ 268 ],
   alphaCSR[ 62 ][ 269 ],
   alphaCSR[ 62 ][ 270 ],
   alphaCSR[ 62 ][ 271 ],
   alphaCSR[ 62 ][ 272 ],
   alphaCSR[ 62 ][ 273 ],
   alphaCSR[ 62 ][ 274 ],
   alphaCSR[ 62 ][ 275 ],
   alphaCSR[ 62 ][ 276 ],
   alphaCSR[ 62 ][ 277 ],
   alphaCSR[ 62 ][ 278 ],
   alphaCSR[ 62 ][ 279 ],
   alphaCSR[ 62 ][ 280 ],
   alphaCSR[ 62 ][ 281 ],
   alphaCSR[ 62 ][ 282 ],
   alphaCSR[ 62 ][ 283 ],
   alphaCSR[ 62 ][ 284 ],
   alphaCSR[ 62 ][ 285 ],
   alphaCSR[ 62 ][ 286 ],
   alphaCSR[ 62 ][ 287 ],
   alphaCSR[ 62 ][ 288 ],
   alphaCSR[ 62 ][ 289 ],
   alphaCSR[ 62 ][ 290 ],
   alphaCSR[ 62 ][ 291 ],
   alphaCSR[ 62 ][ 292 ],
   alphaCSR[ 62 ][ 293 ],
   alphaCSR[ 62 ][ 294 ],
   alphaCSR[ 62 ][ 295 ],
   alphaCSR[ 62 ][ 296 ],
   alphaCSR[ 62 ][ 297 ],
   alphaCSR[ 62 ][ 298 ],
   alphaCSR[ 62 ][ 299 ],
   alphaCSR[ 62 ][ 300 ],
   alphaCSR[ 62 ][ 301 ],
   alphaCSR[ 62 ][ 302 ],
   alphaCSR[ 62 ][ 303 ],
   alphaCSR[ 62 ][ 304 ],
   alphaCSR[ 62 ][ 305 ],
   alphaCSR[ 62 ][ 306 ],
   alphaCSR[ 62 ][ 307 ],
   alphaCSR[ 62 ][ 308 ],
   alphaCSR[ 62 ][ 309 ],
   alphaCSR[ 62 ][ 310 ],
   alphaCSR[ 62 ][ 311 ],
   alphaCSR[ 62 ][ 312 ],
   alphaCSR[ 62 ][ 313 ],
   alphaCSR[ 62 ][ 314 ],
   alphaCSR[ 62 ][ 315 ],
   alphaCSR[ 62 ][ 316 ],
   alphaCSR[ 62 ][ 317 ],
   alphaCSR[ 62 ][ 318 ],
   alphaCSR[ 62 ][ 319 ],
   alphaCSR[ 62 ][ 320 ],
   alphaCSR[ 62 ][ 321 ],
   alphaCSR[ 62 ][ 322 ],
   alphaCSR[ 62 ][ 323 ],
   alphaCSR[ 62 ][ 324 ],
   alphaCSR[ 62 ][ 325 ],
   alphaCSR[ 62 ][ 326 ],
   alphaCSR[ 62 ][ 327 ],
   alphaCSR[ 62 ][ 328 ],
   alphaCSR[ 62 ][ 329 ],
   alphaCSR[ 62 ][ 330 ],
   alphaCSR[ 62 ][ 331 ],
   alphaCSR[ 62 ][ 332 ],
   alphaCSR[ 62 ][ 333 ],
   alphaCSR[ 62 ][ 334 ],
   alphaCSR[ 62 ][ 335 ],
   alphaCSR[ 62 ][ 336 ],
   alphaCSR[ 62 ][ 337 ],
   alphaCSR[ 62 ][ 338 ],
   alphaCSR[ 62 ][ 339 ],
   alphaCSR[ 62 ][ 340 ],
   alphaCSR[ 62 ][ 341 ],
   alphaCSR[ 62 ][ 342 ],
   alphaCSR[ 62 ][ 343 ],
   alphaCSR[ 62 ][ 344 ],
   alphaCSR[ 62 ][ 345 ],
   alphaCSR[ 62 ][ 346 ],
   alphaCSR[ 62 ][ 347 ],
   alphaCSR[ 62 ][ 348 ],
   alphaCSR[ 62 ][ 349 ],
   alphaCSR[ 62 ][ 350 ],
   alphaCSR[ 62 ][ 351 ],
   alphaCSR[ 62 ][ 352 ],
   alphaCSR[ 62 ][ 353 ],
   alphaCSR[ 62 ][ 354 ],
   alphaCSR[ 62 ][ 355 ],
   alphaCSR[ 62 ][ 356 ],
   alphaCSR[ 62 ][ 357 ],
   alphaCSR[ 62 ][ 358 ],
   alphaCSR[ 62 ][ 359 ],
   alphaCSR[ 62 ][ 360 ],
   alphaCSR[ 62 ][ 361 ],
   alphaCSR[ 62 ][ 362 ],
   alphaCSR[ 62 ][ 363 ],
   alphaCSR[ 62 ][ 364 ],
   alphaCSR[ 62 ][ 365 ],
   alphaCSR[ 62 ][ 366 ],
   alphaCSR[ 62 ][ 367 ],
   alphaCSR[ 62 ][ 368 ],
   alphaCSR[ 62 ][ 369 ],
   alphaCSR[ 62 ][ 370 ],
   alphaCSR[ 62 ][ 371 ],
   alphaCSR[ 62 ][ 372 ],
   alphaCSR[ 62 ][ 373 ],
   alphaCSR[ 62 ][ 374 ],
   alphaCSR[ 62 ][ 375 ],
   alphaCSR[ 62 ][ 376 ],
   alphaCSR[ 62 ][ 377 ],
   alphaCSR[ 62 ][ 378 ],
   alphaCSR[ 62 ][ 379 ],
   alphaCSR[ 62 ][ 380 ],
   alphaCSR[ 62 ][ 381 ],
   alphaCSR[ 62 ][ 382 ],
   alphaCSR[ 62 ][ 383 ],
   alphaCSR[ 63 ][ 0 ],
   alphaCSR[ 63 ][ 1 ],
   alphaCSR[ 63 ][ 2 ],
   alphaCSR[ 63 ][ 3 ],
   alphaCSR[ 63 ][ 4 ],
   alphaCSR[ 63 ][ 5 ],
   alphaCSR[ 63 ][ 6 ],
   alphaCSR[ 63 ][ 7 ],
   alphaCSR[ 63 ][ 8 ],
   alphaCSR[ 63 ][ 9 ],
   alphaCSR[ 63 ][ 10 ],
   alphaCSR[ 63 ][ 11 ],
   alphaCSR[ 63 ][ 12 ],
   alphaCSR[ 63 ][ 13 ],
   alphaCSR[ 63 ][ 14 ],
   alphaCSR[ 63 ][ 15 ],
   alphaCSR[ 63 ][ 16 ],
   alphaCSR[ 63 ][ 17 ],
   alphaCSR[ 63 ][ 18 ],
   alphaCSR[ 63 ][ 19 ],
   alphaCSR[ 63 ][ 20 ],
   alphaCSR[ 63 ][ 21 ],
   alphaCSR[ 63 ][ 22 ],
   alphaCSR[ 63 ][ 23 ],
   alphaCSR[ 63 ][ 24 ],
   alphaCSR[ 63 ][ 25 ],
   alphaCSR[ 63 ][ 26 ],
   alphaCSR[ 63 ][ 27 ],
   alphaCSR[ 63 ][ 28 ],
   alphaCSR[ 63 ][ 29 ],
   alphaCSR[ 63 ][ 30 ],
   alphaCSR[ 63 ][ 31 ],
   alphaCSR[ 63 ][ 32 ],
   alphaCSR[ 63 ][ 33 ],
   alphaCSR[ 63 ][ 34 ],
   alphaCSR[ 63 ][ 35 ],
   alphaCSR[ 63 ][ 36 ],
   alphaCSR[ 63 ][ 37 ],
   alphaCSR[ 63 ][ 38 ],
   alphaCSR[ 63 ][ 39 ],
   alphaCSR[ 63 ][ 40 ],
   alphaCSR[ 63 ][ 41 ],
   alphaCSR[ 63 ][ 42 ],
   alphaCSR[ 63 ][ 43 ],
   alphaCSR[ 63 ][ 44 ],
   alphaCSR[ 63 ][ 45 ],
   alphaCSR[ 63 ][ 46 ],
   alphaCSR[ 63 ][ 47 ],
   alphaCSR[ 63 ][ 48 ],
   alphaCSR[ 63 ][ 49 ],
   alphaCSR[ 63 ][ 50 ],
   alphaCSR[ 63 ][ 51 ],
   alphaCSR[ 63 ][ 52 ],
   alphaCSR[ 63 ][ 53 ],
   alphaCSR[ 63 ][ 54 ],
   alphaCSR[ 63 ][ 55 ],
   alphaCSR[ 63 ][ 56 ],
   alphaCSR[ 63 ][ 57 ],
   alphaCSR[ 63 ][ 58 ],
   alphaCSR[ 63 ][ 59 ],
   alphaCSR[ 63 ][ 60 ],
   alphaCSR[ 63 ][ 61 ],
   alphaCSR[ 63 ][ 62 ],
   alphaCSR[ 63 ][ 63 ],
   alphaCSR[ 63 ][ 64 ],
   alphaCSR[ 63 ][ 65 ],
   alphaCSR[ 63 ][ 66 ],
   alphaCSR[ 63 ][ 67 ],
   alphaCSR[ 63 ][ 68 ],
   alphaCSR[ 63 ][ 69 ],
   alphaCSR[ 63 ][ 70 ],
   alphaCSR[ 63 ][ 71 ],
   alphaCSR[ 63 ][ 72 ],
   alphaCSR[ 63 ][ 73 ],
   alphaCSR[ 63 ][ 74 ],
   alphaCSR[ 63 ][ 75 ],
   alphaCSR[ 63 ][ 76 ],
   alphaCSR[ 63 ][ 77 ],
   alphaCSR[ 63 ][ 78 ],
   alphaCSR[ 63 ][ 79 ],
   alphaCSR[ 63 ][ 80 ],
   alphaCSR[ 63 ][ 81 ],
   alphaCSR[ 63 ][ 82 ],
   alphaCSR[ 63 ][ 83 ],
   alphaCSR[ 63 ][ 84 ],
   alphaCSR[ 63 ][ 85 ],
   alphaCSR[ 63 ][ 86 ],
   alphaCSR[ 63 ][ 87 ],
   alphaCSR[ 63 ][ 88 ],
   alphaCSR[ 63 ][ 89 ],
   alphaCSR[ 63 ][ 90 ],
   alphaCSR[ 63 ][ 91 ],
   alphaCSR[ 63 ][ 92 ],
   alphaCSR[ 63 ][ 93 ],
   alphaCSR[ 63 ][ 94 ],
   alphaCSR[ 63 ][ 95 ],
   alphaCSR[ 63 ][ 96 ],
   alphaCSR[ 63 ][ 97 ],
   alphaCSR[ 63 ][ 98 ],
   alphaCSR[ 63 ][ 99 ],
   alphaCSR[ 63 ][ 100 ],
   alphaCSR[ 63 ][ 101 ],
   alphaCSR[ 63 ][ 102 ],
   alphaCSR[ 63 ][ 103 ],
   alphaCSR[ 63 ][ 104 ],
   alphaCSR[ 63 ][ 105 ],
   alphaCSR[ 63 ][ 106 ],
   alphaCSR[ 63 ][ 107 ],
   alphaCSR[ 63 ][ 108 ],
   alphaCSR[ 63 ][ 109 ],
   alphaCSR[ 63 ][ 110 ],
   alphaCSR[ 63 ][ 111 ],
   alphaCSR[ 63 ][ 112 ],
   alphaCSR[ 63 ][ 113 ],
   alphaCSR[ 63 ][ 114 ],
   alphaCSR[ 63 ][ 115 ],
   alphaCSR[ 63 ][ 116 ],
   alphaCSR[ 63 ][ 117 ],
   alphaCSR[ 63 ][ 118 ],
   alphaCSR[ 63 ][ 119 ],
   alphaCSR[ 63 ][ 120 ],
   alphaCSR[ 63 ][ 121 ],
   alphaCSR[ 63 ][ 122 ],
   alphaCSR[ 63 ][ 123 ],
   alphaCSR[ 63 ][ 124 ],
   alphaCSR[ 63 ][ 125 ],
   alphaCSR[ 63 ][ 126 ],
   alphaCSR[ 63 ][ 127 ],
   alphaCSR[ 63 ][ 128 ],
   alphaCSR[ 63 ][ 129 ],
   alphaCSR[ 63 ][ 130 ],
   alphaCSR[ 63 ][ 131 ],
   alphaCSR[ 63 ][ 132 ],
   alphaCSR[ 63 ][ 133 ],
   alphaCSR[ 63 ][ 134 ],
   alphaCSR[ 63 ][ 135 ],
   alphaCSR[ 63 ][ 136 ],
   alphaCSR[ 63 ][ 137 ],
   alphaCSR[ 63 ][ 138 ],
   alphaCSR[ 63 ][ 139 ],
   alphaCSR[ 63 ][ 140 ],
   alphaCSR[ 63 ][ 141 ],
   alphaCSR[ 63 ][ 142 ],
   alphaCSR[ 63 ][ 143 ],
   alphaCSR[ 63 ][ 144 ],
   alphaCSR[ 63 ][ 145 ],
   alphaCSR[ 63 ][ 146 ],
   alphaCSR[ 63 ][ 147 ],
   alphaCSR[ 63 ][ 148 ],
   alphaCSR[ 63 ][ 149 ],
   alphaCSR[ 63 ][ 150 ],
   alphaCSR[ 63 ][ 151 ],
   alphaCSR[ 63 ][ 152 ],
   alphaCSR[ 63 ][ 153 ],
   alphaCSR[ 63 ][ 154 ],
   alphaCSR[ 63 ][ 155 ],
   alphaCSR[ 63 ][ 156 ],
   alphaCSR[ 63 ][ 157 ],
   alphaCSR[ 63 ][ 158 ],
   alphaCSR[ 63 ][ 159 ],
   alphaCSR[ 63 ][ 160 ],
   alphaCSR[ 63 ][ 161 ],
   alphaCSR[ 63 ][ 162 ],
   alphaCSR[ 63 ][ 163 ],
   alphaCSR[ 63 ][ 164 ],
   alphaCSR[ 63 ][ 165 ],
   alphaCSR[ 63 ][ 166 ],
   alphaCSR[ 63 ][ 167 ],
   alphaCSR[ 63 ][ 168 ],
   alphaCSR[ 63 ][ 169 ],
   alphaCSR[ 63 ][ 170 ],
   alphaCSR[ 63 ][ 171 ],
   alphaCSR[ 63 ][ 172 ],
   alphaCSR[ 63 ][ 173 ],
   alphaCSR[ 63 ][ 174 ],
   alphaCSR[ 63 ][ 175 ],
   alphaCSR[ 63 ][ 176 ],
   alphaCSR[ 63 ][ 177 ],
   alphaCSR[ 63 ][ 178 ],
   alphaCSR[ 63 ][ 179 ],
   alphaCSR[ 63 ][ 180 ],
   alphaCSR[ 63 ][ 181 ],
   alphaCSR[ 63 ][ 182 ],
   alphaCSR[ 63 ][ 183 ],
   alphaCSR[ 63 ][ 184 ],
   alphaCSR[ 63 ][ 185 ],
   alphaCSR[ 63 ][ 186 ],
   alphaCSR[ 63 ][ 187 ],
   alphaCSR[ 63 ][ 188 ],
   alphaCSR[ 63 ][ 189 ],
   alphaCSR[ 63 ][ 190 ],
   alphaCSR[ 63 ][ 191 ],
   alphaCSR[ 63 ][ 192 ],
   alphaCSR[ 63 ][ 193 ],
   alphaCSR[ 63 ][ 194 ],
   alphaCSR[ 63 ][ 195 ],
   alphaCSR[ 63 ][ 196 ],
   alphaCSR[ 63 ][ 197 ],
   alphaCSR[ 63 ][ 198 ],
   alphaCSR[ 63 ][ 199 ],
   alphaCSR[ 63 ][ 200 ],
   alphaCSR[ 63 ][ 201 ],
   alphaCSR[ 63 ][ 202 ],
   alphaCSR[ 63 ][ 203 ],
   alphaCSR[ 63 ][ 204 ],
   alphaCSR[ 63 ][ 205 ],
   alphaCSR[ 63 ][ 206 ],
   alphaCSR[ 63 ][ 207 ],
   alphaCSR[ 63 ][ 208 ],
   alphaCSR[ 63 ][ 209 ],
   alphaCSR[ 63 ][ 210 ],
   alphaCSR[ 63 ][ 211 ],
   alphaCSR[ 63 ][ 212 ],
   alphaCSR[ 63 ][ 213 ],
   alphaCSR[ 63 ][ 214 ],
   alphaCSR[ 63 ][ 215 ],
   alphaCSR[ 63 ][ 216 ],
   alphaCSR[ 63 ][ 217 ],
   alphaCSR[ 63 ][ 218 ],
   alphaCSR[ 63 ][ 219 ],
   alphaCSR[ 63 ][ 220 ],
   alphaCSR[ 63 ][ 221 ],
   alphaCSR[ 63 ][ 222 ],
   alphaCSR[ 63 ][ 223 ],
   alphaCSR[ 63 ][ 224 ],
   alphaCSR[ 63 ][ 225 ],
   alphaCSR[ 63 ][ 226 ],
   alphaCSR[ 63 ][ 227 ],
   alphaCSR[ 63 ][ 228 ],
   alphaCSR[ 63 ][ 229 ],
   alphaCSR[ 63 ][ 230 ],
   alphaCSR[ 63 ][ 231 ],
   alphaCSR[ 63 ][ 232 ],
   alphaCSR[ 63 ][ 233 ],
   alphaCSR[ 63 ][ 234 ],
   alphaCSR[ 63 ][ 235 ],
   alphaCSR[ 63 ][ 236 ],
   alphaCSR[ 63 ][ 237 ],
   alphaCSR[ 63 ][ 238 ],
   alphaCSR[ 63 ][ 239 ],
   alphaCSR[ 63 ][ 240 ],
   alphaCSR[ 63 ][ 241 ],
   alphaCSR[ 63 ][ 242 ],
   alphaCSR[ 63 ][ 243 ],
   alphaCSR[ 63 ][ 244 ],
   alphaCSR[ 63 ][ 245 ],
   alphaCSR[ 63 ][ 246 ],
   alphaCSR[ 63 ][ 247 ],
   alphaCSR[ 63 ][ 248 ],
   alphaCSR[ 63 ][ 249 ],
   alphaCSR[ 63 ][ 250 ],
   alphaCSR[ 63 ][ 251 ],
   alphaCSR[ 63 ][ 252 ],
   alphaCSR[ 63 ][ 253 ],
   alphaCSR[ 63 ][ 254 ],
   alphaCSR[ 63 ][ 255 ],
   alphaCSR[ 63 ][ 256 ],
   alphaCSR[ 63 ][ 257 ],
   alphaCSR[ 63 ][ 258 ],
   alphaCSR[ 63 ][ 259 ],
   alphaCSR[ 63 ][ 260 ],
   alphaCSR[ 63 ][ 261 ],
   alphaCSR[ 63 ][ 262 ],
   alphaCSR[ 63 ][ 263 ],
   alphaCSR[ 63 ][ 264 ],
   alphaCSR[ 63 ][ 265 ],
   alphaCSR[ 63 ][ 266 ],
   alphaCSR[ 63 ][ 267 ],
   alphaCSR[ 63 ][ 268 ],
   alphaCSR[ 63 ][ 269 ],
   alphaCSR[ 63 ][ 270 ],
   alphaCSR[ 63 ][ 271 ],
   alphaCSR[ 63 ][ 272 ],
   alphaCSR[ 63 ][ 273 ],
   alphaCSR[ 63 ][ 274 ],
   alphaCSR[ 63 ][ 275 ],
   alphaCSR[ 63 ][ 276 ],
   alphaCSR[ 63 ][ 277 ],
   alphaCSR[ 63 ][ 278 ],
   alphaCSR[ 63 ][ 279 ],
   alphaCSR[ 63 ][ 280 ],
   alphaCSR[ 63 ][ 281 ],
   alphaCSR[ 63 ][ 282 ],
   alphaCSR[ 63 ][ 283 ],
   alphaCSR[ 63 ][ 284 ],
   alphaCSR[ 63 ][ 285 ],
   alphaCSR[ 63 ][ 286 ],
   alphaCSR[ 63 ][ 287 ],
   alphaCSR[ 63 ][ 288 ],
   alphaCSR[ 63 ][ 289 ],
   alphaCSR[ 63 ][ 290 ],
   alphaCSR[ 63 ][ 291 ],
   alphaCSR[ 63 ][ 292 ],
   alphaCSR[ 63 ][ 293 ],
   alphaCSR[ 63 ][ 294 ],
   alphaCSR[ 63 ][ 295 ],
   alphaCSR[ 63 ][ 296 ],
   alphaCSR[ 63 ][ 297 ],
   alphaCSR[ 63 ][ 298 ],
   alphaCSR[ 63 ][ 299 ],
   alphaCSR[ 63 ][ 300 ],
   alphaCSR[ 63 ][ 301 ],
   alphaCSR[ 63 ][ 302 ],
   alphaCSR[ 63 ][ 303 ],
   alphaCSR[ 63 ][ 304 ],
   alphaCSR[ 63 ][ 305 ],
   alphaCSR[ 63 ][ 306 ],
   alphaCSR[ 63 ][ 307 ],
   alphaCSR[ 63 ][ 308 ],
   alphaCSR[ 63 ][ 309 ],
   alphaCSR[ 63 ][ 310 ],
   alphaCSR[ 63 ][ 311 ],
   alphaCSR[ 63 ][ 312 ],
   alphaCSR[ 63 ][ 313 ],
   alphaCSR[ 63 ][ 314 ],
   alphaCSR[ 63 ][ 315 ],
   alphaCSR[ 63 ][ 316 ],
   alphaCSR[ 63 ][ 317 ],
   alphaCSR[ 63 ][ 318 ],
   alphaCSR[ 63 ][ 319 ],
   alphaCSR[ 63 ][ 320 ],
   alphaCSR[ 63 ][ 321 ],
   alphaCSR[ 63 ][ 322 ],
   alphaCSR[ 63 ][ 323 ],
   alphaCSR[ 63 ][ 324 ],
   alphaCSR[ 63 ][ 325 ],
   alphaCSR[ 63 ][ 326 ],
   alphaCSR[ 63 ][ 327 ],
   alphaCSR[ 63 ][ 328 ],
   alphaCSR[ 63 ][ 329 ],
   alphaCSR[ 63 ][ 330 ],
   alphaCSR[ 63 ][ 331 ],
   alphaCSR[ 63 ][ 332 ],
   alphaCSR[ 63 ][ 333 ],
   alphaCSR[ 63 ][ 334 ],
   alphaCSR[ 63 ][ 335 ],
   alphaCSR[ 63 ][ 336 ],
   alphaCSR[ 63 ][ 337 ],
   alphaCSR[ 63 ][ 338 ],
   alphaCSR[ 63 ][ 339 ],
   alphaCSR[ 63 ][ 340 ],
   alphaCSR[ 63 ][ 341 ],
   alphaCSR[ 63 ][ 342 ],
   alphaCSR[ 63 ][ 343 ],
   alphaCSR[ 63 ][ 344 ],
   alphaCSR[ 63 ][ 345 ],
   alphaCSR[ 63 ][ 346 ],
   alphaCSR[ 63 ][ 347 ],
   alphaCSR[ 63 ][ 348 ],
   alphaCSR[ 63 ][ 349 ],
   alphaCSR[ 63 ][ 350 ],
   alphaCSR[ 63 ][ 351 ],
   alphaCSR[ 63 ][ 352 ],
   alphaCSR[ 63 ][ 353 ],
   alphaCSR[ 63 ][ 354 ],
   alphaCSR[ 63 ][ 355 ],
   alphaCSR[ 63 ][ 356 ],
   alphaCSR[ 63 ][ 357 ],
   alphaCSR[ 63 ][ 358 ],
   alphaCSR[ 63 ][ 359 ],
   alphaCSR[ 63 ][ 360 ],
   alphaCSR[ 63 ][ 361 ],
   alphaCSR[ 63 ][ 362 ],
   alphaCSR[ 63 ][ 363 ],
   alphaCSR[ 63 ][ 364 ],
   alphaCSR[ 63 ][ 365 ],
   alphaCSR[ 63 ][ 366 ],
   alphaCSR[ 63 ][ 367 ],
   alphaCSR[ 63 ][ 368 ],
   alphaCSR[ 63 ][ 369 ],
   alphaCSR[ 63 ][ 370 ],
   alphaCSR[ 63 ][ 371 ],
   alphaCSR[ 63 ][ 372 ],
   alphaCSR[ 63 ][ 373 ],
   alphaCSR[ 63 ][ 374 ],
   alphaCSR[ 63 ][ 375 ],
   alphaCSR[ 63 ][ 376 ],
   alphaCSR[ 63 ][ 377 ],
   alphaCSR[ 63 ][ 378 ],
   alphaCSR[ 63 ][ 379 ],
   alphaCSR[ 63 ][ 380 ],
   alphaCSR[ 63 ][ 381 ],
   alphaCSR[ 63 ][ 382 ],
   alphaCSR[ 63 ][ 383 ],
   alphaCSR[ 64 ][ 0 ],
   alphaCSR[ 64 ][ 1 ],
   alphaCSR[ 64 ][ 2 ],
   alphaCSR[ 64 ][ 3 ],
   alphaCSR[ 64 ][ 4 ],
   alphaCSR[ 64 ][ 5 ],
   alphaCSR[ 64 ][ 6 ],
   alphaCSR[ 64 ][ 7 ],
   alphaCSR[ 64 ][ 8 ],
   alphaCSR[ 64 ][ 9 ],
   alphaCSR[ 64 ][ 10 ],
   alphaCSR[ 64 ][ 11 ],
   alphaCSR[ 64 ][ 12 ],
   alphaCSR[ 64 ][ 13 ],
   alphaCSR[ 64 ][ 14 ],
   alphaCSR[ 64 ][ 15 ],
   alphaCSR[ 64 ][ 16 ],
   alphaCSR[ 64 ][ 17 ],
   alphaCSR[ 64 ][ 18 ],
   alphaCSR[ 64 ][ 19 ],
   alphaCSR[ 64 ][ 20 ],
   alphaCSR[ 64 ][ 21 ],
   alphaCSR[ 64 ][ 22 ],
   alphaCSR[ 64 ][ 23 ],
   alphaCSR[ 64 ][ 24 ],
   alphaCSR[ 64 ][ 25 ],
   alphaCSR[ 64 ][ 26 ],
   alphaCSR[ 64 ][ 27 ],
   alphaCSR[ 64 ][ 28 ],
   alphaCSR[ 64 ][ 29 ],
   alphaCSR[ 64 ][ 30 ],
   alphaCSR[ 64 ][ 31 ],
   alphaCSR[ 64 ][ 32 ],
   alphaCSR[ 64 ][ 33 ],
   alphaCSR[ 64 ][ 34 ],
   alphaCSR[ 64 ][ 35 ],
   alphaCSR[ 64 ][ 36 ],
   alphaCSR[ 64 ][ 37 ],
   alphaCSR[ 64 ][ 38 ],
   alphaCSR[ 64 ][ 39 ],
   alphaCSR[ 64 ][ 40 ],
   alphaCSR[ 64 ][ 41 ],
   alphaCSR[ 64 ][ 42 ],
   alphaCSR[ 64 ][ 43 ],
   alphaCSR[ 64 ][ 44 ],
   alphaCSR[ 64 ][ 45 ],
   alphaCSR[ 64 ][ 46 ],
   alphaCSR[ 64 ][ 47 ],
   alphaCSR[ 64 ][ 48 ],
   alphaCSR[ 64 ][ 49 ],
   alphaCSR[ 64 ][ 50 ],
   alphaCSR[ 64 ][ 51 ],
   alphaCSR[ 64 ][ 52 ],
   alphaCSR[ 64 ][ 53 ],
   alphaCSR[ 64 ][ 54 ],
   alphaCSR[ 64 ][ 55 ],
   alphaCSR[ 64 ][ 56 ],
   alphaCSR[ 64 ][ 57 ],
   alphaCSR[ 64 ][ 58 ],
   alphaCSR[ 64 ][ 59 ],
   alphaCSR[ 64 ][ 60 ],
   alphaCSR[ 64 ][ 61 ],
   alphaCSR[ 64 ][ 62 ],
   alphaCSR[ 64 ][ 63 ],
   alphaCSR[ 64 ][ 64 ],
   alphaCSR[ 64 ][ 65 ],
   alphaCSR[ 64 ][ 66 ],
   alphaCSR[ 64 ][ 67 ],
   alphaCSR[ 64 ][ 68 ],
   alphaCSR[ 64 ][ 69 ],
   alphaCSR[ 64 ][ 70 ],
   alphaCSR[ 64 ][ 71 ],
   alphaCSR[ 64 ][ 72 ],
   alphaCSR[ 64 ][ 73 ],
   alphaCSR[ 64 ][ 74 ],
   alphaCSR[ 64 ][ 75 ],
   alphaCSR[ 64 ][ 76 ],
   alphaCSR[ 64 ][ 77 ],
   alphaCSR[ 64 ][ 78 ],
   alphaCSR[ 64 ][ 79 ],
   alphaCSR[ 64 ][ 80 ],
   alphaCSR[ 64 ][ 81 ],
   alphaCSR[ 64 ][ 82 ],
   alphaCSR[ 64 ][ 83 ],
   alphaCSR[ 64 ][ 84 ],
   alphaCSR[ 64 ][ 85 ],
   alphaCSR[ 64 ][ 86 ],
   alphaCSR[ 64 ][ 87 ],
   alphaCSR[ 64 ][ 88 ],
   alphaCSR[ 64 ][ 89 ],
   alphaCSR[ 64 ][ 90 ],
   alphaCSR[ 64 ][ 91 ],
   alphaCSR[ 64 ][ 92 ],
   alphaCSR[ 64 ][ 93 ],
   alphaCSR[ 64 ][ 94 ],
   alphaCSR[ 64 ][ 95 ],
   alphaCSR[ 64 ][ 96 ],
   alphaCSR[ 64 ][ 97 ],
   alphaCSR[ 64 ][ 98 ],
   alphaCSR[ 64 ][ 99 ],
   alphaCSR[ 64 ][ 100 ],
   alphaCSR[ 64 ][ 101 ],
   alphaCSR[ 64 ][ 102 ],
   alphaCSR[ 64 ][ 103 ],
   alphaCSR[ 64 ][ 104 ],
   alphaCSR[ 64 ][ 105 ],
   alphaCSR[ 64 ][ 106 ],
   alphaCSR[ 64 ][ 107 ],
   alphaCSR[ 64 ][ 108 ],
   alphaCSR[ 64 ][ 109 ],
   alphaCSR[ 64 ][ 110 ],
   alphaCSR[ 64 ][ 111 ],
   alphaCSR[ 64 ][ 112 ],
   alphaCSR[ 64 ][ 113 ],
   alphaCSR[ 64 ][ 114 ],
   alphaCSR[ 64 ][ 115 ],
   alphaCSR[ 64 ][ 116 ],
   alphaCSR[ 64 ][ 117 ],
   alphaCSR[ 64 ][ 118 ],
   alphaCSR[ 64 ][ 119 ],
   alphaCSR[ 64 ][ 120 ],
   alphaCSR[ 64 ][ 121 ],
   alphaCSR[ 64 ][ 122 ],
   alphaCSR[ 64 ][ 123 ],
   alphaCSR[ 64 ][ 124 ],
   alphaCSR[ 64 ][ 125 ],
   alphaCSR[ 64 ][ 126 ],
   alphaCSR[ 64 ][ 127 ],
   alphaCSR[ 64 ][ 128 ],
   alphaCSR[ 64 ][ 129 ],
   alphaCSR[ 64 ][ 130 ],
   alphaCSR[ 64 ][ 131 ],
   alphaCSR[ 64 ][ 132 ],
   alphaCSR[ 64 ][ 133 ],
   alphaCSR[ 64 ][ 134 ],
   alphaCSR[ 64 ][ 135 ],
   alphaCSR[ 64 ][ 136 ],
   alphaCSR[ 64 ][ 137 ],
   alphaCSR[ 64 ][ 138 ],
   alphaCSR[ 64 ][ 139 ],
   alphaCSR[ 64 ][ 140 ],
   alphaCSR[ 64 ][ 141 ],
   alphaCSR[ 64 ][ 142 ],
   alphaCSR[ 64 ][ 143 ],
   alphaCSR[ 64 ][ 144 ],
   alphaCSR[ 64 ][ 145 ],
   alphaCSR[ 64 ][ 146 ],
   alphaCSR[ 64 ][ 147 ],
   alphaCSR[ 64 ][ 148 ],
   alphaCSR[ 64 ][ 149 ],
   alphaCSR[ 64 ][ 150 ],
   alphaCSR[ 64 ][ 151 ],
   alphaCSR[ 64 ][ 152 ],
   alphaCSR[ 64 ][ 153 ],
   alphaCSR[ 64 ][ 154 ],
   alphaCSR[ 64 ][ 155 ],
   alphaCSR[ 64 ][ 156 ],
   alphaCSR[ 64 ][ 157 ],
   alphaCSR[ 64 ][ 158 ],
   alphaCSR[ 64 ][ 159 ],
   alphaCSR[ 64 ][ 160 ],
   alphaCSR[ 64 ][ 161 ],
   alphaCSR[ 64 ][ 162 ],
   alphaCSR[ 64 ][ 163 ],
   alphaCSR[ 64 ][ 164 ],
   alphaCSR[ 64 ][ 165 ],
   alphaCSR[ 64 ][ 166 ],
   alphaCSR[ 64 ][ 167 ],
   alphaCSR[ 64 ][ 168 ],
   alphaCSR[ 64 ][ 169 ],
   alphaCSR[ 64 ][ 170 ],
   alphaCSR[ 64 ][ 171 ],
   alphaCSR[ 64 ][ 172 ],
   alphaCSR[ 64 ][ 173 ],
   alphaCSR[ 64 ][ 174 ],
   alphaCSR[ 64 ][ 175 ],
   alphaCSR[ 64 ][ 176 ],
   alphaCSR[ 64 ][ 177 ],
   alphaCSR[ 64 ][ 178 ],
   alphaCSR[ 64 ][ 179 ],
   alphaCSR[ 64 ][ 180 ],
   alphaCSR[ 64 ][ 181 ],
   alphaCSR[ 64 ][ 182 ],
   alphaCSR[ 64 ][ 183 ],
   alphaCSR[ 64 ][ 184 ],
   alphaCSR[ 64 ][ 185 ],
   alphaCSR[ 64 ][ 186 ],
   alphaCSR[ 64 ][ 187 ],
   alphaCSR[ 64 ][ 188 ],
   alphaCSR[ 64 ][ 189 ],
   alphaCSR[ 64 ][ 190 ],
   alphaCSR[ 64 ][ 191 ],
   alphaCSR[ 64 ][ 192 ],
   alphaCSR[ 64 ][ 193 ],
   alphaCSR[ 64 ][ 194 ],
   alphaCSR[ 64 ][ 195 ],
   alphaCSR[ 64 ][ 196 ],
   alphaCSR[ 64 ][ 197 ],
   alphaCSR[ 64 ][ 198 ],
   alphaCSR[ 64 ][ 199 ],
   alphaCSR[ 64 ][ 200 ],
   alphaCSR[ 64 ][ 201 ],
   alphaCSR[ 64 ][ 202 ],
   alphaCSR[ 64 ][ 203 ],
   alphaCSR[ 64 ][ 204 ],
   alphaCSR[ 64 ][ 205 ],
   alphaCSR[ 64 ][ 206 ],
   alphaCSR[ 64 ][ 207 ],
   alphaCSR[ 64 ][ 208 ],
   alphaCSR[ 64 ][ 209 ],
   alphaCSR[ 64 ][ 210 ],
   alphaCSR[ 64 ][ 211 ],
   alphaCSR[ 64 ][ 212 ],
   alphaCSR[ 64 ][ 213 ],
   alphaCSR[ 64 ][ 214 ],
   alphaCSR[ 64 ][ 215 ],
   alphaCSR[ 64 ][ 216 ],
   alphaCSR[ 64 ][ 217 ],
   alphaCSR[ 64 ][ 218 ],
   alphaCSR[ 64 ][ 219 ],
   alphaCSR[ 64 ][ 220 ],
   alphaCSR[ 64 ][ 221 ],
   alphaCSR[ 64 ][ 222 ],
   alphaCSR[ 64 ][ 223 ],
   alphaCSR[ 64 ][ 224 ],
   alphaCSR[ 64 ][ 225 ],
   alphaCSR[ 64 ][ 226 ],
   alphaCSR[ 64 ][ 227 ],
   alphaCSR[ 64 ][ 228 ],
   alphaCSR[ 64 ][ 229 ],
   alphaCSR[ 64 ][ 230 ],
   alphaCSR[ 64 ][ 231 ],
   alphaCSR[ 64 ][ 232 ],
   alphaCSR[ 64 ][ 233 ],
   alphaCSR[ 64 ][ 234 ],
   alphaCSR[ 64 ][ 235 ],
   alphaCSR[ 64 ][ 236 ],
   alphaCSR[ 64 ][ 237 ],
   alphaCSR[ 64 ][ 238 ],
   alphaCSR[ 64 ][ 239 ],
   alphaCSR[ 64 ][ 240 ],
   alphaCSR[ 64 ][ 241 ],
   alphaCSR[ 64 ][ 242 ],
   alphaCSR[ 64 ][ 243 ],
   alphaCSR[ 64 ][ 244 ],
   alphaCSR[ 64 ][ 245 ],
   alphaCSR[ 64 ][ 246 ],
   alphaCSR[ 64 ][ 247 ],
   alphaCSR[ 64 ][ 248 ],
   alphaCSR[ 64 ][ 249 ],
   alphaCSR[ 64 ][ 250 ],
   alphaCSR[ 64 ][ 251 ],
   alphaCSR[ 64 ][ 252 ],
   alphaCSR[ 64 ][ 253 ],
   alphaCSR[ 64 ][ 254 ],
   alphaCSR[ 64 ][ 255 ],
   alphaCSR[ 64 ][ 256 ],
   alphaCSR[ 64 ][ 257 ],
   alphaCSR[ 64 ][ 258 ],
   alphaCSR[ 64 ][ 259 ],
   alphaCSR[ 64 ][ 260 ],
   alphaCSR[ 64 ][ 261 ],
   alphaCSR[ 64 ][ 262 ],
   alphaCSR[ 64 ][ 263 ],
   alphaCSR[ 64 ][ 264 ],
   alphaCSR[ 64 ][ 265 ],
   alphaCSR[ 64 ][ 266 ],
   alphaCSR[ 64 ][ 267 ],
   alphaCSR[ 64 ][ 268 ],
   alphaCSR[ 64 ][ 269 ],
   alphaCSR[ 64 ][ 270 ],
   alphaCSR[ 64 ][ 271 ],
   alphaCSR[ 64 ][ 272 ],
   alphaCSR[ 64 ][ 273 ],
   alphaCSR[ 64 ][ 274 ],
   alphaCSR[ 64 ][ 275 ],
   alphaCSR[ 64 ][ 276 ],
   alphaCSR[ 64 ][ 277 ],
   alphaCSR[ 64 ][ 278 ],
   alphaCSR[ 64 ][ 279 ],
   alphaCSR[ 64 ][ 280 ],
   alphaCSR[ 64 ][ 281 ],
   alphaCSR[ 64 ][ 282 ],
   alphaCSR[ 64 ][ 283 ],
   alphaCSR[ 64 ][ 284 ],
   alphaCSR[ 64 ][ 285 ],
   alphaCSR[ 64 ][ 286 ],
   alphaCSR[ 64 ][ 287 ],
   alphaCSR[ 64 ][ 288 ],
   alphaCSR[ 64 ][ 289 ],
   alphaCSR[ 64 ][ 290 ],
   alphaCSR[ 64 ][ 291 ],
   alphaCSR[ 64 ][ 292 ],
   alphaCSR[ 64 ][ 293 ],
   alphaCSR[ 64 ][ 294 ],
   alphaCSR[ 64 ][ 295 ],
   alphaCSR[ 64 ][ 296 ],
   alphaCSR[ 64 ][ 297 ],
   alphaCSR[ 64 ][ 298 ],
   alphaCSR[ 64 ][ 299 ],
   alphaCSR[ 64 ][ 300 ],
   alphaCSR[ 64 ][ 301 ],
   alphaCSR[ 64 ][ 302 ],
   alphaCSR[ 64 ][ 303 ],
   alphaCSR[ 64 ][ 304 ],
   alphaCSR[ 64 ][ 305 ],
   alphaCSR[ 64 ][ 306 ],
   alphaCSR[ 64 ][ 307 ],
   alphaCSR[ 64 ][ 308 ],
   alphaCSR[ 64 ][ 309 ],
   alphaCSR[ 64 ][ 310 ],
   alphaCSR[ 64 ][ 311 ],
   alphaCSR[ 64 ][ 312 ],
   alphaCSR[ 64 ][ 313 ],
   alphaCSR[ 64 ][ 314 ],
   alphaCSR[ 64 ][ 315 ],
   alphaCSR[ 64 ][ 316 ],
   alphaCSR[ 64 ][ 317 ],
   alphaCSR[ 64 ][ 318 ],
   alphaCSR[ 64 ][ 319 ],
   alphaCSR[ 64 ][ 320 ],
   alphaCSR[ 64 ][ 321 ],
   alphaCSR[ 64 ][ 322 ],
   alphaCSR[ 64 ][ 323 ],
   alphaCSR[ 64 ][ 324 ],
   alphaCSR[ 64 ][ 325 ],
   alphaCSR[ 64 ][ 326 ],
   alphaCSR[ 64 ][ 327 ],
   alphaCSR[ 64 ][ 328 ],
   alphaCSR[ 64 ][ 329 ],
   alphaCSR[ 64 ][ 330 ],
   alphaCSR[ 64 ][ 331 ],
   alphaCSR[ 64 ][ 332 ],
   alphaCSR[ 64 ][ 333 ],
   alphaCSR[ 64 ][ 334 ],
   alphaCSR[ 64 ][ 335 ],
   alphaCSR[ 64 ][ 336 ],
   alphaCSR[ 64 ][ 337 ],
   alphaCSR[ 64 ][ 338 ],
   alphaCSR[ 64 ][ 339 ],
   alphaCSR[ 64 ][ 340 ],
   alphaCSR[ 64 ][ 341 ],
   alphaCSR[ 64 ][ 342 ],
   alphaCSR[ 64 ][ 343 ],
   alphaCSR[ 64 ][ 344 ],
   alphaCSR[ 64 ][ 345 ],
   alphaCSR[ 64 ][ 346 ],
   alphaCSR[ 64 ][ 347 ],
   alphaCSR[ 64 ][ 348 ],
   alphaCSR[ 64 ][ 349 ],
   alphaCSR[ 64 ][ 350 ],
   alphaCSR[ 64 ][ 351 ],
   alphaCSR[ 64 ][ 352 ],
   alphaCSR[ 64 ][ 353 ],
   alphaCSR[ 64 ][ 354 ],
   alphaCSR[ 64 ][ 355 ],
   alphaCSR[ 64 ][ 356 ],
   alphaCSR[ 64 ][ 357 ],
   alphaCSR[ 64 ][ 358 ],
   alphaCSR[ 64 ][ 359 ],
   alphaCSR[ 64 ][ 360 ],
   alphaCSR[ 64 ][ 361 ],
   alphaCSR[ 64 ][ 362 ],
   alphaCSR[ 64 ][ 363 ],
   alphaCSR[ 64 ][ 364 ],
   alphaCSR[ 64 ][ 365 ],
   alphaCSR[ 64 ][ 366 ],
   alphaCSR[ 64 ][ 367 ],
   alphaCSR[ 64 ][ 368 ],
   alphaCSR[ 64 ][ 369 ],
   alphaCSR[ 64 ][ 370 ],
   alphaCSR[ 64 ][ 371 ],
   alphaCSR[ 64 ][ 372 ],
   alphaCSR[ 64 ][ 373 ],
   alphaCSR[ 64 ][ 374 ],
   alphaCSR[ 64 ][ 375 ],
   alphaCSR[ 64 ][ 376 ],
   alphaCSR[ 64 ][ 377 ],
   alphaCSR[ 64 ][ 378 ],
   alphaCSR[ 64 ][ 379 ],
   alphaCSR[ 64 ][ 380 ],
   alphaCSR[ 64 ][ 381 ],
   alphaCSR[ 64 ][ 382 ],
   alphaCSR[ 64 ][ 383 ],
   alphaCSR[ 65 ][ 0 ],
   alphaCSR[ 65 ][ 1 ],
   alphaCSR[ 65 ][ 2 ],
   alphaCSR[ 65 ][ 3 ],
   alphaCSR[ 65 ][ 4 ],
   alphaCSR[ 65 ][ 5 ],
   alphaCSR[ 65 ][ 6 ],
   alphaCSR[ 65 ][ 7 ],
   alphaCSR[ 65 ][ 8 ],
   alphaCSR[ 65 ][ 9 ],
   alphaCSR[ 65 ][ 10 ],
   alphaCSR[ 65 ][ 11 ],
   alphaCSR[ 65 ][ 12 ],
   alphaCSR[ 65 ][ 13 ],
   alphaCSR[ 65 ][ 14 ],
   alphaCSR[ 65 ][ 15 ],
   alphaCSR[ 65 ][ 16 ],
   alphaCSR[ 65 ][ 17 ],
   alphaCSR[ 65 ][ 18 ],
   alphaCSR[ 65 ][ 19 ],
   alphaCSR[ 65 ][ 20 ],
   alphaCSR[ 65 ][ 21 ],
   alphaCSR[ 65 ][ 22 ],
   alphaCSR[ 65 ][ 23 ],
   alphaCSR[ 65 ][ 24 ],
   alphaCSR[ 65 ][ 25 ],
   alphaCSR[ 65 ][ 26 ],
   alphaCSR[ 65 ][ 27 ],
   alphaCSR[ 65 ][ 28 ],
   alphaCSR[ 65 ][ 29 ],
   alphaCSR[ 65 ][ 30 ],
   alphaCSR[ 65 ][ 31 ],
   alphaCSR[ 65 ][ 32 ],
   alphaCSR[ 65 ][ 33 ],
   alphaCSR[ 65 ][ 34 ],
   alphaCSR[ 65 ][ 35 ],
   alphaCSR[ 65 ][ 36 ],
   alphaCSR[ 65 ][ 37 ],
   alphaCSR[ 65 ][ 38 ],
   alphaCSR[ 65 ][ 39 ],
   alphaCSR[ 65 ][ 40 ],
   alphaCSR[ 65 ][ 41 ],
   alphaCSR[ 65 ][ 42 ],
   alphaCSR[ 65 ][ 43 ],
   alphaCSR[ 65 ][ 44 ],
   alphaCSR[ 65 ][ 45 ],
   alphaCSR[ 65 ][ 46 ],
   alphaCSR[ 65 ][ 47 ],
   alphaCSR[ 65 ][ 48 ],
   alphaCSR[ 65 ][ 49 ],
   alphaCSR[ 65 ][ 50 ],
   alphaCSR[ 65 ][ 51 ],
   alphaCSR[ 65 ][ 52 ],
   alphaCSR[ 65 ][ 53 ],
   alphaCSR[ 65 ][ 54 ],
   alphaCSR[ 65 ][ 55 ],
   alphaCSR[ 65 ][ 56 ],
   alphaCSR[ 65 ][ 57 ],
   alphaCSR[ 65 ][ 58 ],
   alphaCSR[ 65 ][ 59 ],
   alphaCSR[ 65 ][ 60 ],
   alphaCSR[ 65 ][ 61 ],
   alphaCSR[ 65 ][ 62 ],
   alphaCSR[ 65 ][ 63 ],
   alphaCSR[ 65 ][ 64 ],
   alphaCSR[ 65 ][ 65 ],
   alphaCSR[ 65 ][ 66 ],
   alphaCSR[ 65 ][ 67 ],
   alphaCSR[ 65 ][ 68 ],
   alphaCSR[ 65 ][ 69 ],
   alphaCSR[ 65 ][ 70 ],
   alphaCSR[ 65 ][ 71 ],
   alphaCSR[ 65 ][ 72 ],
   alphaCSR[ 65 ][ 73 ],
   alphaCSR[ 65 ][ 74 ],
   alphaCSR[ 65 ][ 75 ],
   alphaCSR[ 65 ][ 76 ],
   alphaCSR[ 65 ][ 77 ],
   alphaCSR[ 65 ][ 78 ],
   alphaCSR[ 65 ][ 79 ],
   alphaCSR[ 65 ][ 80 ],
   alphaCSR[ 65 ][ 81 ],
   alphaCSR[ 65 ][ 82 ],
   alphaCSR[ 65 ][ 83 ],
   alphaCSR[ 65 ][ 84 ],
   alphaCSR[ 65 ][ 85 ],
   alphaCSR[ 65 ][ 86 ],
   alphaCSR[ 65 ][ 87 ],
   alphaCSR[ 65 ][ 88 ],
   alphaCSR[ 65 ][ 89 ],
   alphaCSR[ 65 ][ 90 ],
   alphaCSR[ 65 ][ 91 ],
   alphaCSR[ 65 ][ 92 ],
   alphaCSR[ 65 ][ 93 ],
   alphaCSR[ 65 ][ 94 ],
   alphaCSR[ 65 ][ 95 ],
   alphaCSR[ 65 ][ 96 ],
   alphaCSR[ 65 ][ 97 ],
   alphaCSR[ 65 ][ 98 ],
   alphaCSR[ 65 ][ 99 ],
   alphaCSR[ 65 ][ 100 ],
   alphaCSR[ 65 ][ 101 ],
   alphaCSR[ 65 ][ 102 ],
   alphaCSR[ 65 ][ 103 ],
   alphaCSR[ 65 ][ 104 ],
   alphaCSR[ 65 ][ 105 ],
   alphaCSR[ 65 ][ 106 ],
   alphaCSR[ 65 ][ 107 ],
   alphaCSR[ 65 ][ 108 ],
   alphaCSR[ 65 ][ 109 ],
   alphaCSR[ 65 ][ 110 ],
   alphaCSR[ 65 ][ 111 ],
   alphaCSR[ 65 ][ 112 ],
   alphaCSR[ 65 ][ 113 ],
   alphaCSR[ 65 ][ 114 ],
   alphaCSR[ 65 ][ 115 ],
   alphaCSR[ 65 ][ 116 ],
   alphaCSR[ 65 ][ 117 ],
   alphaCSR[ 65 ][ 118 ],
   alphaCSR[ 65 ][ 119 ],
   alphaCSR[ 65 ][ 120 ],
   alphaCSR[ 65 ][ 121 ],
   alphaCSR[ 65 ][ 122 ],
   alphaCSR[ 65 ][ 123 ],
   alphaCSR[ 65 ][ 124 ],
   alphaCSR[ 65 ][ 125 ],
   alphaCSR[ 65 ][ 126 ],
   alphaCSR[ 65 ][ 127 ],
   alphaCSR[ 65 ][ 128 ],
   alphaCSR[ 65 ][ 129 ],
   alphaCSR[ 65 ][ 130 ],
   alphaCSR[ 65 ][ 131 ],
   alphaCSR[ 65 ][ 132 ],
   alphaCSR[ 65 ][ 133 ],
   alphaCSR[ 65 ][ 134 ],
   alphaCSR[ 65 ][ 135 ],
   alphaCSR[ 65 ][ 136 ],
   alphaCSR[ 65 ][ 137 ],
   alphaCSR[ 65 ][ 138 ],
   alphaCSR[ 65 ][ 139 ],
   alphaCSR[ 65 ][ 140 ],
   alphaCSR[ 65 ][ 141 ],
   alphaCSR[ 65 ][ 142 ],
   alphaCSR[ 65 ][ 143 ],
   alphaCSR[ 65 ][ 144 ],
   alphaCSR[ 65 ][ 145 ],
   alphaCSR[ 65 ][ 146 ],
   alphaCSR[ 65 ][ 147 ],
   alphaCSR[ 65 ][ 148 ],
   alphaCSR[ 65 ][ 149 ],
   alphaCSR[ 65 ][ 150 ],
   alphaCSR[ 65 ][ 151 ],
   alphaCSR[ 65 ][ 152 ],
   alphaCSR[ 65 ][ 153 ],
   alphaCSR[ 65 ][ 154 ],
   alphaCSR[ 65 ][ 155 ],
   alphaCSR[ 65 ][ 156 ],
   alphaCSR[ 65 ][ 157 ],
   alphaCSR[ 65 ][ 158 ],
   alphaCSR[ 65 ][ 159 ],
   alphaCSR[ 65 ][ 160 ],
   alphaCSR[ 65 ][ 161 ],
   alphaCSR[ 65 ][ 162 ],
   alphaCSR[ 65 ][ 163 ],
   alphaCSR[ 65 ][ 164 ],
   alphaCSR[ 65 ][ 165 ],
   alphaCSR[ 65 ][ 166 ],
   alphaCSR[ 65 ][ 167 ],
   alphaCSR[ 65 ][ 168 ],
   alphaCSR[ 65 ][ 169 ],
   alphaCSR[ 65 ][ 170 ],
   alphaCSR[ 65 ][ 171 ],
   alphaCSR[ 65 ][ 172 ],
   alphaCSR[ 65 ][ 173 ],
   alphaCSR[ 65 ][ 174 ],
   alphaCSR[ 65 ][ 175 ],
   alphaCSR[ 65 ][ 176 ],
   alphaCSR[ 65 ][ 177 ],
   alphaCSR[ 65 ][ 178 ],
   alphaCSR[ 65 ][ 179 ],
   alphaCSR[ 65 ][ 180 ],
   alphaCSR[ 65 ][ 181 ],
   alphaCSR[ 65 ][ 182 ],
   alphaCSR[ 65 ][ 183 ],
   alphaCSR[ 65 ][ 184 ],
   alphaCSR[ 65 ][ 185 ],
   alphaCSR[ 65 ][ 186 ],
   alphaCSR[ 65 ][ 187 ],
   alphaCSR[ 65 ][ 188 ],
   alphaCSR[ 65 ][ 189 ],
   alphaCSR[ 65 ][ 190 ],
   alphaCSR[ 65 ][ 191 ],
   alphaCSR[ 65 ][ 192 ],
   alphaCSR[ 65 ][ 193 ],
   alphaCSR[ 65 ][ 194 ],
   alphaCSR[ 65 ][ 195 ],
   alphaCSR[ 65 ][ 196 ],
   alphaCSR[ 65 ][ 197 ],
   alphaCSR[ 65 ][ 198 ],
   alphaCSR[ 65 ][ 199 ],
   alphaCSR[ 65 ][ 200 ],
   alphaCSR[ 65 ][ 201 ],
   alphaCSR[ 65 ][ 202 ],
   alphaCSR[ 65 ][ 203 ],
   alphaCSR[ 65 ][ 204 ],
   alphaCSR[ 65 ][ 205 ],
   alphaCSR[ 65 ][ 206 ],
   alphaCSR[ 65 ][ 207 ],
   alphaCSR[ 65 ][ 208 ],
   alphaCSR[ 65 ][ 209 ],
   alphaCSR[ 65 ][ 210 ],
   alphaCSR[ 65 ][ 211 ],
   alphaCSR[ 65 ][ 212 ],
   alphaCSR[ 65 ][ 213 ],
   alphaCSR[ 65 ][ 214 ],
   alphaCSR[ 65 ][ 215 ],
   alphaCSR[ 65 ][ 216 ],
   alphaCSR[ 65 ][ 217 ],
   alphaCSR[ 65 ][ 218 ],
   alphaCSR[ 65 ][ 219 ],
   alphaCSR[ 65 ][ 220 ],
   alphaCSR[ 65 ][ 221 ],
   alphaCSR[ 65 ][ 222 ],
   alphaCSR[ 65 ][ 223 ],
   alphaCSR[ 65 ][ 224 ],
   alphaCSR[ 65 ][ 225 ],
   alphaCSR[ 65 ][ 226 ],
   alphaCSR[ 65 ][ 227 ],
   alphaCSR[ 65 ][ 228 ],
   alphaCSR[ 65 ][ 229 ],
   alphaCSR[ 65 ][ 230 ],
   alphaCSR[ 65 ][ 231 ],
   alphaCSR[ 65 ][ 232 ],
   alphaCSR[ 65 ][ 233 ],
   alphaCSR[ 65 ][ 234 ],
   alphaCSR[ 65 ][ 235 ],
   alphaCSR[ 65 ][ 236 ],
   alphaCSR[ 65 ][ 237 ],
   alphaCSR[ 65 ][ 238 ],
   alphaCSR[ 65 ][ 239 ],
   alphaCSR[ 65 ][ 240 ],
   alphaCSR[ 65 ][ 241 ],
   alphaCSR[ 65 ][ 242 ],
   alphaCSR[ 65 ][ 243 ],
   alphaCSR[ 65 ][ 244 ],
   alphaCSR[ 65 ][ 245 ],
   alphaCSR[ 65 ][ 246 ],
   alphaCSR[ 65 ][ 247 ],
   alphaCSR[ 65 ][ 248 ],
   alphaCSR[ 65 ][ 249 ],
   alphaCSR[ 65 ][ 250 ],
   alphaCSR[ 65 ][ 251 ],
   alphaCSR[ 65 ][ 252 ],
   alphaCSR[ 65 ][ 253 ],
   alphaCSR[ 65 ][ 254 ],
   alphaCSR[ 65 ][ 255 ],
   alphaCSR[ 65 ][ 256 ],
   alphaCSR[ 65 ][ 257 ],
   alphaCSR[ 65 ][ 258 ],
   alphaCSR[ 65 ][ 259 ],
   alphaCSR[ 65 ][ 260 ],
   alphaCSR[ 65 ][ 261 ],
   alphaCSR[ 65 ][ 262 ],
   alphaCSR[ 65 ][ 263 ],
   alphaCSR[ 65 ][ 264 ],
   alphaCSR[ 65 ][ 265 ],
   alphaCSR[ 65 ][ 266 ],
   alphaCSR[ 65 ][ 267 ],
   alphaCSR[ 65 ][ 268 ],
   alphaCSR[ 65 ][ 269 ],
   alphaCSR[ 65 ][ 270 ],
   alphaCSR[ 65 ][ 271 ],
   alphaCSR[ 65 ][ 272 ],
   alphaCSR[ 65 ][ 273 ],
   alphaCSR[ 65 ][ 274 ],
   alphaCSR[ 65 ][ 275 ],
   alphaCSR[ 65 ][ 276 ],
   alphaCSR[ 65 ][ 277 ],
   alphaCSR[ 65 ][ 278 ],
   alphaCSR[ 65 ][ 279 ],
   alphaCSR[ 65 ][ 280 ],
   alphaCSR[ 65 ][ 281 ],
   alphaCSR[ 65 ][ 282 ],
   alphaCSR[ 65 ][ 283 ],
   alphaCSR[ 65 ][ 284 ],
   alphaCSR[ 65 ][ 285 ],
   alphaCSR[ 65 ][ 286 ],
   alphaCSR[ 65 ][ 287 ],
   alphaCSR[ 65 ][ 288 ],
   alphaCSR[ 65 ][ 289 ],
   alphaCSR[ 65 ][ 290 ],
   alphaCSR[ 65 ][ 291 ],
   alphaCSR[ 65 ][ 292 ],
   alphaCSR[ 65 ][ 293 ],
   alphaCSR[ 65 ][ 294 ],
   alphaCSR[ 65 ][ 295 ],
   alphaCSR[ 65 ][ 296 ],
   alphaCSR[ 65 ][ 297 ],
   alphaCSR[ 65 ][ 298 ],
   alphaCSR[ 65 ][ 299 ],
   alphaCSR[ 65 ][ 300 ],
   alphaCSR[ 65 ][ 301 ],
   alphaCSR[ 65 ][ 302 ],
   alphaCSR[ 65 ][ 303 ],
   alphaCSR[ 65 ][ 304 ],
   alphaCSR[ 65 ][ 305 ],
   alphaCSR[ 65 ][ 306 ],
   alphaCSR[ 65 ][ 307 ],
   alphaCSR[ 65 ][ 308 ],
   alphaCSR[ 65 ][ 309 ],
   alphaCSR[ 65 ][ 310 ],
   alphaCSR[ 65 ][ 311 ],
   alphaCSR[ 65 ][ 312 ],
   alphaCSR[ 65 ][ 313 ],
   alphaCSR[ 65 ][ 314 ],
   alphaCSR[ 65 ][ 315 ],
   alphaCSR[ 65 ][ 316 ],
   alphaCSR[ 65 ][ 317 ],
   alphaCSR[ 65 ][ 318 ],
   alphaCSR[ 65 ][ 319 ],
   alphaCSR[ 65 ][ 320 ],
   alphaCSR[ 65 ][ 321 ],
   alphaCSR[ 65 ][ 322 ],
   alphaCSR[ 65 ][ 323 ],
   alphaCSR[ 65 ][ 324 ],
   alphaCSR[ 65 ][ 325 ],
   alphaCSR[ 65 ][ 326 ],
   alphaCSR[ 65 ][ 327 ],
   alphaCSR[ 65 ][ 328 ],
   alphaCSR[ 65 ][ 329 ],
   alphaCSR[ 65 ][ 330 ],
   alphaCSR[ 65 ][ 331 ],
   alphaCSR[ 65 ][ 332 ],
   alphaCSR[ 65 ][ 333 ],
   alphaCSR[ 65 ][ 334 ],
   alphaCSR[ 65 ][ 335 ],
   alphaCSR[ 65 ][ 336 ],
   alphaCSR[ 65 ][ 337 ],
   alphaCSR[ 65 ][ 338 ],
   alphaCSR[ 65 ][ 339 ],
   alphaCSR[ 65 ][ 340 ],
   alphaCSR[ 65 ][ 341 ],
   alphaCSR[ 65 ][ 342 ],
   alphaCSR[ 65 ][ 343 ],
   alphaCSR[ 65 ][ 344 ],
   alphaCSR[ 65 ][ 345 ],
   alphaCSR[ 65 ][ 346 ],
   alphaCSR[ 65 ][ 347 ],
   alphaCSR[ 65 ][ 348 ],
   alphaCSR[ 65 ][ 349 ],
   alphaCSR[ 65 ][ 350 ],
   alphaCSR[ 65 ][ 351 ],
   alphaCSR[ 65 ][ 352 ],
   alphaCSR[ 65 ][ 353 ],
   alphaCSR[ 65 ][ 354 ],
   alphaCSR[ 65 ][ 355 ],
   alphaCSR[ 65 ][ 356 ],
   alphaCSR[ 65 ][ 357 ],
   alphaCSR[ 65 ][ 358 ],
   alphaCSR[ 65 ][ 359 ],
   alphaCSR[ 65 ][ 360 ],
   alphaCSR[ 65 ][ 361 ],
   alphaCSR[ 65 ][ 362 ],
   alphaCSR[ 65 ][ 363 ],
   alphaCSR[ 65 ][ 364 ],
   alphaCSR[ 65 ][ 365 ],
   alphaCSR[ 65 ][ 366 ],
   alphaCSR[ 65 ][ 367 ],
   alphaCSR[ 65 ][ 368 ],
   alphaCSR[ 65 ][ 369 ],
   alphaCSR[ 65 ][ 370 ],
   alphaCSR[ 65 ][ 371 ],
   alphaCSR[ 65 ][ 372 ],
   alphaCSR[ 65 ][ 373 ],
   alphaCSR[ 65 ][ 374 ],
   alphaCSR[ 65 ][ 375 ],
   alphaCSR[ 65 ][ 376 ],
   alphaCSR[ 65 ][ 377 ],
   alphaCSR[ 65 ][ 378 ],
   alphaCSR[ 65 ][ 379 ],
   alphaCSR[ 65 ][ 380 ],
   alphaCSR[ 65 ][ 381 ],
   alphaCSR[ 65 ][ 382 ],
   alphaCSR[ 65 ][ 383 ],
   alphaCSR[ 66 ][ 0 ],
   alphaCSR[ 66 ][ 1 ],
   alphaCSR[ 66 ][ 2 ],
   alphaCSR[ 66 ][ 3 ],
   alphaCSR[ 66 ][ 4 ],
   alphaCSR[ 66 ][ 5 ],
   alphaCSR[ 66 ][ 6 ],
   alphaCSR[ 66 ][ 7 ],
   alphaCSR[ 66 ][ 8 ],
   alphaCSR[ 66 ][ 9 ],
   alphaCSR[ 66 ][ 10 ],
   alphaCSR[ 66 ][ 11 ],
   alphaCSR[ 66 ][ 12 ],
   alphaCSR[ 66 ][ 13 ],
   alphaCSR[ 66 ][ 14 ],
   alphaCSR[ 66 ][ 15 ],
   alphaCSR[ 66 ][ 16 ],
   alphaCSR[ 66 ][ 17 ],
   alphaCSR[ 66 ][ 18 ],
   alphaCSR[ 66 ][ 19 ],
   alphaCSR[ 66 ][ 20 ],
   alphaCSR[ 66 ][ 21 ],
   alphaCSR[ 66 ][ 22 ],
   alphaCSR[ 66 ][ 23 ],
   alphaCSR[ 66 ][ 24 ],
   alphaCSR[ 66 ][ 25 ],
   alphaCSR[ 66 ][ 26 ],
   alphaCSR[ 66 ][ 27 ],
   alphaCSR[ 66 ][ 28 ],
   alphaCSR[ 66 ][ 29 ],
   alphaCSR[ 66 ][ 30 ],
   alphaCSR[ 66 ][ 31 ],
   alphaCSR[ 66 ][ 32 ],
   alphaCSR[ 66 ][ 33 ],
   alphaCSR[ 66 ][ 34 ],
   alphaCSR[ 66 ][ 35 ],
   alphaCSR[ 66 ][ 36 ],
   alphaCSR[ 66 ][ 37 ],
   alphaCSR[ 66 ][ 38 ],
   alphaCSR[ 66 ][ 39 ],
   alphaCSR[ 66 ][ 40 ],
   alphaCSR[ 66 ][ 41 ],
   alphaCSR[ 66 ][ 42 ],
   alphaCSR[ 66 ][ 43 ],
   alphaCSR[ 66 ][ 44 ],
   alphaCSR[ 66 ][ 45 ],
   alphaCSR[ 66 ][ 46 ],
   alphaCSR[ 66 ][ 47 ],
   alphaCSR[ 66 ][ 48 ],
   alphaCSR[ 66 ][ 49 ],
   alphaCSR[ 66 ][ 50 ],
   alphaCSR[ 66 ][ 51 ],
   alphaCSR[ 66 ][ 52 ],
   alphaCSR[ 66 ][ 53 ],
   alphaCSR[ 66 ][ 54 ],
   alphaCSR[ 66 ][ 55 ],
   alphaCSR[ 66 ][ 56 ],
   alphaCSR[ 66 ][ 57 ],
   alphaCSR[ 66 ][ 58 ],
   alphaCSR[ 66 ][ 59 ],
   alphaCSR[ 66 ][ 60 ],
   alphaCSR[ 66 ][ 61 ],
   alphaCSR[ 66 ][ 62 ],
   alphaCSR[ 66 ][ 63 ],
   alphaCSR[ 66 ][ 64 ],
   alphaCSR[ 66 ][ 65 ],
   alphaCSR[ 66 ][ 66 ],
   alphaCSR[ 66 ][ 67 ],
   alphaCSR[ 66 ][ 68 ],
   alphaCSR[ 66 ][ 69 ],
   alphaCSR[ 66 ][ 70 ],
   alphaCSR[ 66 ][ 71 ],
   alphaCSR[ 66 ][ 72 ],
   alphaCSR[ 66 ][ 73 ],
   alphaCSR[ 66 ][ 74 ],
   alphaCSR[ 66 ][ 75 ],
   alphaCSR[ 66 ][ 76 ],
   alphaCSR[ 66 ][ 77 ],
   alphaCSR[ 66 ][ 78 ],
   alphaCSR[ 66 ][ 79 ],
   alphaCSR[ 66 ][ 80 ],
   alphaCSR[ 66 ][ 81 ],
   alphaCSR[ 66 ][ 82 ],
   alphaCSR[ 66 ][ 83 ],
   alphaCSR[ 66 ][ 84 ],
   alphaCSR[ 66 ][ 85 ],
   alphaCSR[ 66 ][ 86 ],
   alphaCSR[ 66 ][ 87 ],
   alphaCSR[ 66 ][ 88 ],
   alphaCSR[ 66 ][ 89 ],
   alphaCSR[ 66 ][ 90 ],
   alphaCSR[ 66 ][ 91 ],
   alphaCSR[ 66 ][ 92 ],
   alphaCSR[ 66 ][ 93 ],
   alphaCSR[ 66 ][ 94 ],
   alphaCSR[ 66 ][ 95 ],
   alphaCSR[ 66 ][ 96 ],
   alphaCSR[ 66 ][ 97 ],
   alphaCSR[ 66 ][ 98 ],
   alphaCSR[ 66 ][ 99 ],
   alphaCSR[ 66 ][ 100 ],
   alphaCSR[ 66 ][ 101 ],
   alphaCSR[ 66 ][ 102 ],
   alphaCSR[ 66 ][ 103 ],
   alphaCSR[ 66 ][ 104 ],
   alphaCSR[ 66 ][ 105 ],
   alphaCSR[ 66 ][ 106 ],
   alphaCSR[ 66 ][ 107 ],
   alphaCSR[ 66 ][ 108 ],
   alphaCSR[ 66 ][ 109 ],
   alphaCSR[ 66 ][ 110 ],
   alphaCSR[ 66 ][ 111 ],
   alphaCSR[ 66 ][ 112 ],
   alphaCSR[ 66 ][ 113 ],
   alphaCSR[ 66 ][ 114 ],
   alphaCSR[ 66 ][ 115 ],
   alphaCSR[ 66 ][ 116 ],
   alphaCSR[ 66 ][ 117 ],
   alphaCSR[ 66 ][ 118 ],
   alphaCSR[ 66 ][ 119 ],
   alphaCSR[ 66 ][ 120 ],
   alphaCSR[ 66 ][ 121 ],
   alphaCSR[ 66 ][ 122 ],
   alphaCSR[ 66 ][ 123 ],
   alphaCSR[ 66 ][ 124 ],
   alphaCSR[ 66 ][ 125 ],
   alphaCSR[ 66 ][ 126 ],
   alphaCSR[ 66 ][ 127 ],
   alphaCSR[ 66 ][ 128 ],
   alphaCSR[ 66 ][ 129 ],
   alphaCSR[ 66 ][ 130 ],
   alphaCSR[ 66 ][ 131 ],
   alphaCSR[ 66 ][ 132 ],
   alphaCSR[ 66 ][ 133 ],
   alphaCSR[ 66 ][ 134 ],
   alphaCSR[ 66 ][ 135 ],
   alphaCSR[ 66 ][ 136 ],
   alphaCSR[ 66 ][ 137 ],
   alphaCSR[ 66 ][ 138 ],
   alphaCSR[ 66 ][ 139 ],
   alphaCSR[ 66 ][ 140 ],
   alphaCSR[ 66 ][ 141 ],
   alphaCSR[ 66 ][ 142 ],
   alphaCSR[ 66 ][ 143 ],
   alphaCSR[ 66 ][ 144 ],
   alphaCSR[ 66 ][ 145 ],
   alphaCSR[ 66 ][ 146 ],
   alphaCSR[ 66 ][ 147 ],
   alphaCSR[ 66 ][ 148 ],
   alphaCSR[ 66 ][ 149 ],
   alphaCSR[ 66 ][ 150 ],
   alphaCSR[ 66 ][ 151 ],
   alphaCSR[ 66 ][ 152 ],
   alphaCSR[ 66 ][ 153 ],
   alphaCSR[ 66 ][ 154 ],
   alphaCSR[ 66 ][ 155 ],
   alphaCSR[ 66 ][ 156 ],
   alphaCSR[ 66 ][ 157 ],
   alphaCSR[ 66 ][ 158 ],
   alphaCSR[ 66 ][ 159 ],
   alphaCSR[ 66 ][ 160 ],
   alphaCSR[ 66 ][ 161 ],
   alphaCSR[ 66 ][ 162 ],
   alphaCSR[ 66 ][ 163 ],
   alphaCSR[ 66 ][ 164 ],
   alphaCSR[ 66 ][ 165 ],
   alphaCSR[ 66 ][ 166 ],
   alphaCSR[ 66 ][ 167 ],
   alphaCSR[ 66 ][ 168 ],
   alphaCSR[ 66 ][ 169 ],
   alphaCSR[ 66 ][ 170 ],
   alphaCSR[ 66 ][ 171 ],
   alphaCSR[ 66 ][ 172 ],
   alphaCSR[ 66 ][ 173 ],
   alphaCSR[ 66 ][ 174 ],
   alphaCSR[ 66 ][ 175 ],
   alphaCSR[ 66 ][ 176 ],
   alphaCSR[ 66 ][ 177 ],
   alphaCSR[ 66 ][ 178 ],
   alphaCSR[ 66 ][ 179 ],
   alphaCSR[ 66 ][ 180 ],
   alphaCSR[ 66 ][ 181 ],
   alphaCSR[ 66 ][ 182 ],
   alphaCSR[ 66 ][ 183 ],
   alphaCSR[ 66 ][ 184 ],
   alphaCSR[ 66 ][ 185 ],
   alphaCSR[ 66 ][ 186 ],
   alphaCSR[ 66 ][ 187 ],
   alphaCSR[ 66 ][ 188 ],
   alphaCSR[ 66 ][ 189 ],
   alphaCSR[ 66 ][ 190 ],
   alphaCSR[ 66 ][ 191 ],
   alphaCSR[ 66 ][ 192 ],
   alphaCSR[ 66 ][ 193 ],
   alphaCSR[ 66 ][ 194 ],
   alphaCSR[ 66 ][ 195 ],
   alphaCSR[ 66 ][ 196 ],
   alphaCSR[ 66 ][ 197 ],
   alphaCSR[ 66 ][ 198 ],
   alphaCSR[ 66 ][ 199 ],
   alphaCSR[ 66 ][ 200 ],
   alphaCSR[ 66 ][ 201 ],
   alphaCSR[ 66 ][ 202 ],
   alphaCSR[ 66 ][ 203 ],
   alphaCSR[ 66 ][ 204 ],
   alphaCSR[ 66 ][ 205 ],
   alphaCSR[ 66 ][ 206 ],
   alphaCSR[ 66 ][ 207 ],
   alphaCSR[ 66 ][ 208 ],
   alphaCSR[ 66 ][ 209 ],
   alphaCSR[ 66 ][ 210 ],
   alphaCSR[ 66 ][ 211 ],
   alphaCSR[ 66 ][ 212 ],
   alphaCSR[ 66 ][ 213 ],
   alphaCSR[ 66 ][ 214 ],
   alphaCSR[ 66 ][ 215 ],
   alphaCSR[ 66 ][ 216 ],
   alphaCSR[ 66 ][ 217 ],
   alphaCSR[ 66 ][ 218 ],
   alphaCSR[ 66 ][ 219 ],
   alphaCSR[ 66 ][ 220 ],
   alphaCSR[ 66 ][ 221 ],
   alphaCSR[ 66 ][ 222 ],
   alphaCSR[ 66 ][ 223 ],
   alphaCSR[ 66 ][ 224 ],
   alphaCSR[ 66 ][ 225 ],
   alphaCSR[ 66 ][ 226 ],
   alphaCSR[ 66 ][ 227 ],
   alphaCSR[ 66 ][ 228 ],
   alphaCSR[ 66 ][ 229 ],
   alphaCSR[ 66 ][ 230 ],
   alphaCSR[ 66 ][ 231 ],
   alphaCSR[ 66 ][ 232 ],
   alphaCSR[ 66 ][ 233 ],
   alphaCSR[ 66 ][ 234 ],
   alphaCSR[ 66 ][ 235 ],
   alphaCSR[ 66 ][ 236 ],
   alphaCSR[ 66 ][ 237 ],
   alphaCSR[ 66 ][ 238 ],
   alphaCSR[ 66 ][ 239 ],
   alphaCSR[ 66 ][ 240 ],
   alphaCSR[ 66 ][ 241 ],
   alphaCSR[ 66 ][ 242 ],
   alphaCSR[ 66 ][ 243 ],
   alphaCSR[ 66 ][ 244 ],
   alphaCSR[ 66 ][ 245 ],
   alphaCSR[ 66 ][ 246 ],
   alphaCSR[ 66 ][ 247 ],
   alphaCSR[ 66 ][ 248 ],
   alphaCSR[ 66 ][ 249 ],
   alphaCSR[ 66 ][ 250 ],
   alphaCSR[ 66 ][ 251 ],
   alphaCSR[ 66 ][ 252 ],
   alphaCSR[ 66 ][ 253 ],
   alphaCSR[ 66 ][ 254 ],
   alphaCSR[ 66 ][ 255 ],
   alphaCSR[ 66 ][ 256 ],
   alphaCSR[ 66 ][ 257 ],
   alphaCSR[ 66 ][ 258 ],
   alphaCSR[ 66 ][ 259 ],
   alphaCSR[ 66 ][ 260 ],
   alphaCSR[ 66 ][ 261 ],
   alphaCSR[ 66 ][ 262 ],
   alphaCSR[ 66 ][ 263 ],
   alphaCSR[ 66 ][ 264 ],
   alphaCSR[ 66 ][ 265 ],
   alphaCSR[ 66 ][ 266 ],
   alphaCSR[ 66 ][ 267 ],
   alphaCSR[ 66 ][ 268 ],
   alphaCSR[ 66 ][ 269 ],
   alphaCSR[ 66 ][ 270 ],
   alphaCSR[ 66 ][ 271 ],
   alphaCSR[ 66 ][ 272 ],
   alphaCSR[ 66 ][ 273 ],
   alphaCSR[ 66 ][ 274 ],
   alphaCSR[ 66 ][ 275 ],
   alphaCSR[ 66 ][ 276 ],
   alphaCSR[ 66 ][ 277 ],
   alphaCSR[ 66 ][ 278 ],
   alphaCSR[ 66 ][ 279 ],
   alphaCSR[ 66 ][ 280 ],
   alphaCSR[ 66 ][ 281 ],
   alphaCSR[ 66 ][ 282 ],
   alphaCSR[ 66 ][ 283 ],
   alphaCSR[ 66 ][ 284 ],
   alphaCSR[ 66 ][ 285 ],
   alphaCSR[ 66 ][ 286 ],
   alphaCSR[ 66 ][ 287 ],
   alphaCSR[ 66 ][ 288 ],
   alphaCSR[ 66 ][ 289 ],
   alphaCSR[ 66 ][ 290 ],
   alphaCSR[ 66 ][ 291 ],
   alphaCSR[ 66 ][ 292 ],
   alphaCSR[ 66 ][ 293 ],
   alphaCSR[ 66 ][ 294 ],
   alphaCSR[ 66 ][ 295 ],
   alphaCSR[ 66 ][ 296 ],
   alphaCSR[ 66 ][ 297 ],
   alphaCSR[ 66 ][ 298 ],
   alphaCSR[ 66 ][ 299 ],
   alphaCSR[ 66 ][ 300 ],
   alphaCSR[ 66 ][ 301 ],
   alphaCSR[ 66 ][ 302 ],
   alphaCSR[ 66 ][ 303 ],
   alphaCSR[ 66 ][ 304 ],
   alphaCSR[ 66 ][ 305 ],
   alphaCSR[ 66 ][ 306 ],
   alphaCSR[ 66 ][ 307 ],
   alphaCSR[ 66 ][ 308 ],
   alphaCSR[ 66 ][ 309 ],
   alphaCSR[ 66 ][ 310 ],
   alphaCSR[ 66 ][ 311 ],
   alphaCSR[ 66 ][ 312 ],
   alphaCSR[ 66 ][ 313 ],
   alphaCSR[ 66 ][ 314 ],
   alphaCSR[ 66 ][ 315 ],
   alphaCSR[ 66 ][ 316 ],
   alphaCSR[ 66 ][ 317 ],
   alphaCSR[ 66 ][ 318 ],
   alphaCSR[ 66 ][ 319 ],
   alphaCSR[ 66 ][ 320 ],
   alphaCSR[ 66 ][ 321 ],
   alphaCSR[ 66 ][ 322 ],
   alphaCSR[ 66 ][ 323 ],
   alphaCSR[ 66 ][ 324 ],
   alphaCSR[ 66 ][ 325 ],
   alphaCSR[ 66 ][ 326 ],
   alphaCSR[ 66 ][ 327 ],
   alphaCSR[ 66 ][ 328 ],
   alphaCSR[ 66 ][ 329 ],
   alphaCSR[ 66 ][ 330 ],
   alphaCSR[ 66 ][ 331 ],
   alphaCSR[ 66 ][ 332 ],
   alphaCSR[ 66 ][ 333 ],
   alphaCSR[ 66 ][ 334 ],
   alphaCSR[ 66 ][ 335 ],
   alphaCSR[ 66 ][ 336 ],
   alphaCSR[ 66 ][ 337 ],
   alphaCSR[ 66 ][ 338 ],
   alphaCSR[ 66 ][ 339 ],
   alphaCSR[ 66 ][ 340 ],
   alphaCSR[ 66 ][ 341 ],
   alphaCSR[ 66 ][ 342 ],
   alphaCSR[ 66 ][ 343 ],
   alphaCSR[ 66 ][ 344 ],
   alphaCSR[ 66 ][ 345 ],
   alphaCSR[ 66 ][ 346 ],
   alphaCSR[ 66 ][ 347 ],
   alphaCSR[ 66 ][ 348 ],
   alphaCSR[ 66 ][ 349 ],
   alphaCSR[ 66 ][ 350 ],
   alphaCSR[ 66 ][ 351 ],
   alphaCSR[ 66 ][ 352 ],
   alphaCSR[ 66 ][ 353 ],
   alphaCSR[ 66 ][ 354 ],
   alphaCSR[ 66 ][ 355 ],
   alphaCSR[ 66 ][ 356 ],
   alphaCSR[ 66 ][ 357 ],
   alphaCSR[ 66 ][ 358 ],
   alphaCSR[ 66 ][ 359 ],
   alphaCSR[ 66 ][ 360 ],
   alphaCSR[ 66 ][ 361 ],
   alphaCSR[ 66 ][ 362 ],
   alphaCSR[ 66 ][ 363 ],
   alphaCSR[ 66 ][ 364 ],
   alphaCSR[ 66 ][ 365 ],
   alphaCSR[ 66 ][ 366 ],
   alphaCSR[ 66 ][ 367 ],
   alphaCSR[ 66 ][ 368 ],
   alphaCSR[ 66 ][ 369 ],
   alphaCSR[ 66 ][ 370 ],
   alphaCSR[ 66 ][ 371 ],
   alphaCSR[ 66 ][ 372 ],
   alphaCSR[ 66 ][ 373 ],
   alphaCSR[ 66 ][ 374 ],
   alphaCSR[ 66 ][ 375 ],
   alphaCSR[ 66 ][ 376 ],
   alphaCSR[ 66 ][ 377 ],
   alphaCSR[ 66 ][ 378 ],
   alphaCSR[ 66 ][ 379 ],
   alphaCSR[ 66 ][ 380 ],
   alphaCSR[ 66 ][ 381 ],
   alphaCSR[ 66 ][ 382 ],
   alphaCSR[ 66 ][ 383 ],
   alphaCSR[ 67 ][ 0 ],
   alphaCSR[ 67 ][ 1 ],
   alphaCSR[ 67 ][ 2 ],
   alphaCSR[ 67 ][ 3 ],
   alphaCSR[ 67 ][ 4 ],
   alphaCSR[ 67 ][ 5 ],
   alphaCSR[ 67 ][ 6 ],
   alphaCSR[ 67 ][ 7 ],
   alphaCSR[ 67 ][ 8 ],
   alphaCSR[ 67 ][ 9 ],
   alphaCSR[ 67 ][ 10 ],
   alphaCSR[ 67 ][ 11 ],
   alphaCSR[ 67 ][ 12 ],
   alphaCSR[ 67 ][ 13 ],
   alphaCSR[ 67 ][ 14 ],
   alphaCSR[ 67 ][ 15 ],
   alphaCSR[ 67 ][ 16 ],
   alphaCSR[ 67 ][ 17 ],
   alphaCSR[ 67 ][ 18 ],
   alphaCSR[ 67 ][ 19 ],
   alphaCSR[ 67 ][ 20 ],
   alphaCSR[ 67 ][ 21 ],
   alphaCSR[ 67 ][ 22 ],
   alphaCSR[ 67 ][ 23 ],
   alphaCSR[ 67 ][ 24 ],
   alphaCSR[ 67 ][ 25 ],
   alphaCSR[ 67 ][ 26 ],
   alphaCSR[ 67 ][ 27 ],
   alphaCSR[ 67 ][ 28 ],
   alphaCSR[ 67 ][ 29 ],
   alphaCSR[ 67 ][ 30 ],
   alphaCSR[ 67 ][ 31 ],
   alphaCSR[ 67 ][ 32 ],
   alphaCSR[ 67 ][ 33 ],
   alphaCSR[ 67 ][ 34 ],
   alphaCSR[ 67 ][ 35 ],
   alphaCSR[ 67 ][ 36 ],
   alphaCSR[ 67 ][ 37 ],
   alphaCSR[ 67 ][ 38 ],
   alphaCSR[ 67 ][ 39 ],
   alphaCSR[ 67 ][ 40 ],
   alphaCSR[ 67 ][ 41 ],
   alphaCSR[ 67 ][ 42 ],
   alphaCSR[ 67 ][ 43 ],
   alphaCSR[ 67 ][ 44 ],
   alphaCSR[ 67 ][ 45 ],
   alphaCSR[ 67 ][ 46 ],
   alphaCSR[ 67 ][ 47 ],
   alphaCSR[ 67 ][ 48 ],
   alphaCSR[ 67 ][ 49 ],
   alphaCSR[ 67 ][ 50 ],
   alphaCSR[ 67 ][ 51 ],
   alphaCSR[ 67 ][ 52 ],
   alphaCSR[ 67 ][ 53 ],
   alphaCSR[ 67 ][ 54 ],
   alphaCSR[ 67 ][ 55 ],
   alphaCSR[ 67 ][ 56 ],
   alphaCSR[ 67 ][ 57 ],
   alphaCSR[ 67 ][ 58 ],
   alphaCSR[ 67 ][ 59 ],
   alphaCSR[ 67 ][ 60 ],
   alphaCSR[ 67 ][ 61 ],
   alphaCSR[ 67 ][ 62 ],
   alphaCSR[ 67 ][ 63 ],
   alphaCSR[ 67 ][ 64 ],
   alphaCSR[ 67 ][ 65 ],
   alphaCSR[ 67 ][ 66 ],
   alphaCSR[ 67 ][ 67 ],
   alphaCSR[ 67 ][ 68 ],
   alphaCSR[ 67 ][ 69 ],
   alphaCSR[ 67 ][ 70 ],
   alphaCSR[ 67 ][ 71 ],
   alphaCSR[ 67 ][ 72 ],
   alphaCSR[ 67 ][ 73 ],
   alphaCSR[ 67 ][ 74 ],
   alphaCSR[ 67 ][ 75 ],
   alphaCSR[ 67 ][ 76 ],
   alphaCSR[ 67 ][ 77 ],
   alphaCSR[ 67 ][ 78 ],
   alphaCSR[ 67 ][ 79 ],
   alphaCSR[ 67 ][ 80 ],
   alphaCSR[ 67 ][ 81 ],
   alphaCSR[ 67 ][ 82 ],
   alphaCSR[ 67 ][ 83 ],
   alphaCSR[ 67 ][ 84 ],
   alphaCSR[ 67 ][ 85 ],
   alphaCSR[ 67 ][ 86 ],
   alphaCSR[ 67 ][ 87 ],
   alphaCSR[ 67 ][ 88 ],
   alphaCSR[ 67 ][ 89 ],
   alphaCSR[ 67 ][ 90 ],
   alphaCSR[ 67 ][ 91 ],
   alphaCSR[ 67 ][ 92 ],
   alphaCSR[ 67 ][ 93 ],
   alphaCSR[ 67 ][ 94 ],
   alphaCSR[ 67 ][ 95 ],
   alphaCSR[ 67 ][ 96 ],
   alphaCSR[ 67 ][ 97 ],
   alphaCSR[ 67 ][ 98 ],
   alphaCSR[ 67 ][ 99 ],
   alphaCSR[ 67 ][ 100 ],
   alphaCSR[ 67 ][ 101 ],
   alphaCSR[ 67 ][ 102 ],
   alphaCSR[ 67 ][ 103 ],
   alphaCSR[ 67 ][ 104 ],
   alphaCSR[ 67 ][ 105 ],
   alphaCSR[ 67 ][ 106 ],
   alphaCSR[ 67 ][ 107 ],
   alphaCSR[ 67 ][ 108 ],
   alphaCSR[ 67 ][ 109 ],
   alphaCSR[ 67 ][ 110 ],
   alphaCSR[ 67 ][ 111 ],
   alphaCSR[ 67 ][ 112 ],
   alphaCSR[ 67 ][ 113 ],
   alphaCSR[ 67 ][ 114 ],
   alphaCSR[ 67 ][ 115 ],
   alphaCSR[ 67 ][ 116 ],
   alphaCSR[ 67 ][ 117 ],
   alphaCSR[ 67 ][ 118 ],
   alphaCSR[ 67 ][ 119 ],
   alphaCSR[ 67 ][ 120 ],
   alphaCSR[ 67 ][ 121 ],
   alphaCSR[ 67 ][ 122 ],
   alphaCSR[ 67 ][ 123 ],
   alphaCSR[ 67 ][ 124 ],
   alphaCSR[ 67 ][ 125 ],
   alphaCSR[ 67 ][ 126 ],
   alphaCSR[ 67 ][ 127 ],
   alphaCSR[ 67 ][ 128 ],
   alphaCSR[ 67 ][ 129 ],
   alphaCSR[ 67 ][ 130 ],
   alphaCSR[ 67 ][ 131 ],
   alphaCSR[ 67 ][ 132 ],
   alphaCSR[ 67 ][ 133 ],
   alphaCSR[ 67 ][ 134 ],
   alphaCSR[ 67 ][ 135 ],
   alphaCSR[ 67 ][ 136 ],
   alphaCSR[ 67 ][ 137 ],
   alphaCSR[ 67 ][ 138 ],
   alphaCSR[ 67 ][ 139 ],
   alphaCSR[ 67 ][ 140 ],
   alphaCSR[ 67 ][ 141 ],
   alphaCSR[ 67 ][ 142 ],
   alphaCSR[ 67 ][ 143 ],
   alphaCSR[ 67 ][ 144 ],
   alphaCSR[ 67 ][ 145 ],
   alphaCSR[ 67 ][ 146 ],
   alphaCSR[ 67 ][ 147 ],
   alphaCSR[ 67 ][ 148 ],
   alphaCSR[ 67 ][ 149 ],
   alphaCSR[ 67 ][ 150 ],
   alphaCSR[ 67 ][ 151 ],
   alphaCSR[ 67 ][ 152 ],
   alphaCSR[ 67 ][ 153 ],
   alphaCSR[ 67 ][ 154 ],
   alphaCSR[ 67 ][ 155 ],
   alphaCSR[ 67 ][ 156 ],
   alphaCSR[ 67 ][ 157 ],
   alphaCSR[ 67 ][ 158 ],
   alphaCSR[ 67 ][ 159 ],
   alphaCSR[ 67 ][ 160 ],
   alphaCSR[ 67 ][ 161 ],
   alphaCSR[ 67 ][ 162 ],
   alphaCSR[ 67 ][ 163 ],
   alphaCSR[ 67 ][ 164 ],
   alphaCSR[ 67 ][ 165 ],
   alphaCSR[ 67 ][ 166 ],
   alphaCSR[ 67 ][ 167 ],
   alphaCSR[ 67 ][ 168 ],
   alphaCSR[ 67 ][ 169 ],
   alphaCSR[ 67 ][ 170 ],
   alphaCSR[ 67 ][ 171 ],
   alphaCSR[ 67 ][ 172 ],
   alphaCSR[ 67 ][ 173 ],
   alphaCSR[ 67 ][ 174 ],
   alphaCSR[ 67 ][ 175 ],
   alphaCSR[ 67 ][ 176 ],
   alphaCSR[ 67 ][ 177 ],
   alphaCSR[ 67 ][ 178 ],
   alphaCSR[ 67 ][ 179 ],
   alphaCSR[ 67 ][ 180 ],
   alphaCSR[ 67 ][ 181 ],
   alphaCSR[ 67 ][ 182 ],
   alphaCSR[ 67 ][ 183 ],
   alphaCSR[ 67 ][ 184 ],
   alphaCSR[ 67 ][ 185 ],
   alphaCSR[ 67 ][ 186 ],
   alphaCSR[ 67 ][ 187 ],
   alphaCSR[ 67 ][ 188 ],
   alphaCSR[ 67 ][ 189 ],
   alphaCSR[ 67 ][ 190 ],
   alphaCSR[ 67 ][ 191 ],
   alphaCSR[ 67 ][ 192 ],
   alphaCSR[ 67 ][ 193 ],
   alphaCSR[ 67 ][ 194 ],
   alphaCSR[ 67 ][ 195 ],
   alphaCSR[ 67 ][ 196 ],
   alphaCSR[ 67 ][ 197 ],
   alphaCSR[ 67 ][ 198 ],
   alphaCSR[ 67 ][ 199 ],
   alphaCSR[ 67 ][ 200 ],
   alphaCSR[ 67 ][ 201 ],
   alphaCSR[ 67 ][ 202 ],
   alphaCSR[ 67 ][ 203 ],
   alphaCSR[ 67 ][ 204 ],
   alphaCSR[ 67 ][ 205 ],
   alphaCSR[ 67 ][ 206 ],
   alphaCSR[ 67 ][ 207 ],
   alphaCSR[ 67 ][ 208 ],
   alphaCSR[ 67 ][ 209 ],
   alphaCSR[ 67 ][ 210 ],
   alphaCSR[ 67 ][ 211 ],
   alphaCSR[ 67 ][ 212 ],
   alphaCSR[ 67 ][ 213 ],
   alphaCSR[ 67 ][ 214 ],
   alphaCSR[ 67 ][ 215 ],
   alphaCSR[ 67 ][ 216 ],
   alphaCSR[ 67 ][ 217 ],
   alphaCSR[ 67 ][ 218 ],
   alphaCSR[ 67 ][ 219 ],
   alphaCSR[ 67 ][ 220 ],
   alphaCSR[ 67 ][ 221 ],
   alphaCSR[ 67 ][ 222 ],
   alphaCSR[ 67 ][ 223 ],
   alphaCSR[ 67 ][ 224 ],
   alphaCSR[ 67 ][ 225 ],
   alphaCSR[ 67 ][ 226 ],
   alphaCSR[ 67 ][ 227 ],
   alphaCSR[ 67 ][ 228 ],
   alphaCSR[ 67 ][ 229 ],
   alphaCSR[ 67 ][ 230 ],
   alphaCSR[ 67 ][ 231 ],
   alphaCSR[ 67 ][ 232 ],
   alphaCSR[ 67 ][ 233 ],
   alphaCSR[ 67 ][ 234 ],
   alphaCSR[ 67 ][ 235 ],
   alphaCSR[ 67 ][ 236 ],
   alphaCSR[ 67 ][ 237 ],
   alphaCSR[ 67 ][ 238 ],
   alphaCSR[ 67 ][ 239 ],
   alphaCSR[ 67 ][ 240 ],
   alphaCSR[ 67 ][ 241 ],
   alphaCSR[ 67 ][ 242 ],
   alphaCSR[ 67 ][ 243 ],
   alphaCSR[ 67 ][ 244 ],
   alphaCSR[ 67 ][ 245 ],
   alphaCSR[ 67 ][ 246 ],
   alphaCSR[ 67 ][ 247 ],
   alphaCSR[ 67 ][ 248 ],
   alphaCSR[ 67 ][ 249 ],
   alphaCSR[ 67 ][ 250 ],
   alphaCSR[ 67 ][ 251 ],
   alphaCSR[ 67 ][ 252 ],
   alphaCSR[ 67 ][ 253 ],
   alphaCSR[ 67 ][ 254 ],
   alphaCSR[ 67 ][ 255 ],
   alphaCSR[ 67 ][ 256 ],
   alphaCSR[ 67 ][ 257 ],
   alphaCSR[ 67 ][ 258 ],
   alphaCSR[ 67 ][ 259 ],
   alphaCSR[ 67 ][ 260 ],
   alphaCSR[ 67 ][ 261 ],
   alphaCSR[ 67 ][ 262 ],
   alphaCSR[ 67 ][ 263 ],
   alphaCSR[ 67 ][ 264 ],
   alphaCSR[ 67 ][ 265 ],
   alphaCSR[ 67 ][ 266 ],
   alphaCSR[ 67 ][ 267 ],
   alphaCSR[ 67 ][ 268 ],
   alphaCSR[ 67 ][ 269 ],
   alphaCSR[ 67 ][ 270 ],
   alphaCSR[ 67 ][ 271 ],
   alphaCSR[ 67 ][ 272 ],
   alphaCSR[ 67 ][ 273 ],
   alphaCSR[ 67 ][ 274 ],
   alphaCSR[ 67 ][ 275 ],
   alphaCSR[ 67 ][ 276 ],
   alphaCSR[ 67 ][ 277 ],
   alphaCSR[ 67 ][ 278 ],
   alphaCSR[ 67 ][ 279 ],
   alphaCSR[ 67 ][ 280 ],
   alphaCSR[ 67 ][ 281 ],
   alphaCSR[ 67 ][ 282 ],
   alphaCSR[ 67 ][ 283 ],
   alphaCSR[ 67 ][ 284 ],
   alphaCSR[ 67 ][ 285 ],
   alphaCSR[ 67 ][ 286 ],
   alphaCSR[ 67 ][ 287 ],
   alphaCSR[ 67 ][ 288 ],
   alphaCSR[ 67 ][ 289 ],
   alphaCSR[ 67 ][ 290 ],
   alphaCSR[ 67 ][ 291 ],
   alphaCSR[ 67 ][ 292 ],
   alphaCSR[ 67 ][ 293 ],
   alphaCSR[ 67 ][ 294 ],
   alphaCSR[ 67 ][ 295 ],
   alphaCSR[ 67 ][ 296 ],
   alphaCSR[ 67 ][ 297 ],
   alphaCSR[ 67 ][ 298 ],
   alphaCSR[ 67 ][ 299 ],
   alphaCSR[ 67 ][ 300 ],
   alphaCSR[ 67 ][ 301 ],
   alphaCSR[ 67 ][ 302 ],
   alphaCSR[ 67 ][ 303 ],
   alphaCSR[ 67 ][ 304 ],
   alphaCSR[ 67 ][ 305 ],
   alphaCSR[ 67 ][ 306 ],
   alphaCSR[ 67 ][ 307 ],
   alphaCSR[ 67 ][ 308 ],
   alphaCSR[ 67 ][ 309 ],
   alphaCSR[ 67 ][ 310 ],
   alphaCSR[ 67 ][ 311 ],
   alphaCSR[ 67 ][ 312 ],
   alphaCSR[ 67 ][ 313 ],
   alphaCSR[ 67 ][ 314 ],
   alphaCSR[ 67 ][ 315 ],
   alphaCSR[ 67 ][ 316 ],
   alphaCSR[ 67 ][ 317 ],
   alphaCSR[ 67 ][ 318 ],
   alphaCSR[ 67 ][ 319 ],
   alphaCSR[ 67 ][ 320 ],
   alphaCSR[ 67 ][ 321 ],
   alphaCSR[ 67 ][ 322 ],
   alphaCSR[ 67 ][ 323 ],
   alphaCSR[ 67 ][ 324 ],
   alphaCSR[ 67 ][ 325 ],
   alphaCSR[ 67 ][ 326 ],
   alphaCSR[ 67 ][ 327 ],
   alphaCSR[ 67 ][ 328 ],
   alphaCSR[ 67 ][ 329 ],
   alphaCSR[ 67 ][ 330 ],
   alphaCSR[ 67 ][ 331 ],
   alphaCSR[ 67 ][ 332 ],
   alphaCSR[ 67 ][ 333 ],
   alphaCSR[ 67 ][ 334 ],
   alphaCSR[ 67 ][ 335 ],
   alphaCSR[ 67 ][ 336 ],
   alphaCSR[ 67 ][ 337 ],
   alphaCSR[ 67 ][ 338 ],
   alphaCSR[ 67 ][ 339 ],
   alphaCSR[ 67 ][ 340 ],
   alphaCSR[ 67 ][ 341 ],
   alphaCSR[ 67 ][ 342 ],
   alphaCSR[ 67 ][ 343 ],
   alphaCSR[ 67 ][ 344 ],
   alphaCSR[ 67 ][ 345 ],
   alphaCSR[ 67 ][ 346 ],
   alphaCSR[ 67 ][ 347 ],
   alphaCSR[ 67 ][ 348 ],
   alphaCSR[ 67 ][ 349 ],
   alphaCSR[ 67 ][ 350 ],
   alphaCSR[ 67 ][ 351 ],
   alphaCSR[ 67 ][ 352 ],
   alphaCSR[ 67 ][ 353 ],
   alphaCSR[ 67 ][ 354 ],
   alphaCSR[ 67 ][ 355 ],
   alphaCSR[ 67 ][ 356 ],
   alphaCSR[ 67 ][ 357 ],
   alphaCSR[ 67 ][ 358 ],
   alphaCSR[ 67 ][ 359 ],
   alphaCSR[ 67 ][ 360 ],
   alphaCSR[ 67 ][ 361 ],
   alphaCSR[ 67 ][ 362 ],
   alphaCSR[ 67 ][ 363 ],
   alphaCSR[ 67 ][ 364 ],
   alphaCSR[ 67 ][ 365 ],
   alphaCSR[ 67 ][ 366 ],
   alphaCSR[ 67 ][ 367 ],
   alphaCSR[ 67 ][ 368 ],
   alphaCSR[ 67 ][ 369 ],
   alphaCSR[ 67 ][ 370 ],
   alphaCSR[ 67 ][ 371 ],
   alphaCSR[ 67 ][ 372 ],
   alphaCSR[ 67 ][ 373 ],
   alphaCSR[ 67 ][ 374 ],
   alphaCSR[ 67 ][ 375 ],
   alphaCSR[ 67 ][ 376 ],
   alphaCSR[ 67 ][ 377 ],
   alphaCSR[ 67 ][ 378 ],
   alphaCSR[ 67 ][ 379 ],
   alphaCSR[ 67 ][ 380 ],
   alphaCSR[ 67 ][ 381 ],
   alphaCSR[ 67 ][ 382 ],
   alphaCSR[ 67 ][ 383 ],
   alphaCSR[ 68 ][ 0 ],
   alphaCSR[ 68 ][ 1 ],
   alphaCSR[ 68 ][ 2 ],
   alphaCSR[ 68 ][ 3 ],
   alphaCSR[ 68 ][ 4 ],
   alphaCSR[ 68 ][ 5 ],
   alphaCSR[ 68 ][ 6 ],
   alphaCSR[ 68 ][ 7 ],
   alphaCSR[ 68 ][ 8 ],
   alphaCSR[ 68 ][ 9 ],
   alphaCSR[ 68 ][ 10 ],
   alphaCSR[ 68 ][ 11 ],
   alphaCSR[ 68 ][ 12 ],
   alphaCSR[ 68 ][ 13 ],
   alphaCSR[ 68 ][ 14 ],
   alphaCSR[ 68 ][ 15 ],
   alphaCSR[ 68 ][ 16 ],
   alphaCSR[ 68 ][ 17 ],
   alphaCSR[ 68 ][ 18 ],
   alphaCSR[ 68 ][ 19 ],
   alphaCSR[ 68 ][ 20 ],
   alphaCSR[ 68 ][ 21 ],
   alphaCSR[ 68 ][ 22 ],
   alphaCSR[ 68 ][ 23 ],
   alphaCSR[ 68 ][ 24 ],
   alphaCSR[ 68 ][ 25 ],
   alphaCSR[ 68 ][ 26 ],
   alphaCSR[ 68 ][ 27 ],
   alphaCSR[ 68 ][ 28 ],
   alphaCSR[ 68 ][ 29 ],
   alphaCSR[ 68 ][ 30 ],
   alphaCSR[ 68 ][ 31 ],
   alphaCSR[ 68 ][ 32 ],
   alphaCSR[ 68 ][ 33 ],
   alphaCSR[ 68 ][ 34 ],
   alphaCSR[ 68 ][ 35 ],
   alphaCSR[ 68 ][ 36 ],
   alphaCSR[ 68 ][ 37 ],
   alphaCSR[ 68 ][ 38 ],
   alphaCSR[ 68 ][ 39 ],
   alphaCSR[ 68 ][ 40 ],
   alphaCSR[ 68 ][ 41 ],
   alphaCSR[ 68 ][ 42 ],
   alphaCSR[ 68 ][ 43 ],
   alphaCSR[ 68 ][ 44 ],
   alphaCSR[ 68 ][ 45 ],
   alphaCSR[ 68 ][ 46 ],
   alphaCSR[ 68 ][ 47 ],
   alphaCSR[ 68 ][ 48 ],
   alphaCSR[ 68 ][ 49 ],
   alphaCSR[ 68 ][ 50 ],
   alphaCSR[ 68 ][ 51 ],
   alphaCSR[ 68 ][ 52 ],
   alphaCSR[ 68 ][ 53 ],
   alphaCSR[ 68 ][ 54 ],
   alphaCSR[ 68 ][ 55 ],
   alphaCSR[ 68 ][ 56 ],
   alphaCSR[ 68 ][ 57 ],
   alphaCSR[ 68 ][ 58 ],
   alphaCSR[ 68 ][ 59 ],
   alphaCSR[ 68 ][ 60 ],
   alphaCSR[ 68 ][ 61 ],
   alphaCSR[ 68 ][ 62 ],
   alphaCSR[ 68 ][ 63 ],
   alphaCSR[ 68 ][ 64 ],
   alphaCSR[ 68 ][ 65 ],
   alphaCSR[ 68 ][ 66 ],
   alphaCSR[ 68 ][ 67 ],
   alphaCSR[ 68 ][ 68 ],
   alphaCSR[ 68 ][ 69 ],
   alphaCSR[ 68 ][ 70 ],
   alphaCSR[ 68 ][ 71 ],
   alphaCSR[ 68 ][ 72 ],
   alphaCSR[ 68 ][ 73 ],
   alphaCSR[ 68 ][ 74 ],
   alphaCSR[ 68 ][ 75 ],
   alphaCSR[ 68 ][ 76 ],
   alphaCSR[ 68 ][ 77 ],
   alphaCSR[ 68 ][ 78 ],
   alphaCSR[ 68 ][ 79 ],
   alphaCSR[ 68 ][ 80 ],
   alphaCSR[ 68 ][ 81 ],
   alphaCSR[ 68 ][ 82 ],
   alphaCSR[ 68 ][ 83 ],
   alphaCSR[ 68 ][ 84 ],
   alphaCSR[ 68 ][ 85 ],
   alphaCSR[ 68 ][ 86 ],
   alphaCSR[ 68 ][ 87 ],
   alphaCSR[ 68 ][ 88 ],
   alphaCSR[ 68 ][ 89 ],
   alphaCSR[ 68 ][ 90 ],
   alphaCSR[ 68 ][ 91 ],
   alphaCSR[ 68 ][ 92 ],
   alphaCSR[ 68 ][ 93 ],
   alphaCSR[ 68 ][ 94 ],
   alphaCSR[ 68 ][ 95 ],
   alphaCSR[ 68 ][ 96 ],
   alphaCSR[ 68 ][ 97 ],
   alphaCSR[ 68 ][ 98 ],
   alphaCSR[ 68 ][ 99 ],
   alphaCSR[ 68 ][ 100 ],
   alphaCSR[ 68 ][ 101 ],
   alphaCSR[ 68 ][ 102 ],
   alphaCSR[ 68 ][ 103 ],
   alphaCSR[ 68 ][ 104 ],
   alphaCSR[ 68 ][ 105 ],
   alphaCSR[ 68 ][ 106 ],
   alphaCSR[ 68 ][ 107 ],
   alphaCSR[ 68 ][ 108 ],
   alphaCSR[ 68 ][ 109 ],
   alphaCSR[ 68 ][ 110 ],
   alphaCSR[ 68 ][ 111 ],
   alphaCSR[ 68 ][ 112 ],
   alphaCSR[ 68 ][ 113 ],
   alphaCSR[ 68 ][ 114 ],
   alphaCSR[ 68 ][ 115 ],
   alphaCSR[ 68 ][ 116 ],
   alphaCSR[ 68 ][ 117 ],
   alphaCSR[ 68 ][ 118 ],
   alphaCSR[ 68 ][ 119 ],
   alphaCSR[ 68 ][ 120 ],
   alphaCSR[ 68 ][ 121 ],
   alphaCSR[ 68 ][ 122 ],
   alphaCSR[ 68 ][ 123 ],
   alphaCSR[ 68 ][ 124 ],
   alphaCSR[ 68 ][ 125 ],
   alphaCSR[ 68 ][ 126 ],
   alphaCSR[ 68 ][ 127 ],
   alphaCSR[ 68 ][ 128 ],
   alphaCSR[ 68 ][ 129 ],
   alphaCSR[ 68 ][ 130 ],
   alphaCSR[ 68 ][ 131 ],
   alphaCSR[ 68 ][ 132 ],
   alphaCSR[ 68 ][ 133 ],
   alphaCSR[ 68 ][ 134 ],
   alphaCSR[ 68 ][ 135 ],
   alphaCSR[ 68 ][ 136 ],
   alphaCSR[ 68 ][ 137 ],
   alphaCSR[ 68 ][ 138 ],
   alphaCSR[ 68 ][ 139 ],
   alphaCSR[ 68 ][ 140 ],
   alphaCSR[ 68 ][ 141 ],
   alphaCSR[ 68 ][ 142 ],
   alphaCSR[ 68 ][ 143 ],
   alphaCSR[ 68 ][ 144 ],
   alphaCSR[ 68 ][ 145 ],
   alphaCSR[ 68 ][ 146 ],
   alphaCSR[ 68 ][ 147 ],
   alphaCSR[ 68 ][ 148 ],
   alphaCSR[ 68 ][ 149 ],
   alphaCSR[ 68 ][ 150 ],
   alphaCSR[ 68 ][ 151 ],
   alphaCSR[ 68 ][ 152 ],
   alphaCSR[ 68 ][ 153 ],
   alphaCSR[ 68 ][ 154 ],
   alphaCSR[ 68 ][ 155 ],
   alphaCSR[ 68 ][ 156 ],
   alphaCSR[ 68 ][ 157 ],
   alphaCSR[ 68 ][ 158 ],
   alphaCSR[ 68 ][ 159 ],
   alphaCSR[ 68 ][ 160 ],
   alphaCSR[ 68 ][ 161 ],
   alphaCSR[ 68 ][ 162 ],
   alphaCSR[ 68 ][ 163 ],
   alphaCSR[ 68 ][ 164 ],
   alphaCSR[ 68 ][ 165 ],
   alphaCSR[ 68 ][ 166 ],
   alphaCSR[ 68 ][ 167 ],
   alphaCSR[ 68 ][ 168 ],
   alphaCSR[ 68 ][ 169 ],
   alphaCSR[ 68 ][ 170 ],
   alphaCSR[ 68 ][ 171 ],
   alphaCSR[ 68 ][ 172 ],
   alphaCSR[ 68 ][ 173 ],
   alphaCSR[ 68 ][ 174 ],
   alphaCSR[ 68 ][ 175 ],
   alphaCSR[ 68 ][ 176 ],
   alphaCSR[ 68 ][ 177 ],
   alphaCSR[ 68 ][ 178 ],
   alphaCSR[ 68 ][ 179 ],
   alphaCSR[ 68 ][ 180 ],
   alphaCSR[ 68 ][ 181 ],
   alphaCSR[ 68 ][ 182 ],
   alphaCSR[ 68 ][ 183 ],
   alphaCSR[ 68 ][ 184 ],
   alphaCSR[ 68 ][ 185 ],
   alphaCSR[ 68 ][ 186 ],
   alphaCSR[ 68 ][ 187 ],
   alphaCSR[ 68 ][ 188 ],
   alphaCSR[ 68 ][ 189 ],
   alphaCSR[ 68 ][ 190 ],
   alphaCSR[ 68 ][ 191 ],
   alphaCSR[ 68 ][ 192 ],
   alphaCSR[ 68 ][ 193 ],
   alphaCSR[ 68 ][ 194 ],
   alphaCSR[ 68 ][ 195 ],
   alphaCSR[ 68 ][ 196 ],
   alphaCSR[ 68 ][ 197 ],
   alphaCSR[ 68 ][ 198 ],
   alphaCSR[ 68 ][ 199 ],
   alphaCSR[ 68 ][ 200 ],
   alphaCSR[ 68 ][ 201 ],
   alphaCSR[ 68 ][ 202 ],
   alphaCSR[ 68 ][ 203 ],
   alphaCSR[ 68 ][ 204 ],
   alphaCSR[ 68 ][ 205 ],
   alphaCSR[ 68 ][ 206 ],
   alphaCSR[ 68 ][ 207 ],
   alphaCSR[ 68 ][ 208 ],
   alphaCSR[ 68 ][ 209 ],
   alphaCSR[ 68 ][ 210 ],
   alphaCSR[ 68 ][ 211 ],
   alphaCSR[ 68 ][ 212 ],
   alphaCSR[ 68 ][ 213 ],
   alphaCSR[ 68 ][ 214 ],
   alphaCSR[ 68 ][ 215 ],
   alphaCSR[ 68 ][ 216 ],
   alphaCSR[ 68 ][ 217 ],
   alphaCSR[ 68 ][ 218 ],
   alphaCSR[ 68 ][ 219 ],
   alphaCSR[ 68 ][ 220 ],
   alphaCSR[ 68 ][ 221 ],
   alphaCSR[ 68 ][ 222 ],
   alphaCSR[ 68 ][ 223 ],
   alphaCSR[ 68 ][ 224 ],
   alphaCSR[ 68 ][ 225 ],
   alphaCSR[ 68 ][ 226 ],
   alphaCSR[ 68 ][ 227 ],
   alphaCSR[ 68 ][ 228 ],
   alphaCSR[ 68 ][ 229 ],
   alphaCSR[ 68 ][ 230 ],
   alphaCSR[ 68 ][ 231 ],
   alphaCSR[ 68 ][ 232 ],
   alphaCSR[ 68 ][ 233 ],
   alphaCSR[ 68 ][ 234 ],
   alphaCSR[ 68 ][ 235 ],
   alphaCSR[ 68 ][ 236 ],
   alphaCSR[ 68 ][ 237 ],
   alphaCSR[ 68 ][ 238 ],
   alphaCSR[ 68 ][ 239 ],
   alphaCSR[ 68 ][ 240 ],
   alphaCSR[ 68 ][ 241 ],
   alphaCSR[ 68 ][ 242 ],
   alphaCSR[ 68 ][ 243 ],
   alphaCSR[ 68 ][ 244 ],
   alphaCSR[ 68 ][ 245 ],
   alphaCSR[ 68 ][ 246 ],
   alphaCSR[ 68 ][ 247 ],
   alphaCSR[ 68 ][ 248 ],
   alphaCSR[ 68 ][ 249 ],
   alphaCSR[ 68 ][ 250 ],
   alphaCSR[ 68 ][ 251 ],
   alphaCSR[ 68 ][ 252 ],
   alphaCSR[ 68 ][ 253 ],
   alphaCSR[ 68 ][ 254 ],
   alphaCSR[ 68 ][ 255 ],
   alphaCSR[ 68 ][ 256 ],
   alphaCSR[ 68 ][ 257 ],
   alphaCSR[ 68 ][ 258 ],
   alphaCSR[ 68 ][ 259 ],
   alphaCSR[ 68 ][ 260 ],
   alphaCSR[ 68 ][ 261 ],
   alphaCSR[ 68 ][ 262 ],
   alphaCSR[ 68 ][ 263 ],
   alphaCSR[ 68 ][ 264 ],
   alphaCSR[ 68 ][ 265 ],
   alphaCSR[ 68 ][ 266 ],
   alphaCSR[ 68 ][ 267 ],
   alphaCSR[ 68 ][ 268 ],
   alphaCSR[ 68 ][ 269 ],
   alphaCSR[ 68 ][ 270 ],
   alphaCSR[ 68 ][ 271 ],
   alphaCSR[ 68 ][ 272 ],
   alphaCSR[ 68 ][ 273 ],
   alphaCSR[ 68 ][ 274 ],
   alphaCSR[ 68 ][ 275 ],
   alphaCSR[ 68 ][ 276 ],
   alphaCSR[ 68 ][ 277 ],
   alphaCSR[ 68 ][ 278 ],
   alphaCSR[ 68 ][ 279 ],
   alphaCSR[ 68 ][ 280 ],
   alphaCSR[ 68 ][ 281 ],
   alphaCSR[ 68 ][ 282 ],
   alphaCSR[ 68 ][ 283 ],
   alphaCSR[ 68 ][ 284 ],
   alphaCSR[ 68 ][ 285 ],
   alphaCSR[ 68 ][ 286 ],
   alphaCSR[ 68 ][ 287 ],
   alphaCSR[ 68 ][ 288 ],
   alphaCSR[ 68 ][ 289 ],
   alphaCSR[ 68 ][ 290 ],
   alphaCSR[ 68 ][ 291 ],
   alphaCSR[ 68 ][ 292 ],
   alphaCSR[ 68 ][ 293 ],
   alphaCSR[ 68 ][ 294 ],
   alphaCSR[ 68 ][ 295 ],
   alphaCSR[ 68 ][ 296 ],
   alphaCSR[ 68 ][ 297 ],
   alphaCSR[ 68 ][ 298 ],
   alphaCSR[ 68 ][ 299 ],
   alphaCSR[ 68 ][ 300 ],
   alphaCSR[ 68 ][ 301 ],
   alphaCSR[ 68 ][ 302 ],
   alphaCSR[ 68 ][ 303 ],
   alphaCSR[ 68 ][ 304 ],
   alphaCSR[ 68 ][ 305 ],
   alphaCSR[ 68 ][ 306 ],
   alphaCSR[ 68 ][ 307 ],
   alphaCSR[ 68 ][ 308 ],
   alphaCSR[ 68 ][ 309 ],
   alphaCSR[ 68 ][ 310 ],
   alphaCSR[ 68 ][ 311 ],
   alphaCSR[ 68 ][ 312 ],
   alphaCSR[ 68 ][ 313 ],
   alphaCSR[ 68 ][ 314 ],
   alphaCSR[ 68 ][ 315 ],
   alphaCSR[ 68 ][ 316 ],
   alphaCSR[ 68 ][ 317 ],
   alphaCSR[ 68 ][ 318 ],
   alphaCSR[ 68 ][ 319 ],
   alphaCSR[ 68 ][ 320 ],
   alphaCSR[ 68 ][ 321 ],
   alphaCSR[ 68 ][ 322 ],
   alphaCSR[ 68 ][ 323 ],
   alphaCSR[ 68 ][ 324 ],
   alphaCSR[ 68 ][ 325 ],
   alphaCSR[ 68 ][ 326 ],
   alphaCSR[ 68 ][ 327 ],
   alphaCSR[ 68 ][ 328 ],
   alphaCSR[ 68 ][ 329 ],
   alphaCSR[ 68 ][ 330 ],
   alphaCSR[ 68 ][ 331 ],
   alphaCSR[ 68 ][ 332 ],
   alphaCSR[ 68 ][ 333 ],
   alphaCSR[ 68 ][ 334 ],
   alphaCSR[ 68 ][ 335 ],
   alphaCSR[ 68 ][ 336 ],
   alphaCSR[ 68 ][ 337 ],
   alphaCSR[ 68 ][ 338 ],
   alphaCSR[ 68 ][ 339 ],
   alphaCSR[ 68 ][ 340 ],
   alphaCSR[ 68 ][ 341 ],
   alphaCSR[ 68 ][ 342 ],
   alphaCSR[ 68 ][ 343 ],
   alphaCSR[ 68 ][ 344 ],
   alphaCSR[ 68 ][ 345 ],
   alphaCSR[ 68 ][ 346 ],
   alphaCSR[ 68 ][ 347 ],
   alphaCSR[ 68 ][ 348 ],
   alphaCSR[ 68 ][ 349 ],
   alphaCSR[ 68 ][ 350 ],
   alphaCSR[ 68 ][ 351 ],
   alphaCSR[ 68 ][ 352 ],
   alphaCSR[ 68 ][ 353 ],
   alphaCSR[ 68 ][ 354 ],
   alphaCSR[ 68 ][ 355 ],
   alphaCSR[ 68 ][ 356 ],
   alphaCSR[ 68 ][ 357 ],
   alphaCSR[ 68 ][ 358 ],
   alphaCSR[ 68 ][ 359 ],
   alphaCSR[ 68 ][ 360 ],
   alphaCSR[ 68 ][ 361 ],
   alphaCSR[ 68 ][ 362 ],
   alphaCSR[ 68 ][ 363 ],
   alphaCSR[ 68 ][ 364 ],
   alphaCSR[ 68 ][ 365 ],
   alphaCSR[ 68 ][ 366 ],
   alphaCSR[ 68 ][ 367 ],
   alphaCSR[ 68 ][ 368 ],
   alphaCSR[ 68 ][ 369 ],
   alphaCSR[ 68 ][ 370 ],
   alphaCSR[ 68 ][ 371 ],
   alphaCSR[ 68 ][ 372 ],
   alphaCSR[ 68 ][ 373 ],
   alphaCSR[ 68 ][ 374 ],
   alphaCSR[ 68 ][ 375 ],
   alphaCSR[ 68 ][ 376 ],
   alphaCSR[ 68 ][ 377 ],
   alphaCSR[ 68 ][ 378 ],
   alphaCSR[ 68 ][ 379 ],
   alphaCSR[ 68 ][ 380 ],
   alphaCSR[ 68 ][ 381 ],
   alphaCSR[ 68 ][ 382 ],
   alphaCSR[ 68 ][ 383 ],
   alphaCSR[ 69 ][ 0 ],
   alphaCSR[ 69 ][ 1 ],
   alphaCSR[ 69 ][ 2 ],
   alphaCSR[ 69 ][ 3 ],
   alphaCSR[ 69 ][ 4 ],
   alphaCSR[ 69 ][ 5 ],
   alphaCSR[ 69 ][ 6 ],
   alphaCSR[ 69 ][ 7 ],
   alphaCSR[ 69 ][ 8 ],
   alphaCSR[ 69 ][ 9 ],
   alphaCSR[ 69 ][ 10 ],
   alphaCSR[ 69 ][ 11 ],
   alphaCSR[ 69 ][ 12 ],
   alphaCSR[ 69 ][ 13 ],
   alphaCSR[ 69 ][ 14 ],
   alphaCSR[ 69 ][ 15 ],
   alphaCSR[ 69 ][ 16 ],
   alphaCSR[ 69 ][ 17 ],
   alphaCSR[ 69 ][ 18 ],
   alphaCSR[ 69 ][ 19 ],
   alphaCSR[ 69 ][ 20 ],
   alphaCSR[ 69 ][ 21 ],
   alphaCSR[ 69 ][ 22 ],
   alphaCSR[ 69 ][ 23 ],
   alphaCSR[ 69 ][ 24 ],
   alphaCSR[ 69 ][ 25 ],
   alphaCSR[ 69 ][ 26 ],
   alphaCSR[ 69 ][ 27 ],
   alphaCSR[ 69 ][ 28 ],
   alphaCSR[ 69 ][ 29 ],
   alphaCSR[ 69 ][ 30 ],
   alphaCSR[ 69 ][ 31 ],
   alphaCSR[ 69 ][ 32 ],
   alphaCSR[ 69 ][ 33 ],
   alphaCSR[ 69 ][ 34 ],
   alphaCSR[ 69 ][ 35 ],
   alphaCSR[ 69 ][ 36 ],
   alphaCSR[ 69 ][ 37 ],
   alphaCSR[ 69 ][ 38 ],
   alphaCSR[ 69 ][ 39 ],
   alphaCSR[ 69 ][ 40 ],
   alphaCSR[ 69 ][ 41 ],
   alphaCSR[ 69 ][ 42 ],
   alphaCSR[ 69 ][ 43 ],
   alphaCSR[ 69 ][ 44 ],
   alphaCSR[ 69 ][ 45 ],
   alphaCSR[ 69 ][ 46 ],
   alphaCSR[ 69 ][ 47 ],
   alphaCSR[ 69 ][ 48 ],
   alphaCSR[ 69 ][ 49 ],
   alphaCSR[ 69 ][ 50 ],
   alphaCSR[ 69 ][ 51 ],
   alphaCSR[ 69 ][ 52 ],
   alphaCSR[ 69 ][ 53 ],
   alphaCSR[ 69 ][ 54 ],
   alphaCSR[ 69 ][ 55 ],
   alphaCSR[ 69 ][ 56 ],
   alphaCSR[ 69 ][ 57 ],
   alphaCSR[ 69 ][ 58 ],
   alphaCSR[ 69 ][ 59 ],
   alphaCSR[ 69 ][ 60 ],
   alphaCSR[ 69 ][ 61 ],
   alphaCSR[ 69 ][ 62 ],
   alphaCSR[ 69 ][ 63 ],
   alphaCSR[ 69 ][ 64 ],
   alphaCSR[ 69 ][ 65 ],
   alphaCSR[ 69 ][ 66 ],
   alphaCSR[ 69 ][ 67 ],
   alphaCSR[ 69 ][ 68 ],
   alphaCSR[ 69 ][ 69 ],
   alphaCSR[ 69 ][ 70 ],
   alphaCSR[ 69 ][ 71 ],
   alphaCSR[ 69 ][ 72 ],
   alphaCSR[ 69 ][ 73 ],
   alphaCSR[ 69 ][ 74 ],
   alphaCSR[ 69 ][ 75 ],
   alphaCSR[ 69 ][ 76 ],
   alphaCSR[ 69 ][ 77 ],
   alphaCSR[ 69 ][ 78 ],
   alphaCSR[ 69 ][ 79 ],
   alphaCSR[ 69 ][ 80 ],
   alphaCSR[ 69 ][ 81 ],
   alphaCSR[ 69 ][ 82 ],
   alphaCSR[ 69 ][ 83 ],
   alphaCSR[ 69 ][ 84 ],
   alphaCSR[ 69 ][ 85 ],
   alphaCSR[ 69 ][ 86 ],
   alphaCSR[ 69 ][ 87 ],
   alphaCSR[ 69 ][ 88 ],
   alphaCSR[ 69 ][ 89 ],
   alphaCSR[ 69 ][ 90 ],
   alphaCSR[ 69 ][ 91 ],
   alphaCSR[ 69 ][ 92 ],
   alphaCSR[ 69 ][ 93 ],
   alphaCSR[ 69 ][ 94 ],
   alphaCSR[ 69 ][ 95 ],
   alphaCSR[ 69 ][ 96 ],
   alphaCSR[ 69 ][ 97 ],
   alphaCSR[ 69 ][ 98 ],
   alphaCSR[ 69 ][ 99 ],
   alphaCSR[ 69 ][ 100 ],
   alphaCSR[ 69 ][ 101 ],
   alphaCSR[ 69 ][ 102 ],
   alphaCSR[ 69 ][ 103 ],
   alphaCSR[ 69 ][ 104 ],
   alphaCSR[ 69 ][ 105 ],
   alphaCSR[ 69 ][ 106 ],
   alphaCSR[ 69 ][ 107 ],
   alphaCSR[ 69 ][ 108 ],
   alphaCSR[ 69 ][ 109 ],
   alphaCSR[ 69 ][ 110 ],
   alphaCSR[ 69 ][ 111 ],
   alphaCSR[ 69 ][ 112 ],
   alphaCSR[ 69 ][ 113 ],
   alphaCSR[ 69 ][ 114 ],
   alphaCSR[ 69 ][ 115 ],
   alphaCSR[ 69 ][ 116 ],
   alphaCSR[ 69 ][ 117 ],
   alphaCSR[ 69 ][ 118 ],
   alphaCSR[ 69 ][ 119 ],
   alphaCSR[ 69 ][ 120 ],
   alphaCSR[ 69 ][ 121 ],
   alphaCSR[ 69 ][ 122 ],
   alphaCSR[ 69 ][ 123 ],
   alphaCSR[ 69 ][ 124 ],
   alphaCSR[ 69 ][ 125 ],
   alphaCSR[ 69 ][ 126 ],
   alphaCSR[ 69 ][ 127 ],
   alphaCSR[ 69 ][ 128 ],
   alphaCSR[ 69 ][ 129 ],
   alphaCSR[ 69 ][ 130 ],
   alphaCSR[ 69 ][ 131 ],
   alphaCSR[ 69 ][ 132 ],
   alphaCSR[ 69 ][ 133 ],
   alphaCSR[ 69 ][ 134 ],
   alphaCSR[ 69 ][ 135 ],
   alphaCSR[ 69 ][ 136 ],
   alphaCSR[ 69 ][ 137 ],
   alphaCSR[ 69 ][ 138 ],
   alphaCSR[ 69 ][ 139 ],
   alphaCSR[ 69 ][ 140 ],
   alphaCSR[ 69 ][ 141 ],
   alphaCSR[ 69 ][ 142 ],
   alphaCSR[ 69 ][ 143 ],
   alphaCSR[ 69 ][ 144 ],
   alphaCSR[ 69 ][ 145 ],
   alphaCSR[ 69 ][ 146 ],
   alphaCSR[ 69 ][ 147 ],
   alphaCSR[ 69 ][ 148 ],
   alphaCSR[ 69 ][ 149 ],
   alphaCSR[ 69 ][ 150 ],
   alphaCSR[ 69 ][ 151 ],
   alphaCSR[ 69 ][ 152 ],
   alphaCSR[ 69 ][ 153 ],
   alphaCSR[ 69 ][ 154 ],
   alphaCSR[ 69 ][ 155 ],
   alphaCSR[ 69 ][ 156 ],
   alphaCSR[ 69 ][ 157 ],
   alphaCSR[ 69 ][ 158 ],
   alphaCSR[ 69 ][ 159 ],
   alphaCSR[ 69 ][ 160 ],
   alphaCSR[ 69 ][ 161 ],
   alphaCSR[ 69 ][ 162 ],
   alphaCSR[ 69 ][ 163 ],
   alphaCSR[ 69 ][ 164 ],
   alphaCSR[ 69 ][ 165 ],
   alphaCSR[ 69 ][ 166 ],
   alphaCSR[ 69 ][ 167 ],
   alphaCSR[ 69 ][ 168 ],
   alphaCSR[ 69 ][ 169 ],
   alphaCSR[ 69 ][ 170 ],
   alphaCSR[ 69 ][ 171 ],
   alphaCSR[ 69 ][ 172 ],
   alphaCSR[ 69 ][ 173 ],
   alphaCSR[ 69 ][ 174 ],
   alphaCSR[ 69 ][ 175 ],
   alphaCSR[ 69 ][ 176 ],
   alphaCSR[ 69 ][ 177 ],
   alphaCSR[ 69 ][ 178 ],
   alphaCSR[ 69 ][ 179 ],
   alphaCSR[ 69 ][ 180 ],
   alphaCSR[ 69 ][ 181 ],
   alphaCSR[ 69 ][ 182 ],
   alphaCSR[ 69 ][ 183 ],
   alphaCSR[ 69 ][ 184 ],
   alphaCSR[ 69 ][ 185 ],
   alphaCSR[ 69 ][ 186 ],
   alphaCSR[ 69 ][ 187 ],
   alphaCSR[ 69 ][ 188 ],
   alphaCSR[ 69 ][ 189 ],
   alphaCSR[ 69 ][ 190 ],
   alphaCSR[ 69 ][ 191 ],
   alphaCSR[ 69 ][ 192 ],
   alphaCSR[ 69 ][ 193 ],
   alphaCSR[ 69 ][ 194 ],
   alphaCSR[ 69 ][ 195 ],
   alphaCSR[ 69 ][ 196 ],
   alphaCSR[ 69 ][ 197 ],
   alphaCSR[ 69 ][ 198 ],
   alphaCSR[ 69 ][ 199 ],
   alphaCSR[ 69 ][ 200 ],
   alphaCSR[ 69 ][ 201 ],
   alphaCSR[ 69 ][ 202 ],
   alphaCSR[ 69 ][ 203 ],
   alphaCSR[ 69 ][ 204 ],
   alphaCSR[ 69 ][ 205 ],
   alphaCSR[ 69 ][ 206 ],
   alphaCSR[ 69 ][ 207 ],
   alphaCSR[ 69 ][ 208 ],
   alphaCSR[ 69 ][ 209 ],
   alphaCSR[ 69 ][ 210 ],
   alphaCSR[ 69 ][ 211 ],
   alphaCSR[ 69 ][ 212 ],
   alphaCSR[ 69 ][ 213 ],
   alphaCSR[ 69 ][ 214 ],
   alphaCSR[ 69 ][ 215 ],
   alphaCSR[ 69 ][ 216 ],
   alphaCSR[ 69 ][ 217 ],
   alphaCSR[ 69 ][ 218 ],
   alphaCSR[ 69 ][ 219 ],
   alphaCSR[ 69 ][ 220 ],
   alphaCSR[ 69 ][ 221 ],
   alphaCSR[ 69 ][ 222 ],
   alphaCSR[ 69 ][ 223 ],
   alphaCSR[ 69 ][ 224 ],
   alphaCSR[ 69 ][ 225 ],
   alphaCSR[ 69 ][ 226 ],
   alphaCSR[ 69 ][ 227 ],
   alphaCSR[ 69 ][ 228 ],
   alphaCSR[ 69 ][ 229 ],
   alphaCSR[ 69 ][ 230 ],
   alphaCSR[ 69 ][ 231 ],
   alphaCSR[ 69 ][ 232 ],
   alphaCSR[ 69 ][ 233 ],
   alphaCSR[ 69 ][ 234 ],
   alphaCSR[ 69 ][ 235 ],
   alphaCSR[ 69 ][ 236 ],
   alphaCSR[ 69 ][ 237 ],
   alphaCSR[ 69 ][ 238 ],
   alphaCSR[ 69 ][ 239 ],
   alphaCSR[ 69 ][ 240 ],
   alphaCSR[ 69 ][ 241 ],
   alphaCSR[ 69 ][ 242 ],
   alphaCSR[ 69 ][ 243 ],
   alphaCSR[ 69 ][ 244 ],
   alphaCSR[ 69 ][ 245 ],
   alphaCSR[ 69 ][ 246 ],
   alphaCSR[ 69 ][ 247 ],
   alphaCSR[ 69 ][ 248 ],
   alphaCSR[ 69 ][ 249 ],
   alphaCSR[ 69 ][ 250 ],
   alphaCSR[ 69 ][ 251 ],
   alphaCSR[ 69 ][ 252 ],
   alphaCSR[ 69 ][ 253 ],
   alphaCSR[ 69 ][ 254 ],
   alphaCSR[ 69 ][ 255 ],
   alphaCSR[ 69 ][ 256 ],
   alphaCSR[ 69 ][ 257 ],
   alphaCSR[ 69 ][ 258 ],
   alphaCSR[ 69 ][ 259 ],
   alphaCSR[ 69 ][ 260 ],
   alphaCSR[ 69 ][ 261 ],
   alphaCSR[ 69 ][ 262 ],
   alphaCSR[ 69 ][ 263 ],
   alphaCSR[ 69 ][ 264 ],
   alphaCSR[ 69 ][ 265 ],
   alphaCSR[ 69 ][ 266 ],
   alphaCSR[ 69 ][ 267 ],
   alphaCSR[ 69 ][ 268 ],
   alphaCSR[ 69 ][ 269 ],
   alphaCSR[ 69 ][ 270 ],
   alphaCSR[ 69 ][ 271 ],
   alphaCSR[ 69 ][ 272 ],
   alphaCSR[ 69 ][ 273 ],
   alphaCSR[ 69 ][ 274 ],
   alphaCSR[ 69 ][ 275 ],
   alphaCSR[ 69 ][ 276 ],
   alphaCSR[ 69 ][ 277 ],
   alphaCSR[ 69 ][ 278 ],
   alphaCSR[ 69 ][ 279 ],
   alphaCSR[ 69 ][ 280 ],
   alphaCSR[ 69 ][ 281 ],
   alphaCSR[ 69 ][ 282 ],
   alphaCSR[ 69 ][ 283 ],
   alphaCSR[ 69 ][ 284 ],
   alphaCSR[ 69 ][ 285 ],
   alphaCSR[ 69 ][ 286 ],
   alphaCSR[ 69 ][ 287 ],
   alphaCSR[ 69 ][ 288 ],
   alphaCSR[ 69 ][ 289 ],
   alphaCSR[ 69 ][ 290 ],
   alphaCSR[ 69 ][ 291 ],
   alphaCSR[ 69 ][ 292 ],
   alphaCSR[ 69 ][ 293 ],
   alphaCSR[ 69 ][ 294 ],
   alphaCSR[ 69 ][ 295 ],
   alphaCSR[ 69 ][ 296 ],
   alphaCSR[ 69 ][ 297 ],
   alphaCSR[ 69 ][ 298 ],
   alphaCSR[ 69 ][ 299 ],
   alphaCSR[ 69 ][ 300 ],
   alphaCSR[ 69 ][ 301 ],
   alphaCSR[ 69 ][ 302 ],
   alphaCSR[ 69 ][ 303 ],
   alphaCSR[ 69 ][ 304 ],
   alphaCSR[ 69 ][ 305 ],
   alphaCSR[ 69 ][ 306 ],
   alphaCSR[ 69 ][ 307 ],
   alphaCSR[ 69 ][ 308 ],
   alphaCSR[ 69 ][ 309 ],
   alphaCSR[ 69 ][ 310 ],
   alphaCSR[ 69 ][ 311 ],
   alphaCSR[ 69 ][ 312 ],
   alphaCSR[ 69 ][ 313 ],
   alphaCSR[ 69 ][ 314 ],
   alphaCSR[ 69 ][ 315 ],
   alphaCSR[ 69 ][ 316 ],
   alphaCSR[ 69 ][ 317 ],
   alphaCSR[ 69 ][ 318 ],
   alphaCSR[ 69 ][ 319 ],
   alphaCSR[ 69 ][ 320 ],
   alphaCSR[ 69 ][ 321 ],
   alphaCSR[ 69 ][ 322 ],
   alphaCSR[ 69 ][ 323 ],
   alphaCSR[ 69 ][ 324 ],
   alphaCSR[ 69 ][ 325 ],
   alphaCSR[ 69 ][ 326 ],
   alphaCSR[ 69 ][ 327 ],
   alphaCSR[ 69 ][ 328 ],
   alphaCSR[ 69 ][ 329 ],
   alphaCSR[ 69 ][ 330 ],
   alphaCSR[ 69 ][ 331 ],
   alphaCSR[ 69 ][ 332 ],
   alphaCSR[ 69 ][ 333 ],
   alphaCSR[ 69 ][ 334 ],
   alphaCSR[ 69 ][ 335 ],
   alphaCSR[ 69 ][ 336 ],
   alphaCSR[ 69 ][ 337 ],
   alphaCSR[ 69 ][ 338 ],
   alphaCSR[ 69 ][ 339 ],
   alphaCSR[ 69 ][ 340 ],
   alphaCSR[ 69 ][ 341 ],
   alphaCSR[ 69 ][ 342 ],
   alphaCSR[ 69 ][ 343 ],
   alphaCSR[ 69 ][ 344 ],
   alphaCSR[ 69 ][ 345 ],
   alphaCSR[ 69 ][ 346 ],
   alphaCSR[ 69 ][ 347 ],
   alphaCSR[ 69 ][ 348 ],
   alphaCSR[ 69 ][ 349 ],
   alphaCSR[ 69 ][ 350 ],
   alphaCSR[ 69 ][ 351 ],
   alphaCSR[ 69 ][ 352 ],
   alphaCSR[ 69 ][ 353 ],
   alphaCSR[ 69 ][ 354 ],
   alphaCSR[ 69 ][ 355 ],
   alphaCSR[ 69 ][ 356 ],
   alphaCSR[ 69 ][ 357 ],
   alphaCSR[ 69 ][ 358 ],
   alphaCSR[ 69 ][ 359 ],
   alphaCSR[ 69 ][ 360 ],
   alphaCSR[ 69 ][ 361 ],
   alphaCSR[ 69 ][ 362 ],
   alphaCSR[ 69 ][ 363 ],
   alphaCSR[ 69 ][ 364 ],
   alphaCSR[ 69 ][ 365 ],
   alphaCSR[ 69 ][ 366 ],
   alphaCSR[ 69 ][ 367 ],
   alphaCSR[ 69 ][ 368 ],
   alphaCSR[ 69 ][ 369 ],
   alphaCSR[ 69 ][ 370 ],
   alphaCSR[ 69 ][ 371 ],
   alphaCSR[ 69 ][ 372 ],
   alphaCSR[ 69 ][ 373 ],
   alphaCSR[ 69 ][ 374 ],
   alphaCSR[ 69 ][ 375 ],
   alphaCSR[ 69 ][ 376 ],
   alphaCSR[ 69 ][ 377 ],
   alphaCSR[ 69 ][ 378 ],
   alphaCSR[ 69 ][ 379 ],
   alphaCSR[ 69 ][ 380 ],
   alphaCSR[ 69 ][ 381 ],
   alphaCSR[ 69 ][ 382 ],
   alphaCSR[ 69 ][ 383 ],
   alphaCSR[ 70 ][ 0 ],
   alphaCSR[ 70 ][ 1 ],
   alphaCSR[ 70 ][ 2 ],
   alphaCSR[ 70 ][ 3 ],
   alphaCSR[ 70 ][ 4 ],
   alphaCSR[ 70 ][ 5 ],
   alphaCSR[ 70 ][ 6 ],
   alphaCSR[ 70 ][ 7 ],
   alphaCSR[ 70 ][ 8 ],
   alphaCSR[ 70 ][ 9 ],
   alphaCSR[ 70 ][ 10 ],
   alphaCSR[ 70 ][ 11 ],
   alphaCSR[ 70 ][ 12 ],
   alphaCSR[ 70 ][ 13 ],
   alphaCSR[ 70 ][ 14 ],
   alphaCSR[ 70 ][ 15 ],
   alphaCSR[ 70 ][ 16 ],
   alphaCSR[ 70 ][ 17 ],
   alphaCSR[ 70 ][ 18 ],
   alphaCSR[ 70 ][ 19 ],
   alphaCSR[ 70 ][ 20 ],
   alphaCSR[ 70 ][ 21 ],
   alphaCSR[ 70 ][ 22 ],
   alphaCSR[ 70 ][ 23 ],
   alphaCSR[ 70 ][ 24 ],
   alphaCSR[ 70 ][ 25 ],
   alphaCSR[ 70 ][ 26 ],
   alphaCSR[ 70 ][ 27 ],
   alphaCSR[ 70 ][ 28 ],
   alphaCSR[ 70 ][ 29 ],
   alphaCSR[ 70 ][ 30 ],
   alphaCSR[ 70 ][ 31 ],
   alphaCSR[ 70 ][ 32 ],
   alphaCSR[ 70 ][ 33 ],
   alphaCSR[ 70 ][ 34 ],
   alphaCSR[ 70 ][ 35 ],
   alphaCSR[ 70 ][ 36 ],
   alphaCSR[ 70 ][ 37 ],
   alphaCSR[ 70 ][ 38 ],
   alphaCSR[ 70 ][ 39 ],
   alphaCSR[ 70 ][ 40 ],
   alphaCSR[ 70 ][ 41 ],
   alphaCSR[ 70 ][ 42 ],
   alphaCSR[ 70 ][ 43 ],
   alphaCSR[ 70 ][ 44 ],
   alphaCSR[ 70 ][ 45 ],
   alphaCSR[ 70 ][ 46 ],
   alphaCSR[ 70 ][ 47 ],
   alphaCSR[ 70 ][ 48 ],
   alphaCSR[ 70 ][ 49 ],
   alphaCSR[ 70 ][ 50 ],
   alphaCSR[ 70 ][ 51 ],
   alphaCSR[ 70 ][ 52 ],
   alphaCSR[ 70 ][ 53 ],
   alphaCSR[ 70 ][ 54 ],
   alphaCSR[ 70 ][ 55 ],
   alphaCSR[ 70 ][ 56 ],
   alphaCSR[ 70 ][ 57 ],
   alphaCSR[ 70 ][ 58 ],
   alphaCSR[ 70 ][ 59 ],
   alphaCSR[ 70 ][ 60 ],
   alphaCSR[ 70 ][ 61 ],
   alphaCSR[ 70 ][ 62 ],
   alphaCSR[ 70 ][ 63 ],
   alphaCSR[ 70 ][ 64 ],
   alphaCSR[ 70 ][ 65 ],
   alphaCSR[ 70 ][ 66 ],
   alphaCSR[ 70 ][ 67 ],
   alphaCSR[ 70 ][ 68 ],
   alphaCSR[ 70 ][ 69 ],
   alphaCSR[ 70 ][ 70 ],
   alphaCSR[ 70 ][ 71 ],
   alphaCSR[ 70 ][ 72 ],
   alphaCSR[ 70 ][ 73 ],
   alphaCSR[ 70 ][ 74 ],
   alphaCSR[ 70 ][ 75 ],
   alphaCSR[ 70 ][ 76 ],
   alphaCSR[ 70 ][ 77 ],
   alphaCSR[ 70 ][ 78 ],
   alphaCSR[ 70 ][ 79 ],
   alphaCSR[ 70 ][ 80 ],
   alphaCSR[ 70 ][ 81 ],
   alphaCSR[ 70 ][ 82 ],
   alphaCSR[ 70 ][ 83 ],
   alphaCSR[ 70 ][ 84 ],
   alphaCSR[ 70 ][ 85 ],
   alphaCSR[ 70 ][ 86 ],
   alphaCSR[ 70 ][ 87 ],
   alphaCSR[ 70 ][ 88 ],
   alphaCSR[ 70 ][ 89 ],
   alphaCSR[ 70 ][ 90 ],
   alphaCSR[ 70 ][ 91 ],
   alphaCSR[ 70 ][ 92 ],
   alphaCSR[ 70 ][ 93 ],
   alphaCSR[ 70 ][ 94 ],
   alphaCSR[ 70 ][ 95 ],
   alphaCSR[ 70 ][ 96 ],
   alphaCSR[ 70 ][ 97 ],
   alphaCSR[ 70 ][ 98 ],
   alphaCSR[ 70 ][ 99 ],
   alphaCSR[ 70 ][ 100 ],
   alphaCSR[ 70 ][ 101 ],
   alphaCSR[ 70 ][ 102 ],
   alphaCSR[ 70 ][ 103 ],
   alphaCSR[ 70 ][ 104 ],
   alphaCSR[ 70 ][ 105 ],
   alphaCSR[ 70 ][ 106 ],
   alphaCSR[ 70 ][ 107 ],
   alphaCSR[ 70 ][ 108 ],
   alphaCSR[ 70 ][ 109 ],
   alphaCSR[ 70 ][ 110 ],
   alphaCSR[ 70 ][ 111 ],
   alphaCSR[ 70 ][ 112 ],
   alphaCSR[ 70 ][ 113 ],
   alphaCSR[ 70 ][ 114 ],
   alphaCSR[ 70 ][ 115 ],
   alphaCSR[ 70 ][ 116 ],
   alphaCSR[ 70 ][ 117 ],
   alphaCSR[ 70 ][ 118 ],
   alphaCSR[ 70 ][ 119 ],
   alphaCSR[ 70 ][ 120 ],
   alphaCSR[ 70 ][ 121 ],
   alphaCSR[ 70 ][ 122 ],
   alphaCSR[ 70 ][ 123 ],
   alphaCSR[ 70 ][ 124 ],
   alphaCSR[ 70 ][ 125 ],
   alphaCSR[ 70 ][ 126 ],
   alphaCSR[ 70 ][ 127 ],
   alphaCSR[ 70 ][ 128 ],
   alphaCSR[ 70 ][ 129 ],
   alphaCSR[ 70 ][ 130 ],
   alphaCSR[ 70 ][ 131 ],
   alphaCSR[ 70 ][ 132 ],
   alphaCSR[ 70 ][ 133 ],
   alphaCSR[ 70 ][ 134 ],
   alphaCSR[ 70 ][ 135 ],
   alphaCSR[ 70 ][ 136 ],
   alphaCSR[ 70 ][ 137 ],
   alphaCSR[ 70 ][ 138 ],
   alphaCSR[ 70 ][ 139 ],
   alphaCSR[ 70 ][ 140 ],
   alphaCSR[ 70 ][ 141 ],
   alphaCSR[ 70 ][ 142 ],
   alphaCSR[ 70 ][ 143 ],
   alphaCSR[ 70 ][ 144 ],
   alphaCSR[ 70 ][ 145 ],
   alphaCSR[ 70 ][ 146 ],
   alphaCSR[ 70 ][ 147 ],
   alphaCSR[ 70 ][ 148 ],
   alphaCSR[ 70 ][ 149 ],
   alphaCSR[ 70 ][ 150 ],
   alphaCSR[ 70 ][ 151 ],
   alphaCSR[ 70 ][ 152 ],
   alphaCSR[ 70 ][ 153 ],
   alphaCSR[ 70 ][ 154 ],
   alphaCSR[ 70 ][ 155 ],
   alphaCSR[ 70 ][ 156 ],
   alphaCSR[ 70 ][ 157 ],
   alphaCSR[ 70 ][ 158 ],
   alphaCSR[ 70 ][ 159 ],
   alphaCSR[ 70 ][ 160 ],
   alphaCSR[ 70 ][ 161 ],
   alphaCSR[ 70 ][ 162 ],
   alphaCSR[ 70 ][ 163 ],
   alphaCSR[ 70 ][ 164 ],
   alphaCSR[ 70 ][ 165 ],
   alphaCSR[ 70 ][ 166 ],
   alphaCSR[ 70 ][ 167 ],
   alphaCSR[ 70 ][ 168 ],
   alphaCSR[ 70 ][ 169 ],
   alphaCSR[ 70 ][ 170 ],
   alphaCSR[ 70 ][ 171 ],
   alphaCSR[ 70 ][ 172 ],
   alphaCSR[ 70 ][ 173 ],
   alphaCSR[ 70 ][ 174 ],
   alphaCSR[ 70 ][ 175 ],
   alphaCSR[ 70 ][ 176 ],
   alphaCSR[ 70 ][ 177 ],
   alphaCSR[ 70 ][ 178 ],
   alphaCSR[ 70 ][ 179 ],
   alphaCSR[ 70 ][ 180 ],
   alphaCSR[ 70 ][ 181 ],
   alphaCSR[ 70 ][ 182 ],
   alphaCSR[ 70 ][ 183 ],
   alphaCSR[ 70 ][ 184 ],
   alphaCSR[ 70 ][ 185 ],
   alphaCSR[ 70 ][ 186 ],
   alphaCSR[ 70 ][ 187 ],
   alphaCSR[ 70 ][ 188 ],
   alphaCSR[ 70 ][ 189 ],
   alphaCSR[ 70 ][ 190 ],
   alphaCSR[ 70 ][ 191 ],
   alphaCSR[ 70 ][ 192 ],
   alphaCSR[ 70 ][ 193 ],
   alphaCSR[ 70 ][ 194 ],
   alphaCSR[ 70 ][ 195 ],
   alphaCSR[ 70 ][ 196 ],
   alphaCSR[ 70 ][ 197 ],
   alphaCSR[ 70 ][ 198 ],
   alphaCSR[ 70 ][ 199 ],
   alphaCSR[ 70 ][ 200 ],
   alphaCSR[ 70 ][ 201 ],
   alphaCSR[ 70 ][ 202 ],
   alphaCSR[ 70 ][ 203 ],
   alphaCSR[ 70 ][ 204 ],
   alphaCSR[ 70 ][ 205 ],
   alphaCSR[ 70 ][ 206 ],
   alphaCSR[ 70 ][ 207 ],
   alphaCSR[ 70 ][ 208 ],
   alphaCSR[ 70 ][ 209 ],
   alphaCSR[ 70 ][ 210 ],
   alphaCSR[ 70 ][ 211 ],
   alphaCSR[ 70 ][ 212 ],
   alphaCSR[ 70 ][ 213 ],
   alphaCSR[ 70 ][ 214 ],
   alphaCSR[ 70 ][ 215 ],
   alphaCSR[ 70 ][ 216 ],
   alphaCSR[ 70 ][ 217 ],
   alphaCSR[ 70 ][ 218 ],
   alphaCSR[ 70 ][ 219 ],
   alphaCSR[ 70 ][ 220 ],
   alphaCSR[ 70 ][ 221 ],
   alphaCSR[ 70 ][ 222 ],
   alphaCSR[ 70 ][ 223 ],
   alphaCSR[ 70 ][ 224 ],
   alphaCSR[ 70 ][ 225 ],
   alphaCSR[ 70 ][ 226 ],
   alphaCSR[ 70 ][ 227 ],
   alphaCSR[ 70 ][ 228 ],
   alphaCSR[ 70 ][ 229 ],
   alphaCSR[ 70 ][ 230 ],
   alphaCSR[ 70 ][ 231 ],
   alphaCSR[ 70 ][ 232 ],
   alphaCSR[ 70 ][ 233 ],
   alphaCSR[ 70 ][ 234 ],
   alphaCSR[ 70 ][ 235 ],
   alphaCSR[ 70 ][ 236 ],
   alphaCSR[ 70 ][ 237 ],
   alphaCSR[ 70 ][ 238 ],
   alphaCSR[ 70 ][ 239 ],
   alphaCSR[ 70 ][ 240 ],
   alphaCSR[ 70 ][ 241 ],
   alphaCSR[ 70 ][ 242 ],
   alphaCSR[ 70 ][ 243 ],
   alphaCSR[ 70 ][ 244 ],
   alphaCSR[ 70 ][ 245 ],
   alphaCSR[ 70 ][ 246 ],
   alphaCSR[ 70 ][ 247 ],
   alphaCSR[ 70 ][ 248 ],
   alphaCSR[ 70 ][ 249 ],
   alphaCSR[ 70 ][ 250 ],
   alphaCSR[ 70 ][ 251 ],
   alphaCSR[ 70 ][ 252 ],
   alphaCSR[ 70 ][ 253 ],
   alphaCSR[ 70 ][ 254 ],
   alphaCSR[ 70 ][ 255 ],
   alphaCSR[ 70 ][ 256 ],
   alphaCSR[ 70 ][ 257 ],
   alphaCSR[ 70 ][ 258 ],
   alphaCSR[ 70 ][ 259 ],
   alphaCSR[ 70 ][ 260 ],
   alphaCSR[ 70 ][ 261 ],
   alphaCSR[ 70 ][ 262 ],
   alphaCSR[ 70 ][ 263 ],
   alphaCSR[ 70 ][ 264 ],
   alphaCSR[ 70 ][ 265 ],
   alphaCSR[ 70 ][ 266 ],
   alphaCSR[ 70 ][ 267 ],
   alphaCSR[ 70 ][ 268 ],
   alphaCSR[ 70 ][ 269 ],
   alphaCSR[ 70 ][ 270 ],
   alphaCSR[ 70 ][ 271 ],
   alphaCSR[ 70 ][ 272 ],
   alphaCSR[ 70 ][ 273 ],
   alphaCSR[ 70 ][ 274 ],
   alphaCSR[ 70 ][ 275 ],
   alphaCSR[ 70 ][ 276 ],
   alphaCSR[ 70 ][ 277 ],
   alphaCSR[ 70 ][ 278 ],
   alphaCSR[ 70 ][ 279 ],
   alphaCSR[ 70 ][ 280 ],
   alphaCSR[ 70 ][ 281 ],
   alphaCSR[ 70 ][ 282 ],
   alphaCSR[ 70 ][ 283 ],
   alphaCSR[ 70 ][ 284 ],
   alphaCSR[ 70 ][ 285 ],
   alphaCSR[ 70 ][ 286 ],
   alphaCSR[ 70 ][ 287 ],
   alphaCSR[ 70 ][ 288 ],
   alphaCSR[ 70 ][ 289 ],
   alphaCSR[ 70 ][ 290 ],
   alphaCSR[ 70 ][ 291 ],
   alphaCSR[ 70 ][ 292 ],
   alphaCSR[ 70 ][ 293 ],
   alphaCSR[ 70 ][ 294 ],
   alphaCSR[ 70 ][ 295 ],
   alphaCSR[ 70 ][ 296 ],
   alphaCSR[ 70 ][ 297 ],
   alphaCSR[ 70 ][ 298 ],
   alphaCSR[ 70 ][ 299 ],
   alphaCSR[ 70 ][ 300 ],
   alphaCSR[ 70 ][ 301 ],
   alphaCSR[ 70 ][ 302 ],
   alphaCSR[ 70 ][ 303 ],
   alphaCSR[ 70 ][ 304 ],
   alphaCSR[ 70 ][ 305 ],
   alphaCSR[ 70 ][ 306 ],
   alphaCSR[ 70 ][ 307 ],
   alphaCSR[ 70 ][ 308 ],
   alphaCSR[ 70 ][ 309 ],
   alphaCSR[ 70 ][ 310 ],
   alphaCSR[ 70 ][ 311 ],
   alphaCSR[ 70 ][ 312 ],
   alphaCSR[ 70 ][ 313 ],
   alphaCSR[ 70 ][ 314 ],
   alphaCSR[ 70 ][ 315 ],
   alphaCSR[ 70 ][ 316 ],
   alphaCSR[ 70 ][ 317 ],
   alphaCSR[ 70 ][ 318 ],
   alphaCSR[ 70 ][ 319 ],
   alphaCSR[ 70 ][ 320 ],
   alphaCSR[ 70 ][ 321 ],
   alphaCSR[ 70 ][ 322 ],
   alphaCSR[ 70 ][ 323 ],
   alphaCSR[ 70 ][ 324 ],
   alphaCSR[ 70 ][ 325 ],
   alphaCSR[ 70 ][ 326 ],
   alphaCSR[ 70 ][ 327 ],
   alphaCSR[ 70 ][ 328 ],
   alphaCSR[ 70 ][ 329 ],
   alphaCSR[ 70 ][ 330 ],
   alphaCSR[ 70 ][ 331 ],
   alphaCSR[ 70 ][ 332 ],
   alphaCSR[ 70 ][ 333 ],
   alphaCSR[ 70 ][ 334 ],
   alphaCSR[ 70 ][ 335 ],
   alphaCSR[ 70 ][ 336 ],
   alphaCSR[ 70 ][ 337 ],
   alphaCSR[ 70 ][ 338 ],
   alphaCSR[ 70 ][ 339 ],
   alphaCSR[ 70 ][ 340 ],
   alphaCSR[ 70 ][ 341 ],
   alphaCSR[ 70 ][ 342 ],
   alphaCSR[ 70 ][ 343 ],
   alphaCSR[ 70 ][ 344 ],
   alphaCSR[ 70 ][ 345 ],
   alphaCSR[ 70 ][ 346 ],
   alphaCSR[ 70 ][ 347 ],
   alphaCSR[ 70 ][ 348 ],
   alphaCSR[ 70 ][ 349 ],
   alphaCSR[ 70 ][ 350 ],
   alphaCSR[ 70 ][ 351 ],
   alphaCSR[ 70 ][ 352 ],
   alphaCSR[ 70 ][ 353 ],
   alphaCSR[ 70 ][ 354 ],
   alphaCSR[ 70 ][ 355 ],
   alphaCSR[ 70 ][ 356 ],
   alphaCSR[ 70 ][ 357 ],
   alphaCSR[ 70 ][ 358 ],
   alphaCSR[ 70 ][ 359 ],
   alphaCSR[ 70 ][ 360 ],
   alphaCSR[ 70 ][ 361 ],
   alphaCSR[ 70 ][ 362 ],
   alphaCSR[ 70 ][ 363 ],
   alphaCSR[ 70 ][ 364 ],
   alphaCSR[ 70 ][ 365 ],
   alphaCSR[ 70 ][ 366 ],
   alphaCSR[ 70 ][ 367 ],
   alphaCSR[ 70 ][ 368 ],
   alphaCSR[ 70 ][ 369 ],
   alphaCSR[ 70 ][ 370 ],
   alphaCSR[ 70 ][ 371 ],
   alphaCSR[ 70 ][ 372 ],
   alphaCSR[ 70 ][ 373 ],
   alphaCSR[ 70 ][ 374 ],
   alphaCSR[ 70 ][ 375 ],
   alphaCSR[ 70 ][ 376 ],
   alphaCSR[ 70 ][ 377 ],
   alphaCSR[ 70 ][ 378 ],
   alphaCSR[ 70 ][ 379 ],
   alphaCSR[ 70 ][ 380 ],
   alphaCSR[ 70 ][ 381 ],
   alphaCSR[ 70 ][ 382 ],
   alphaCSR[ 70 ][ 383 ],
   alphaCSR[ 71 ][ 0 ],
   alphaCSR[ 71 ][ 1 ],
   alphaCSR[ 71 ][ 2 ],
   alphaCSR[ 71 ][ 3 ],
   alphaCSR[ 71 ][ 4 ],
   alphaCSR[ 71 ][ 5 ],
   alphaCSR[ 71 ][ 6 ],
   alphaCSR[ 71 ][ 7 ],
   alphaCSR[ 71 ][ 8 ],
   alphaCSR[ 71 ][ 9 ],
   alphaCSR[ 71 ][ 10 ],
   alphaCSR[ 71 ][ 11 ],
   alphaCSR[ 71 ][ 12 ],
   alphaCSR[ 71 ][ 13 ],
   alphaCSR[ 71 ][ 14 ],
   alphaCSR[ 71 ][ 15 ],
   alphaCSR[ 71 ][ 16 ],
   alphaCSR[ 71 ][ 17 ],
   alphaCSR[ 71 ][ 18 ],
   alphaCSR[ 71 ][ 19 ],
   alphaCSR[ 71 ][ 20 ],
   alphaCSR[ 71 ][ 21 ],
   alphaCSR[ 71 ][ 22 ],
   alphaCSR[ 71 ][ 23 ],
   alphaCSR[ 71 ][ 24 ],
   alphaCSR[ 71 ][ 25 ],
   alphaCSR[ 71 ][ 26 ],
   alphaCSR[ 71 ][ 27 ],
   alphaCSR[ 71 ][ 28 ],
   alphaCSR[ 71 ][ 29 ],
   alphaCSR[ 71 ][ 30 ],
   alphaCSR[ 71 ][ 31 ],
   alphaCSR[ 71 ][ 32 ],
   alphaCSR[ 71 ][ 33 ],
   alphaCSR[ 71 ][ 34 ],
   alphaCSR[ 71 ][ 35 ],
   alphaCSR[ 71 ][ 36 ],
   alphaCSR[ 71 ][ 37 ],
   alphaCSR[ 71 ][ 38 ],
   alphaCSR[ 71 ][ 39 ],
   alphaCSR[ 71 ][ 40 ],
   alphaCSR[ 71 ][ 41 ],
   alphaCSR[ 71 ][ 42 ],
   alphaCSR[ 71 ][ 43 ],
   alphaCSR[ 71 ][ 44 ],
   alphaCSR[ 71 ][ 45 ],
   alphaCSR[ 71 ][ 46 ],
   alphaCSR[ 71 ][ 47 ],
   alphaCSR[ 71 ][ 48 ],
   alphaCSR[ 71 ][ 49 ],
   alphaCSR[ 71 ][ 50 ],
   alphaCSR[ 71 ][ 51 ],
   alphaCSR[ 71 ][ 52 ],
   alphaCSR[ 71 ][ 53 ],
   alphaCSR[ 71 ][ 54 ],
   alphaCSR[ 71 ][ 55 ],
   alphaCSR[ 71 ][ 56 ],
   alphaCSR[ 71 ][ 57 ],
   alphaCSR[ 71 ][ 58 ],
   alphaCSR[ 71 ][ 59 ],
   alphaCSR[ 71 ][ 60 ],
   alphaCSR[ 71 ][ 61 ],
   alphaCSR[ 71 ][ 62 ],
   alphaCSR[ 71 ][ 63 ],
   alphaCSR[ 71 ][ 64 ],
   alphaCSR[ 71 ][ 65 ],
   alphaCSR[ 71 ][ 66 ],
   alphaCSR[ 71 ][ 67 ],
   alphaCSR[ 71 ][ 68 ],
   alphaCSR[ 71 ][ 69 ],
   alphaCSR[ 71 ][ 70 ],
   alphaCSR[ 71 ][ 71 ],
   alphaCSR[ 71 ][ 72 ],
   alphaCSR[ 71 ][ 73 ],
   alphaCSR[ 71 ][ 74 ],
   alphaCSR[ 71 ][ 75 ],
   alphaCSR[ 71 ][ 76 ],
   alphaCSR[ 71 ][ 77 ],
   alphaCSR[ 71 ][ 78 ],
   alphaCSR[ 71 ][ 79 ],
   alphaCSR[ 71 ][ 80 ],
   alphaCSR[ 71 ][ 81 ],
   alphaCSR[ 71 ][ 82 ],
   alphaCSR[ 71 ][ 83 ],
   alphaCSR[ 71 ][ 84 ],
   alphaCSR[ 71 ][ 85 ],
   alphaCSR[ 71 ][ 86 ],
   alphaCSR[ 71 ][ 87 ],
   alphaCSR[ 71 ][ 88 ],
   alphaCSR[ 71 ][ 89 ],
   alphaCSR[ 71 ][ 90 ],
   alphaCSR[ 71 ][ 91 ],
   alphaCSR[ 71 ][ 92 ],
   alphaCSR[ 71 ][ 93 ],
   alphaCSR[ 71 ][ 94 ],
   alphaCSR[ 71 ][ 95 ],
   alphaCSR[ 71 ][ 96 ],
   alphaCSR[ 71 ][ 97 ],
   alphaCSR[ 71 ][ 98 ],
   alphaCSR[ 71 ][ 99 ],
   alphaCSR[ 71 ][ 100 ],
   alphaCSR[ 71 ][ 101 ],
   alphaCSR[ 71 ][ 102 ],
   alphaCSR[ 71 ][ 103 ],
   alphaCSR[ 71 ][ 104 ],
   alphaCSR[ 71 ][ 105 ],
   alphaCSR[ 71 ][ 106 ],
   alphaCSR[ 71 ][ 107 ],
   alphaCSR[ 71 ][ 108 ],
   alphaCSR[ 71 ][ 109 ],
   alphaCSR[ 71 ][ 110 ],
   alphaCSR[ 71 ][ 111 ],
   alphaCSR[ 71 ][ 112 ],
   alphaCSR[ 71 ][ 113 ],
   alphaCSR[ 71 ][ 114 ],
   alphaCSR[ 71 ][ 115 ],
   alphaCSR[ 71 ][ 116 ],
   alphaCSR[ 71 ][ 117 ],
   alphaCSR[ 71 ][ 118 ],
   alphaCSR[ 71 ][ 119 ],
   alphaCSR[ 71 ][ 120 ],
   alphaCSR[ 71 ][ 121 ],
   alphaCSR[ 71 ][ 122 ],
   alphaCSR[ 71 ][ 123 ],
   alphaCSR[ 71 ][ 124 ],
   alphaCSR[ 71 ][ 125 ],
   alphaCSR[ 71 ][ 126 ],
   alphaCSR[ 71 ][ 127 ],
   alphaCSR[ 71 ][ 128 ],
   alphaCSR[ 71 ][ 129 ],
   alphaCSR[ 71 ][ 130 ],
   alphaCSR[ 71 ][ 131 ],
   alphaCSR[ 71 ][ 132 ],
   alphaCSR[ 71 ][ 133 ],
   alphaCSR[ 71 ][ 134 ],
   alphaCSR[ 71 ][ 135 ],
   alphaCSR[ 71 ][ 136 ],
   alphaCSR[ 71 ][ 137 ],
   alphaCSR[ 71 ][ 138 ],
   alphaCSR[ 71 ][ 139 ],
   alphaCSR[ 71 ][ 140 ],
   alphaCSR[ 71 ][ 141 ],
   alphaCSR[ 71 ][ 142 ],
   alphaCSR[ 71 ][ 143 ],
   alphaCSR[ 71 ][ 144 ],
   alphaCSR[ 71 ][ 145 ],
   alphaCSR[ 71 ][ 146 ],
   alphaCSR[ 71 ][ 147 ],
   alphaCSR[ 71 ][ 148 ],
   alphaCSR[ 71 ][ 149 ],
   alphaCSR[ 71 ][ 150 ],
   alphaCSR[ 71 ][ 151 ],
   alphaCSR[ 71 ][ 152 ],
   alphaCSR[ 71 ][ 153 ],
   alphaCSR[ 71 ][ 154 ],
   alphaCSR[ 71 ][ 155 ],
   alphaCSR[ 71 ][ 156 ],
   alphaCSR[ 71 ][ 157 ],
   alphaCSR[ 71 ][ 158 ],
   alphaCSR[ 71 ][ 159 ],
   alphaCSR[ 71 ][ 160 ],
   alphaCSR[ 71 ][ 161 ],
   alphaCSR[ 71 ][ 162 ],
   alphaCSR[ 71 ][ 163 ],
   alphaCSR[ 71 ][ 164 ],
   alphaCSR[ 71 ][ 165 ],
   alphaCSR[ 71 ][ 166 ],
   alphaCSR[ 71 ][ 167 ],
   alphaCSR[ 71 ][ 168 ],
   alphaCSR[ 71 ][ 169 ],
   alphaCSR[ 71 ][ 170 ],
   alphaCSR[ 71 ][ 171 ],
   alphaCSR[ 71 ][ 172 ],
   alphaCSR[ 71 ][ 173 ],
   alphaCSR[ 71 ][ 174 ],
   alphaCSR[ 71 ][ 175 ],
   alphaCSR[ 71 ][ 176 ],
   alphaCSR[ 71 ][ 177 ],
   alphaCSR[ 71 ][ 178 ],
   alphaCSR[ 71 ][ 179 ],
   alphaCSR[ 71 ][ 180 ],
   alphaCSR[ 71 ][ 181 ],
   alphaCSR[ 71 ][ 182 ],
   alphaCSR[ 71 ][ 183 ],
   alphaCSR[ 71 ][ 184 ],
   alphaCSR[ 71 ][ 185 ],
   alphaCSR[ 71 ][ 186 ],
   alphaCSR[ 71 ][ 187 ],
   alphaCSR[ 71 ][ 188 ],
   alphaCSR[ 71 ][ 189 ],
   alphaCSR[ 71 ][ 190 ],
   alphaCSR[ 71 ][ 191 ],
   alphaCSR[ 71 ][ 192 ],
   alphaCSR[ 71 ][ 193 ],
   alphaCSR[ 71 ][ 194 ],
   alphaCSR[ 71 ][ 195 ],
   alphaCSR[ 71 ][ 196 ],
   alphaCSR[ 71 ][ 197 ],
   alphaCSR[ 71 ][ 198 ],
   alphaCSR[ 71 ][ 199 ],
   alphaCSR[ 71 ][ 200 ],
   alphaCSR[ 71 ][ 201 ],
   alphaCSR[ 71 ][ 202 ],
   alphaCSR[ 71 ][ 203 ],
   alphaCSR[ 71 ][ 204 ],
   alphaCSR[ 71 ][ 205 ],
   alphaCSR[ 71 ][ 206 ],
   alphaCSR[ 71 ][ 207 ],
   alphaCSR[ 71 ][ 208 ],
   alphaCSR[ 71 ][ 209 ],
   alphaCSR[ 71 ][ 210 ],
   alphaCSR[ 71 ][ 211 ],
   alphaCSR[ 71 ][ 212 ],
   alphaCSR[ 71 ][ 213 ],
   alphaCSR[ 71 ][ 214 ],
   alphaCSR[ 71 ][ 215 ],
   alphaCSR[ 71 ][ 216 ],
   alphaCSR[ 71 ][ 217 ],
   alphaCSR[ 71 ][ 218 ],
   alphaCSR[ 71 ][ 219 ],
   alphaCSR[ 71 ][ 220 ],
   alphaCSR[ 71 ][ 221 ],
   alphaCSR[ 71 ][ 222 ],
   alphaCSR[ 71 ][ 223 ],
   alphaCSR[ 71 ][ 224 ],
   alphaCSR[ 71 ][ 225 ],
   alphaCSR[ 71 ][ 226 ],
   alphaCSR[ 71 ][ 227 ],
   alphaCSR[ 71 ][ 228 ],
   alphaCSR[ 71 ][ 229 ],
   alphaCSR[ 71 ][ 230 ],
   alphaCSR[ 71 ][ 231 ],
   alphaCSR[ 71 ][ 232 ],
   alphaCSR[ 71 ][ 233 ],
   alphaCSR[ 71 ][ 234 ],
   alphaCSR[ 71 ][ 235 ],
   alphaCSR[ 71 ][ 236 ],
   alphaCSR[ 71 ][ 237 ],
   alphaCSR[ 71 ][ 238 ],
   alphaCSR[ 71 ][ 239 ],
   alphaCSR[ 71 ][ 240 ],
   alphaCSR[ 71 ][ 241 ],
   alphaCSR[ 71 ][ 242 ],
   alphaCSR[ 71 ][ 243 ],
   alphaCSR[ 71 ][ 244 ],
   alphaCSR[ 71 ][ 245 ],
   alphaCSR[ 71 ][ 246 ],
   alphaCSR[ 71 ][ 247 ],
   alphaCSR[ 71 ][ 248 ],
   alphaCSR[ 71 ][ 249 ],
   alphaCSR[ 71 ][ 250 ],
   alphaCSR[ 71 ][ 251 ],
   alphaCSR[ 71 ][ 252 ],
   alphaCSR[ 71 ][ 253 ],
   alphaCSR[ 71 ][ 254 ],
   alphaCSR[ 71 ][ 255 ],
   alphaCSR[ 71 ][ 256 ],
   alphaCSR[ 71 ][ 257 ],
   alphaCSR[ 71 ][ 258 ],
   alphaCSR[ 71 ][ 259 ],
   alphaCSR[ 71 ][ 260 ],
   alphaCSR[ 71 ][ 261 ],
   alphaCSR[ 71 ][ 262 ],
   alphaCSR[ 71 ][ 263 ],
   alphaCSR[ 71 ][ 264 ],
   alphaCSR[ 71 ][ 265 ],
   alphaCSR[ 71 ][ 266 ],
   alphaCSR[ 71 ][ 267 ],
   alphaCSR[ 71 ][ 268 ],
   alphaCSR[ 71 ][ 269 ],
   alphaCSR[ 71 ][ 270 ],
   alphaCSR[ 71 ][ 271 ],
   alphaCSR[ 71 ][ 272 ],
   alphaCSR[ 71 ][ 273 ],
   alphaCSR[ 71 ][ 274 ],
   alphaCSR[ 71 ][ 275 ],
   alphaCSR[ 71 ][ 276 ],
   alphaCSR[ 71 ][ 277 ],
   alphaCSR[ 71 ][ 278 ],
   alphaCSR[ 71 ][ 279 ],
   alphaCSR[ 71 ][ 280 ],
   alphaCSR[ 71 ][ 281 ],
   alphaCSR[ 71 ][ 282 ],
   alphaCSR[ 71 ][ 283 ],
   alphaCSR[ 71 ][ 284 ],
   alphaCSR[ 71 ][ 285 ],
   alphaCSR[ 71 ][ 286 ],
   alphaCSR[ 71 ][ 287 ],
   alphaCSR[ 71 ][ 288 ],
   alphaCSR[ 71 ][ 289 ],
   alphaCSR[ 71 ][ 290 ],
   alphaCSR[ 71 ][ 291 ],
   alphaCSR[ 71 ][ 292 ],
   alphaCSR[ 71 ][ 293 ],
   alphaCSR[ 71 ][ 294 ],
   alphaCSR[ 71 ][ 295 ],
   alphaCSR[ 71 ][ 296 ],
   alphaCSR[ 71 ][ 297 ],
   alphaCSR[ 71 ][ 298 ],
   alphaCSR[ 71 ][ 299 ],
   alphaCSR[ 71 ][ 300 ],
   alphaCSR[ 71 ][ 301 ],
   alphaCSR[ 71 ][ 302 ],
   alphaCSR[ 71 ][ 303 ],
   alphaCSR[ 71 ][ 304 ],
   alphaCSR[ 71 ][ 305 ],
   alphaCSR[ 71 ][ 306 ],
   alphaCSR[ 71 ][ 307 ],
   alphaCSR[ 71 ][ 308 ],
   alphaCSR[ 71 ][ 309 ],
   alphaCSR[ 71 ][ 310 ],
   alphaCSR[ 71 ][ 311 ],
   alphaCSR[ 71 ][ 312 ],
   alphaCSR[ 71 ][ 313 ],
   alphaCSR[ 71 ][ 314 ],
   alphaCSR[ 71 ][ 315 ],
   alphaCSR[ 71 ][ 316 ],
   alphaCSR[ 71 ][ 317 ],
   alphaCSR[ 71 ][ 318 ],
   alphaCSR[ 71 ][ 319 ],
   alphaCSR[ 71 ][ 320 ],
   alphaCSR[ 71 ][ 321 ],
   alphaCSR[ 71 ][ 322 ],
   alphaCSR[ 71 ][ 323 ],
   alphaCSR[ 71 ][ 324 ],
   alphaCSR[ 71 ][ 325 ],
   alphaCSR[ 71 ][ 326 ],
   alphaCSR[ 71 ][ 327 ],
   alphaCSR[ 71 ][ 328 ],
   alphaCSR[ 71 ][ 329 ],
   alphaCSR[ 71 ][ 330 ],
   alphaCSR[ 71 ][ 331 ],
   alphaCSR[ 71 ][ 332 ],
   alphaCSR[ 71 ][ 333 ],
   alphaCSR[ 71 ][ 334 ],
   alphaCSR[ 71 ][ 335 ],
   alphaCSR[ 71 ][ 336 ],
   alphaCSR[ 71 ][ 337 ],
   alphaCSR[ 71 ][ 338 ],
   alphaCSR[ 71 ][ 339 ],
   alphaCSR[ 71 ][ 340 ],
   alphaCSR[ 71 ][ 341 ],
   alphaCSR[ 71 ][ 342 ],
   alphaCSR[ 71 ][ 343 ],
   alphaCSR[ 71 ][ 344 ],
   alphaCSR[ 71 ][ 345 ],
   alphaCSR[ 71 ][ 346 ],
   alphaCSR[ 71 ][ 347 ],
   alphaCSR[ 71 ][ 348 ],
   alphaCSR[ 71 ][ 349 ],
   alphaCSR[ 71 ][ 350 ],
   alphaCSR[ 71 ][ 351 ],
   alphaCSR[ 71 ][ 352 ],
   alphaCSR[ 71 ][ 353 ],
   alphaCSR[ 71 ][ 354 ],
   alphaCSR[ 71 ][ 355 ],
   alphaCSR[ 71 ][ 356 ],
   alphaCSR[ 71 ][ 357 ],
   alphaCSR[ 71 ][ 358 ],
   alphaCSR[ 71 ][ 359 ],
   alphaCSR[ 71 ][ 360 ],
   alphaCSR[ 71 ][ 361 ],
   alphaCSR[ 71 ][ 362 ],
   alphaCSR[ 71 ][ 363 ],
   alphaCSR[ 71 ][ 364 ],
   alphaCSR[ 71 ][ 365 ],
   alphaCSR[ 71 ][ 366 ],
   alphaCSR[ 71 ][ 367 ],
   alphaCSR[ 71 ][ 368 ],
   alphaCSR[ 71 ][ 369 ],
   alphaCSR[ 71 ][ 370 ],
   alphaCSR[ 71 ][ 371 ],
   alphaCSR[ 71 ][ 372 ],
   alphaCSR[ 71 ][ 373 ],
   alphaCSR[ 71 ][ 374 ],
   alphaCSR[ 71 ][ 375 ],
   alphaCSR[ 71 ][ 376 ],
   alphaCSR[ 71 ][ 377 ],
   alphaCSR[ 71 ][ 378 ],
   alphaCSR[ 71 ][ 379 ],
   alphaCSR[ 71 ][ 380 ],
   alphaCSR[ 71 ][ 381 ],
   alphaCSR[ 71 ][ 382 ],
   alphaCSR[ 71 ][ 383 ],
   alphaCSR[ 72 ][ 0 ],
   alphaCSR[ 72 ][ 1 ],
   alphaCSR[ 72 ][ 2 ],
   alphaCSR[ 72 ][ 3 ],
   alphaCSR[ 72 ][ 4 ],
   alphaCSR[ 72 ][ 5 ],
   alphaCSR[ 72 ][ 6 ],
   alphaCSR[ 72 ][ 7 ],
   alphaCSR[ 72 ][ 8 ],
   alphaCSR[ 72 ][ 9 ],
   alphaCSR[ 72 ][ 10 ],
   alphaCSR[ 72 ][ 11 ],
   alphaCSR[ 72 ][ 12 ],
   alphaCSR[ 72 ][ 13 ],
   alphaCSR[ 72 ][ 14 ],
   alphaCSR[ 72 ][ 15 ],
   alphaCSR[ 72 ][ 16 ],
   alphaCSR[ 72 ][ 17 ],
   alphaCSR[ 72 ][ 18 ],
   alphaCSR[ 72 ][ 19 ],
   alphaCSR[ 72 ][ 20 ],
   alphaCSR[ 72 ][ 21 ],
   alphaCSR[ 72 ][ 22 ],
   alphaCSR[ 72 ][ 23 ],
   alphaCSR[ 72 ][ 24 ],
   alphaCSR[ 72 ][ 25 ],
   alphaCSR[ 72 ][ 26 ],
   alphaCSR[ 72 ][ 27 ],
   alphaCSR[ 72 ][ 28 ],
   alphaCSR[ 72 ][ 29 ],
   alphaCSR[ 72 ][ 30 ],
   alphaCSR[ 72 ][ 31 ],
   alphaCSR[ 72 ][ 32 ],
   alphaCSR[ 72 ][ 33 ],
   alphaCSR[ 72 ][ 34 ],
   alphaCSR[ 72 ][ 35 ],
   alphaCSR[ 72 ][ 36 ],
   alphaCSR[ 72 ][ 37 ],
   alphaCSR[ 72 ][ 38 ],
   alphaCSR[ 72 ][ 39 ],
   alphaCSR[ 72 ][ 40 ],
   alphaCSR[ 72 ][ 41 ],
   alphaCSR[ 72 ][ 42 ],
   alphaCSR[ 72 ][ 43 ],
   alphaCSR[ 72 ][ 44 ],
   alphaCSR[ 72 ][ 45 ],
   alphaCSR[ 72 ][ 46 ],
   alphaCSR[ 72 ][ 47 ],
   alphaCSR[ 72 ][ 48 ],
   alphaCSR[ 72 ][ 49 ],
   alphaCSR[ 72 ][ 50 ],
   alphaCSR[ 72 ][ 51 ],
   alphaCSR[ 72 ][ 52 ],
   alphaCSR[ 72 ][ 53 ],
   alphaCSR[ 72 ][ 54 ],
   alphaCSR[ 72 ][ 55 ],
   alphaCSR[ 72 ][ 56 ],
   alphaCSR[ 72 ][ 57 ],
   alphaCSR[ 72 ][ 58 ],
   alphaCSR[ 72 ][ 59 ],
   alphaCSR[ 72 ][ 60 ],
   alphaCSR[ 72 ][ 61 ],
   alphaCSR[ 72 ][ 62 ],
   alphaCSR[ 72 ][ 63 ],
   alphaCSR[ 72 ][ 64 ],
   alphaCSR[ 72 ][ 65 ],
   alphaCSR[ 72 ][ 66 ],
   alphaCSR[ 72 ][ 67 ],
   alphaCSR[ 72 ][ 68 ],
   alphaCSR[ 72 ][ 69 ],
   alphaCSR[ 72 ][ 70 ],
   alphaCSR[ 72 ][ 71 ],
   alphaCSR[ 72 ][ 72 ],
   alphaCSR[ 72 ][ 73 ],
   alphaCSR[ 72 ][ 74 ],
   alphaCSR[ 72 ][ 75 ],
   alphaCSR[ 72 ][ 76 ],
   alphaCSR[ 72 ][ 77 ],
   alphaCSR[ 72 ][ 78 ],
   alphaCSR[ 72 ][ 79 ],
   alphaCSR[ 72 ][ 80 ],
   alphaCSR[ 72 ][ 81 ],
   alphaCSR[ 72 ][ 82 ],
   alphaCSR[ 72 ][ 83 ],
   alphaCSR[ 72 ][ 84 ],
   alphaCSR[ 72 ][ 85 ],
   alphaCSR[ 72 ][ 86 ],
   alphaCSR[ 72 ][ 87 ],
   alphaCSR[ 72 ][ 88 ],
   alphaCSR[ 72 ][ 89 ],
   alphaCSR[ 72 ][ 90 ],
   alphaCSR[ 72 ][ 91 ],
   alphaCSR[ 72 ][ 92 ],
   alphaCSR[ 72 ][ 93 ],
   alphaCSR[ 72 ][ 94 ],
   alphaCSR[ 72 ][ 95 ],
   alphaCSR[ 72 ][ 96 ],
   alphaCSR[ 72 ][ 97 ],
   alphaCSR[ 72 ][ 98 ],
   alphaCSR[ 72 ][ 99 ],
   alphaCSR[ 72 ][ 100 ],
   alphaCSR[ 72 ][ 101 ],
   alphaCSR[ 72 ][ 102 ],
   alphaCSR[ 72 ][ 103 ],
   alphaCSR[ 72 ][ 104 ],
   alphaCSR[ 72 ][ 105 ],
   alphaCSR[ 72 ][ 106 ],
   alphaCSR[ 72 ][ 107 ],
   alphaCSR[ 72 ][ 108 ],
   alphaCSR[ 72 ][ 109 ],
   alphaCSR[ 72 ][ 110 ],
   alphaCSR[ 72 ][ 111 ],
   alphaCSR[ 72 ][ 112 ],
   alphaCSR[ 72 ][ 113 ],
   alphaCSR[ 72 ][ 114 ],
   alphaCSR[ 72 ][ 115 ],
   alphaCSR[ 72 ][ 116 ],
   alphaCSR[ 72 ][ 117 ],
   alphaCSR[ 72 ][ 118 ],
   alphaCSR[ 72 ][ 119 ],
   alphaCSR[ 72 ][ 120 ],
   alphaCSR[ 72 ][ 121 ],
   alphaCSR[ 72 ][ 122 ],
   alphaCSR[ 72 ][ 123 ],
   alphaCSR[ 72 ][ 124 ],
   alphaCSR[ 72 ][ 125 ],
   alphaCSR[ 72 ][ 126 ],
   alphaCSR[ 72 ][ 127 ],
   alphaCSR[ 72 ][ 128 ],
   alphaCSR[ 72 ][ 129 ],
   alphaCSR[ 72 ][ 130 ],
   alphaCSR[ 72 ][ 131 ],
   alphaCSR[ 72 ][ 132 ],
   alphaCSR[ 72 ][ 133 ],
   alphaCSR[ 72 ][ 134 ],
   alphaCSR[ 72 ][ 135 ],
   alphaCSR[ 72 ][ 136 ],
   alphaCSR[ 72 ][ 137 ],
   alphaCSR[ 72 ][ 138 ],
   alphaCSR[ 72 ][ 139 ],
   alphaCSR[ 72 ][ 140 ],
   alphaCSR[ 72 ][ 141 ],
   alphaCSR[ 72 ][ 142 ],
   alphaCSR[ 72 ][ 143 ],
   alphaCSR[ 72 ][ 144 ],
   alphaCSR[ 72 ][ 145 ],
   alphaCSR[ 72 ][ 146 ],
   alphaCSR[ 72 ][ 147 ],
   alphaCSR[ 72 ][ 148 ],
   alphaCSR[ 72 ][ 149 ],
   alphaCSR[ 72 ][ 150 ],
   alphaCSR[ 72 ][ 151 ],
   alphaCSR[ 72 ][ 152 ],
   alphaCSR[ 72 ][ 153 ],
   alphaCSR[ 72 ][ 154 ],
   alphaCSR[ 72 ][ 155 ],
   alphaCSR[ 72 ][ 156 ],
   alphaCSR[ 72 ][ 157 ],
   alphaCSR[ 72 ][ 158 ],
   alphaCSR[ 72 ][ 159 ],
   alphaCSR[ 72 ][ 160 ],
   alphaCSR[ 72 ][ 161 ],
   alphaCSR[ 72 ][ 162 ],
   alphaCSR[ 72 ][ 163 ],
   alphaCSR[ 72 ][ 164 ],
   alphaCSR[ 72 ][ 165 ],
   alphaCSR[ 72 ][ 166 ],
   alphaCSR[ 72 ][ 167 ],
   alphaCSR[ 72 ][ 168 ],
   alphaCSR[ 72 ][ 169 ],
   alphaCSR[ 72 ][ 170 ],
   alphaCSR[ 72 ][ 171 ],
   alphaCSR[ 72 ][ 172 ],
   alphaCSR[ 72 ][ 173 ],
   alphaCSR[ 72 ][ 174 ],
   alphaCSR[ 72 ][ 175 ],
   alphaCSR[ 72 ][ 176 ],
   alphaCSR[ 72 ][ 177 ],
   alphaCSR[ 72 ][ 178 ],
   alphaCSR[ 72 ][ 179 ],
   alphaCSR[ 72 ][ 180 ],
   alphaCSR[ 72 ][ 181 ],
   alphaCSR[ 72 ][ 182 ],
   alphaCSR[ 72 ][ 183 ],
   alphaCSR[ 72 ][ 184 ],
   alphaCSR[ 72 ][ 185 ],
   alphaCSR[ 72 ][ 186 ],
   alphaCSR[ 72 ][ 187 ],
   alphaCSR[ 72 ][ 188 ],
   alphaCSR[ 72 ][ 189 ],
   alphaCSR[ 72 ][ 190 ],
   alphaCSR[ 72 ][ 191 ],
   alphaCSR[ 72 ][ 192 ],
   alphaCSR[ 72 ][ 193 ],
   alphaCSR[ 72 ][ 194 ],
   alphaCSR[ 72 ][ 195 ],
   alphaCSR[ 72 ][ 196 ],
   alphaCSR[ 72 ][ 197 ],
   alphaCSR[ 72 ][ 198 ],
   alphaCSR[ 72 ][ 199 ],
   alphaCSR[ 72 ][ 200 ],
   alphaCSR[ 72 ][ 201 ],
   alphaCSR[ 72 ][ 202 ],
   alphaCSR[ 72 ][ 203 ],
   alphaCSR[ 72 ][ 204 ],
   alphaCSR[ 72 ][ 205 ],
   alphaCSR[ 72 ][ 206 ],
   alphaCSR[ 72 ][ 207 ],
   alphaCSR[ 72 ][ 208 ],
   alphaCSR[ 72 ][ 209 ],
   alphaCSR[ 72 ][ 210 ],
   alphaCSR[ 72 ][ 211 ],
   alphaCSR[ 72 ][ 212 ],
   alphaCSR[ 72 ][ 213 ],
   alphaCSR[ 72 ][ 214 ],
   alphaCSR[ 72 ][ 215 ],
   alphaCSR[ 72 ][ 216 ],
   alphaCSR[ 72 ][ 217 ],
   alphaCSR[ 72 ][ 218 ],
   alphaCSR[ 72 ][ 219 ],
   alphaCSR[ 72 ][ 220 ],
   alphaCSR[ 72 ][ 221 ],
   alphaCSR[ 72 ][ 222 ],
   alphaCSR[ 72 ][ 223 ],
   alphaCSR[ 72 ][ 224 ],
   alphaCSR[ 72 ][ 225 ],
   alphaCSR[ 72 ][ 226 ],
   alphaCSR[ 72 ][ 227 ],
   alphaCSR[ 72 ][ 228 ],
   alphaCSR[ 72 ][ 229 ],
   alphaCSR[ 72 ][ 230 ],
   alphaCSR[ 72 ][ 231 ],
   alphaCSR[ 72 ][ 232 ],
   alphaCSR[ 72 ][ 233 ],
   alphaCSR[ 72 ][ 234 ],
   alphaCSR[ 72 ][ 235 ],
   alphaCSR[ 72 ][ 236 ],
   alphaCSR[ 72 ][ 237 ],
   alphaCSR[ 72 ][ 238 ],
   alphaCSR[ 72 ][ 239 ],
   alphaCSR[ 72 ][ 240 ],
   alphaCSR[ 72 ][ 241 ],
   alphaCSR[ 72 ][ 242 ],
   alphaCSR[ 72 ][ 243 ],
   alphaCSR[ 72 ][ 244 ],
   alphaCSR[ 72 ][ 245 ],
   alphaCSR[ 72 ][ 246 ],
   alphaCSR[ 72 ][ 247 ],
   alphaCSR[ 72 ][ 248 ],
   alphaCSR[ 72 ][ 249 ],
   alphaCSR[ 72 ][ 250 ],
   alphaCSR[ 72 ][ 251 ],
   alphaCSR[ 72 ][ 252 ],
   alphaCSR[ 72 ][ 253 ],
   alphaCSR[ 72 ][ 254 ],
   alphaCSR[ 72 ][ 255 ],
   alphaCSR[ 72 ][ 256 ],
   alphaCSR[ 72 ][ 257 ],
   alphaCSR[ 72 ][ 258 ],
   alphaCSR[ 72 ][ 259 ],
   alphaCSR[ 72 ][ 260 ],
   alphaCSR[ 72 ][ 261 ],
   alphaCSR[ 72 ][ 262 ],
   alphaCSR[ 72 ][ 263 ],
   alphaCSR[ 72 ][ 264 ],
   alphaCSR[ 72 ][ 265 ],
   alphaCSR[ 72 ][ 266 ],
   alphaCSR[ 72 ][ 267 ],
   alphaCSR[ 72 ][ 268 ],
   alphaCSR[ 72 ][ 269 ],
   alphaCSR[ 72 ][ 270 ],
   alphaCSR[ 72 ][ 271 ],
   alphaCSR[ 72 ][ 272 ],
   alphaCSR[ 72 ][ 273 ],
   alphaCSR[ 72 ][ 274 ],
   alphaCSR[ 72 ][ 275 ],
   alphaCSR[ 72 ][ 276 ],
   alphaCSR[ 72 ][ 277 ],
   alphaCSR[ 72 ][ 278 ],
   alphaCSR[ 72 ][ 279 ],
   alphaCSR[ 72 ][ 280 ],
   alphaCSR[ 72 ][ 281 ],
   alphaCSR[ 72 ][ 282 ],
   alphaCSR[ 72 ][ 283 ],
   alphaCSR[ 72 ][ 284 ],
   alphaCSR[ 72 ][ 285 ],
   alphaCSR[ 72 ][ 286 ],
   alphaCSR[ 72 ][ 287 ],
   alphaCSR[ 72 ][ 288 ],
   alphaCSR[ 72 ][ 289 ],
   alphaCSR[ 72 ][ 290 ],
   alphaCSR[ 72 ][ 291 ],
   alphaCSR[ 72 ][ 292 ],
   alphaCSR[ 72 ][ 293 ],
   alphaCSR[ 72 ][ 294 ],
   alphaCSR[ 72 ][ 295 ],
   alphaCSR[ 72 ][ 296 ],
   alphaCSR[ 72 ][ 297 ],
   alphaCSR[ 72 ][ 298 ],
   alphaCSR[ 72 ][ 299 ],
   alphaCSR[ 72 ][ 300 ],
   alphaCSR[ 72 ][ 301 ],
   alphaCSR[ 72 ][ 302 ],
   alphaCSR[ 72 ][ 303 ],
   alphaCSR[ 72 ][ 304 ],
   alphaCSR[ 72 ][ 305 ],
   alphaCSR[ 72 ][ 306 ],
   alphaCSR[ 72 ][ 307 ],
   alphaCSR[ 72 ][ 308 ],
   alphaCSR[ 72 ][ 309 ],
   alphaCSR[ 72 ][ 310 ],
   alphaCSR[ 72 ][ 311 ],
   alphaCSR[ 72 ][ 312 ],
   alphaCSR[ 72 ][ 313 ],
   alphaCSR[ 72 ][ 314 ],
   alphaCSR[ 72 ][ 315 ],
   alphaCSR[ 72 ][ 316 ],
   alphaCSR[ 72 ][ 317 ],
   alphaCSR[ 72 ][ 318 ],
   alphaCSR[ 72 ][ 319 ],
   alphaCSR[ 72 ][ 320 ],
   alphaCSR[ 72 ][ 321 ],
   alphaCSR[ 72 ][ 322 ],
   alphaCSR[ 72 ][ 323 ],
   alphaCSR[ 72 ][ 324 ],
   alphaCSR[ 72 ][ 325 ],
   alphaCSR[ 72 ][ 326 ],
   alphaCSR[ 72 ][ 327 ],
   alphaCSR[ 72 ][ 328 ],
   alphaCSR[ 72 ][ 329 ],
   alphaCSR[ 72 ][ 330 ],
   alphaCSR[ 72 ][ 331 ],
   alphaCSR[ 72 ][ 332 ],
   alphaCSR[ 72 ][ 333 ],
   alphaCSR[ 72 ][ 334 ],
   alphaCSR[ 72 ][ 335 ],
   alphaCSR[ 72 ][ 336 ],
   alphaCSR[ 72 ][ 337 ],
   alphaCSR[ 72 ][ 338 ],
   alphaCSR[ 72 ][ 339 ],
   alphaCSR[ 72 ][ 340 ],
   alphaCSR[ 72 ][ 341 ],
   alphaCSR[ 72 ][ 342 ],
   alphaCSR[ 72 ][ 343 ],
   alphaCSR[ 72 ][ 344 ],
   alphaCSR[ 72 ][ 345 ],
   alphaCSR[ 72 ][ 346 ],
   alphaCSR[ 72 ][ 347 ],
   alphaCSR[ 72 ][ 348 ],
   alphaCSR[ 72 ][ 349 ],
   alphaCSR[ 72 ][ 350 ],
   alphaCSR[ 72 ][ 351 ],
   alphaCSR[ 72 ][ 352 ],
   alphaCSR[ 72 ][ 353 ],
   alphaCSR[ 72 ][ 354 ],
   alphaCSR[ 72 ][ 355 ],
   alphaCSR[ 72 ][ 356 ],
   alphaCSR[ 72 ][ 357 ],
   alphaCSR[ 72 ][ 358 ],
   alphaCSR[ 72 ][ 359 ],
   alphaCSR[ 72 ][ 360 ],
   alphaCSR[ 72 ][ 361 ],
   alphaCSR[ 72 ][ 362 ],
   alphaCSR[ 72 ][ 363 ],
   alphaCSR[ 72 ][ 364 ],
   alphaCSR[ 72 ][ 365 ],
   alphaCSR[ 72 ][ 366 ],
   alphaCSR[ 72 ][ 367 ],
   alphaCSR[ 72 ][ 368 ],
   alphaCSR[ 72 ][ 369 ],
   alphaCSR[ 72 ][ 370 ],
   alphaCSR[ 72 ][ 371 ],
   alphaCSR[ 72 ][ 372 ],
   alphaCSR[ 72 ][ 373 ],
   alphaCSR[ 72 ][ 374 ],
   alphaCSR[ 72 ][ 375 ],
   alphaCSR[ 72 ][ 376 ],
   alphaCSR[ 72 ][ 377 ],
   alphaCSR[ 72 ][ 378 ],
   alphaCSR[ 72 ][ 379 ],
   alphaCSR[ 72 ][ 380 ],
   alphaCSR[ 72 ][ 381 ],
   alphaCSR[ 72 ][ 382 ],
   alphaCSR[ 72 ][ 383 ],
   alphaCSR[ 73 ][ 0 ],
   alphaCSR[ 73 ][ 1 ],
   alphaCSR[ 73 ][ 2 ],
   alphaCSR[ 73 ][ 3 ],
   alphaCSR[ 73 ][ 4 ],
   alphaCSR[ 73 ][ 5 ],
   alphaCSR[ 73 ][ 6 ],
   alphaCSR[ 73 ][ 7 ],
   alphaCSR[ 73 ][ 8 ],
   alphaCSR[ 73 ][ 9 ],
   alphaCSR[ 73 ][ 10 ],
   alphaCSR[ 73 ][ 11 ],
   alphaCSR[ 73 ][ 12 ],
   alphaCSR[ 73 ][ 13 ],
   alphaCSR[ 73 ][ 14 ],
   alphaCSR[ 73 ][ 15 ],
   alphaCSR[ 73 ][ 16 ],
   alphaCSR[ 73 ][ 17 ],
   alphaCSR[ 73 ][ 18 ],
   alphaCSR[ 73 ][ 19 ],
   alphaCSR[ 73 ][ 20 ],
   alphaCSR[ 73 ][ 21 ],
   alphaCSR[ 73 ][ 22 ],
   alphaCSR[ 73 ][ 23 ],
   alphaCSR[ 73 ][ 24 ],
   alphaCSR[ 73 ][ 25 ],
   alphaCSR[ 73 ][ 26 ],
   alphaCSR[ 73 ][ 27 ],
   alphaCSR[ 73 ][ 28 ],
   alphaCSR[ 73 ][ 29 ],
   alphaCSR[ 73 ][ 30 ],
   alphaCSR[ 73 ][ 31 ],
   alphaCSR[ 73 ][ 32 ],
   alphaCSR[ 73 ][ 33 ],
   alphaCSR[ 73 ][ 34 ],
   alphaCSR[ 73 ][ 35 ],
   alphaCSR[ 73 ][ 36 ],
   alphaCSR[ 73 ][ 37 ],
   alphaCSR[ 73 ][ 38 ],
   alphaCSR[ 73 ][ 39 ],
   alphaCSR[ 73 ][ 40 ],
   alphaCSR[ 73 ][ 41 ],
   alphaCSR[ 73 ][ 42 ],
   alphaCSR[ 73 ][ 43 ],
   alphaCSR[ 73 ][ 44 ],
   alphaCSR[ 73 ][ 45 ],
   alphaCSR[ 73 ][ 46 ],
   alphaCSR[ 73 ][ 47 ],
   alphaCSR[ 73 ][ 48 ],
   alphaCSR[ 73 ][ 49 ],
   alphaCSR[ 73 ][ 50 ],
   alphaCSR[ 73 ][ 51 ],
   alphaCSR[ 73 ][ 52 ],
   alphaCSR[ 73 ][ 53 ],
   alphaCSR[ 73 ][ 54 ],
   alphaCSR[ 73 ][ 55 ],
   alphaCSR[ 73 ][ 56 ],
   alphaCSR[ 73 ][ 57 ],
   alphaCSR[ 73 ][ 58 ],
   alphaCSR[ 73 ][ 59 ],
   alphaCSR[ 73 ][ 60 ],
   alphaCSR[ 73 ][ 61 ],
   alphaCSR[ 73 ][ 62 ],
   alphaCSR[ 73 ][ 63 ],
   alphaCSR[ 73 ][ 64 ],
   alphaCSR[ 73 ][ 65 ],
   alphaCSR[ 73 ][ 66 ],
   alphaCSR[ 73 ][ 67 ],
   alphaCSR[ 73 ][ 68 ],
   alphaCSR[ 73 ][ 69 ],
   alphaCSR[ 73 ][ 70 ],
   alphaCSR[ 73 ][ 71 ],
   alphaCSR[ 73 ][ 72 ],
   alphaCSR[ 73 ][ 73 ],
   alphaCSR[ 73 ][ 74 ],
   alphaCSR[ 73 ][ 75 ],
   alphaCSR[ 73 ][ 76 ],
   alphaCSR[ 73 ][ 77 ],
   alphaCSR[ 73 ][ 78 ],
   alphaCSR[ 73 ][ 79 ],
   alphaCSR[ 73 ][ 80 ],
   alphaCSR[ 73 ][ 81 ],
   alphaCSR[ 73 ][ 82 ],
   alphaCSR[ 73 ][ 83 ],
   alphaCSR[ 73 ][ 84 ],
   alphaCSR[ 73 ][ 85 ],
   alphaCSR[ 73 ][ 86 ],
   alphaCSR[ 73 ][ 87 ],
   alphaCSR[ 73 ][ 88 ],
   alphaCSR[ 73 ][ 89 ],
   alphaCSR[ 73 ][ 90 ],
   alphaCSR[ 73 ][ 91 ],
   alphaCSR[ 73 ][ 92 ],
   alphaCSR[ 73 ][ 93 ],
   alphaCSR[ 73 ][ 94 ],
   alphaCSR[ 73 ][ 95 ],
   alphaCSR[ 73 ][ 96 ],
   alphaCSR[ 73 ][ 97 ],
   alphaCSR[ 73 ][ 98 ],
   alphaCSR[ 73 ][ 99 ],
   alphaCSR[ 73 ][ 100 ],
   alphaCSR[ 73 ][ 101 ],
   alphaCSR[ 73 ][ 102 ],
   alphaCSR[ 73 ][ 103 ],
   alphaCSR[ 73 ][ 104 ],
   alphaCSR[ 73 ][ 105 ],
   alphaCSR[ 73 ][ 106 ],
   alphaCSR[ 73 ][ 107 ],
   alphaCSR[ 73 ][ 108 ],
   alphaCSR[ 73 ][ 109 ],
   alphaCSR[ 73 ][ 110 ],
   alphaCSR[ 73 ][ 111 ],
   alphaCSR[ 73 ][ 112 ],
   alphaCSR[ 73 ][ 113 ],
   alphaCSR[ 73 ][ 114 ],
   alphaCSR[ 73 ][ 115 ],
   alphaCSR[ 73 ][ 116 ],
   alphaCSR[ 73 ][ 117 ],
   alphaCSR[ 73 ][ 118 ],
   alphaCSR[ 73 ][ 119 ],
   alphaCSR[ 73 ][ 120 ],
   alphaCSR[ 73 ][ 121 ],
   alphaCSR[ 73 ][ 122 ],
   alphaCSR[ 73 ][ 123 ],
   alphaCSR[ 73 ][ 124 ],
   alphaCSR[ 73 ][ 125 ],
   alphaCSR[ 73 ][ 126 ],
   alphaCSR[ 73 ][ 127 ],
   alphaCSR[ 73 ][ 128 ],
   alphaCSR[ 73 ][ 129 ],
   alphaCSR[ 73 ][ 130 ],
   alphaCSR[ 73 ][ 131 ],
   alphaCSR[ 73 ][ 132 ],
   alphaCSR[ 73 ][ 133 ],
   alphaCSR[ 73 ][ 134 ],
   alphaCSR[ 73 ][ 135 ],
   alphaCSR[ 73 ][ 136 ],
   alphaCSR[ 73 ][ 137 ],
   alphaCSR[ 73 ][ 138 ],
   alphaCSR[ 73 ][ 139 ],
   alphaCSR[ 73 ][ 140 ],
   alphaCSR[ 73 ][ 141 ],
   alphaCSR[ 73 ][ 142 ],
   alphaCSR[ 73 ][ 143 ],
   alphaCSR[ 73 ][ 144 ],
   alphaCSR[ 73 ][ 145 ],
   alphaCSR[ 73 ][ 146 ],
   alphaCSR[ 73 ][ 147 ],
   alphaCSR[ 73 ][ 148 ],
   alphaCSR[ 73 ][ 149 ],
   alphaCSR[ 73 ][ 150 ],
   alphaCSR[ 73 ][ 151 ],
   alphaCSR[ 73 ][ 152 ],
   alphaCSR[ 73 ][ 153 ],
   alphaCSR[ 73 ][ 154 ],
   alphaCSR[ 73 ][ 155 ],
   alphaCSR[ 73 ][ 156 ],
   alphaCSR[ 73 ][ 157 ],
   alphaCSR[ 73 ][ 158 ],
   alphaCSR[ 73 ][ 159 ],
   alphaCSR[ 73 ][ 160 ],
   alphaCSR[ 73 ][ 161 ],
   alphaCSR[ 73 ][ 162 ],
   alphaCSR[ 73 ][ 163 ],
   alphaCSR[ 73 ][ 164 ],
   alphaCSR[ 73 ][ 165 ],
   alphaCSR[ 73 ][ 166 ],
   alphaCSR[ 73 ][ 167 ],
   alphaCSR[ 73 ][ 168 ],
   alphaCSR[ 73 ][ 169 ],
   alphaCSR[ 73 ][ 170 ],
   alphaCSR[ 73 ][ 171 ],
   alphaCSR[ 73 ][ 172 ],
   alphaCSR[ 73 ][ 173 ],
   alphaCSR[ 73 ][ 174 ],
   alphaCSR[ 73 ][ 175 ],
   alphaCSR[ 73 ][ 176 ],
   alphaCSR[ 73 ][ 177 ],
   alphaCSR[ 73 ][ 178 ],
   alphaCSR[ 73 ][ 179 ],
   alphaCSR[ 73 ][ 180 ],
   alphaCSR[ 73 ][ 181 ],
   alphaCSR[ 73 ][ 182 ],
   alphaCSR[ 73 ][ 183 ],
   alphaCSR[ 73 ][ 184 ],
   alphaCSR[ 73 ][ 185 ],
   alphaCSR[ 73 ][ 186 ],
   alphaCSR[ 73 ][ 187 ],
   alphaCSR[ 73 ][ 188 ],
   alphaCSR[ 73 ][ 189 ],
   alphaCSR[ 73 ][ 190 ],
   alphaCSR[ 73 ][ 191 ],
   alphaCSR[ 73 ][ 192 ],
   alphaCSR[ 73 ][ 193 ],
   alphaCSR[ 73 ][ 194 ],
   alphaCSR[ 73 ][ 195 ],
   alphaCSR[ 73 ][ 196 ],
   alphaCSR[ 73 ][ 197 ],
   alphaCSR[ 73 ][ 198 ],
   alphaCSR[ 73 ][ 199 ],
   alphaCSR[ 73 ][ 200 ],
   alphaCSR[ 73 ][ 201 ],
   alphaCSR[ 73 ][ 202 ],
   alphaCSR[ 73 ][ 203 ],
   alphaCSR[ 73 ][ 204 ],
   alphaCSR[ 73 ][ 205 ],
   alphaCSR[ 73 ][ 206 ],
   alphaCSR[ 73 ][ 207 ],
   alphaCSR[ 73 ][ 208 ],
   alphaCSR[ 73 ][ 209 ],
   alphaCSR[ 73 ][ 210 ],
   alphaCSR[ 73 ][ 211 ],
   alphaCSR[ 73 ][ 212 ],
   alphaCSR[ 73 ][ 213 ],
   alphaCSR[ 73 ][ 214 ],
   alphaCSR[ 73 ][ 215 ],
   alphaCSR[ 73 ][ 216 ],
   alphaCSR[ 73 ][ 217 ],
   alphaCSR[ 73 ][ 218 ],
   alphaCSR[ 73 ][ 219 ],
   alphaCSR[ 73 ][ 220 ],
   alphaCSR[ 73 ][ 221 ],
   alphaCSR[ 73 ][ 222 ],
   alphaCSR[ 73 ][ 223 ],
   alphaCSR[ 73 ][ 224 ],
   alphaCSR[ 73 ][ 225 ],
   alphaCSR[ 73 ][ 226 ],
   alphaCSR[ 73 ][ 227 ],
   alphaCSR[ 73 ][ 228 ],
   alphaCSR[ 73 ][ 229 ],
   alphaCSR[ 73 ][ 230 ],
   alphaCSR[ 73 ][ 231 ],
   alphaCSR[ 73 ][ 232 ],
   alphaCSR[ 73 ][ 233 ],
   alphaCSR[ 73 ][ 234 ],
   alphaCSR[ 73 ][ 235 ],
   alphaCSR[ 73 ][ 236 ],
   alphaCSR[ 73 ][ 237 ],
   alphaCSR[ 73 ][ 238 ],
   alphaCSR[ 73 ][ 239 ],
   alphaCSR[ 73 ][ 240 ],
   alphaCSR[ 73 ][ 241 ],
   alphaCSR[ 73 ][ 242 ],
   alphaCSR[ 73 ][ 243 ],
   alphaCSR[ 73 ][ 244 ],
   alphaCSR[ 73 ][ 245 ],
   alphaCSR[ 73 ][ 246 ],
   alphaCSR[ 73 ][ 247 ],
   alphaCSR[ 73 ][ 248 ],
   alphaCSR[ 73 ][ 249 ],
   alphaCSR[ 73 ][ 250 ],
   alphaCSR[ 73 ][ 251 ],
   alphaCSR[ 73 ][ 252 ],
   alphaCSR[ 73 ][ 253 ],
   alphaCSR[ 73 ][ 254 ],
   alphaCSR[ 73 ][ 255 ],
   alphaCSR[ 73 ][ 256 ],
   alphaCSR[ 73 ][ 257 ],
   alphaCSR[ 73 ][ 258 ],
   alphaCSR[ 73 ][ 259 ],
   alphaCSR[ 73 ][ 260 ],
   alphaCSR[ 73 ][ 261 ],
   alphaCSR[ 73 ][ 262 ],
   alphaCSR[ 73 ][ 263 ],
   alphaCSR[ 73 ][ 264 ],
   alphaCSR[ 73 ][ 265 ],
   alphaCSR[ 73 ][ 266 ],
   alphaCSR[ 73 ][ 267 ],
   alphaCSR[ 73 ][ 268 ],
   alphaCSR[ 73 ][ 269 ],
   alphaCSR[ 73 ][ 270 ],
   alphaCSR[ 73 ][ 271 ],
   alphaCSR[ 73 ][ 272 ],
   alphaCSR[ 73 ][ 273 ],
   alphaCSR[ 73 ][ 274 ],
   alphaCSR[ 73 ][ 275 ],
   alphaCSR[ 73 ][ 276 ],
   alphaCSR[ 73 ][ 277 ],
   alphaCSR[ 73 ][ 278 ],
   alphaCSR[ 73 ][ 279 ],
   alphaCSR[ 73 ][ 280 ],
   alphaCSR[ 73 ][ 281 ],
   alphaCSR[ 73 ][ 282 ],
   alphaCSR[ 73 ][ 283 ],
   alphaCSR[ 73 ][ 284 ],
   alphaCSR[ 73 ][ 285 ],
   alphaCSR[ 73 ][ 286 ],
   alphaCSR[ 73 ][ 287 ],
   alphaCSR[ 73 ][ 288 ],
   alphaCSR[ 73 ][ 289 ],
   alphaCSR[ 73 ][ 290 ],
   alphaCSR[ 73 ][ 291 ],
   alphaCSR[ 73 ][ 292 ],
   alphaCSR[ 73 ][ 293 ],
   alphaCSR[ 73 ][ 294 ],
   alphaCSR[ 73 ][ 295 ],
   alphaCSR[ 73 ][ 296 ],
   alphaCSR[ 73 ][ 297 ],
   alphaCSR[ 73 ][ 298 ],
   alphaCSR[ 73 ][ 299 ],
   alphaCSR[ 73 ][ 300 ],
   alphaCSR[ 73 ][ 301 ],
   alphaCSR[ 73 ][ 302 ],
   alphaCSR[ 73 ][ 303 ],
   alphaCSR[ 73 ][ 304 ],
   alphaCSR[ 73 ][ 305 ],
   alphaCSR[ 73 ][ 306 ],
   alphaCSR[ 73 ][ 307 ],
   alphaCSR[ 73 ][ 308 ],
   alphaCSR[ 73 ][ 309 ],
   alphaCSR[ 73 ][ 310 ],
   alphaCSR[ 73 ][ 311 ],
   alphaCSR[ 73 ][ 312 ],
   alphaCSR[ 73 ][ 313 ],
   alphaCSR[ 73 ][ 314 ],
   alphaCSR[ 73 ][ 315 ],
   alphaCSR[ 73 ][ 316 ],
   alphaCSR[ 73 ][ 317 ],
   alphaCSR[ 73 ][ 318 ],
   alphaCSR[ 73 ][ 319 ],
   alphaCSR[ 73 ][ 320 ],
   alphaCSR[ 73 ][ 321 ],
   alphaCSR[ 73 ][ 322 ],
   alphaCSR[ 73 ][ 323 ],
   alphaCSR[ 73 ][ 324 ],
   alphaCSR[ 73 ][ 325 ],
   alphaCSR[ 73 ][ 326 ],
   alphaCSR[ 73 ][ 327 ],
   alphaCSR[ 73 ][ 328 ],
   alphaCSR[ 73 ][ 329 ],
   alphaCSR[ 73 ][ 330 ],
   alphaCSR[ 73 ][ 331 ],
   alphaCSR[ 73 ][ 332 ],
   alphaCSR[ 73 ][ 333 ],
   alphaCSR[ 73 ][ 334 ],
   alphaCSR[ 73 ][ 335 ],
   alphaCSR[ 73 ][ 336 ],
   alphaCSR[ 73 ][ 337 ],
   alphaCSR[ 73 ][ 338 ],
   alphaCSR[ 73 ][ 339 ],
   alphaCSR[ 73 ][ 340 ],
   alphaCSR[ 73 ][ 341 ],
   alphaCSR[ 73 ][ 342 ],
   alphaCSR[ 73 ][ 343 ],
   alphaCSR[ 73 ][ 344 ],
   alphaCSR[ 73 ][ 345 ],
   alphaCSR[ 73 ][ 346 ],
   alphaCSR[ 73 ][ 347 ],
   alphaCSR[ 73 ][ 348 ],
   alphaCSR[ 73 ][ 349 ],
   alphaCSR[ 73 ][ 350 ],
   alphaCSR[ 73 ][ 351 ],
   alphaCSR[ 73 ][ 352 ],
   alphaCSR[ 73 ][ 353 ],
   alphaCSR[ 73 ][ 354 ],
   alphaCSR[ 73 ][ 355 ],
   alphaCSR[ 73 ][ 356 ],
   alphaCSR[ 73 ][ 357 ],
   alphaCSR[ 73 ][ 358 ],
   alphaCSR[ 73 ][ 359 ],
   alphaCSR[ 73 ][ 360 ],
   alphaCSR[ 73 ][ 361 ],
   alphaCSR[ 73 ][ 362 ],
   alphaCSR[ 73 ][ 363 ],
   alphaCSR[ 73 ][ 364 ],
   alphaCSR[ 73 ][ 365 ],
   alphaCSR[ 73 ][ 366 ],
   alphaCSR[ 73 ][ 367 ],
   alphaCSR[ 73 ][ 368 ],
   alphaCSR[ 73 ][ 369 ],
   alphaCSR[ 73 ][ 370 ],
   alphaCSR[ 73 ][ 371 ],
   alphaCSR[ 73 ][ 372 ],
   alphaCSR[ 73 ][ 373 ],
   alphaCSR[ 73 ][ 374 ],
   alphaCSR[ 73 ][ 375 ],
   alphaCSR[ 73 ][ 376 ],
   alphaCSR[ 73 ][ 377 ],
   alphaCSR[ 73 ][ 378 ],
   alphaCSR[ 73 ][ 379 ],
   alphaCSR[ 73 ][ 380 ],
   alphaCSR[ 73 ][ 381 ],
   alphaCSR[ 73 ][ 382 ],
   alphaCSR[ 73 ][ 383 ],
   alphaCSR[ 74 ][ 0 ],
   alphaCSR[ 74 ][ 1 ],
   alphaCSR[ 74 ][ 2 ],
   alphaCSR[ 74 ][ 3 ],
   alphaCSR[ 74 ][ 4 ],
   alphaCSR[ 74 ][ 5 ],
   alphaCSR[ 74 ][ 6 ],
   alphaCSR[ 74 ][ 7 ],
   alphaCSR[ 74 ][ 8 ],
   alphaCSR[ 74 ][ 9 ],
   alphaCSR[ 74 ][ 10 ],
   alphaCSR[ 74 ][ 11 ],
   alphaCSR[ 74 ][ 12 ],
   alphaCSR[ 74 ][ 13 ],
   alphaCSR[ 74 ][ 14 ],
   alphaCSR[ 74 ][ 15 ],
   alphaCSR[ 74 ][ 16 ],
   alphaCSR[ 74 ][ 17 ],
   alphaCSR[ 74 ][ 18 ],
   alphaCSR[ 74 ][ 19 ],
   alphaCSR[ 74 ][ 20 ],
   alphaCSR[ 74 ][ 21 ],
   alphaCSR[ 74 ][ 22 ],
   alphaCSR[ 74 ][ 23 ],
   alphaCSR[ 74 ][ 24 ],
   alphaCSR[ 74 ][ 25 ],
   alphaCSR[ 74 ][ 26 ],
   alphaCSR[ 74 ][ 27 ],
   alphaCSR[ 74 ][ 28 ],
   alphaCSR[ 74 ][ 29 ],
   alphaCSR[ 74 ][ 30 ],
   alphaCSR[ 74 ][ 31 ],
   alphaCSR[ 74 ][ 32 ],
   alphaCSR[ 74 ][ 33 ],
   alphaCSR[ 74 ][ 34 ],
   alphaCSR[ 74 ][ 35 ],
   alphaCSR[ 74 ][ 36 ],
   alphaCSR[ 74 ][ 37 ],
   alphaCSR[ 74 ][ 38 ],
   alphaCSR[ 74 ][ 39 ],
   alphaCSR[ 74 ][ 40 ],
   alphaCSR[ 74 ][ 41 ],
   alphaCSR[ 74 ][ 42 ],
   alphaCSR[ 74 ][ 43 ],
   alphaCSR[ 74 ][ 44 ],
   alphaCSR[ 74 ][ 45 ],
   alphaCSR[ 74 ][ 46 ],
   alphaCSR[ 74 ][ 47 ],
   alphaCSR[ 74 ][ 48 ],
   alphaCSR[ 74 ][ 49 ],
   alphaCSR[ 74 ][ 50 ],
   alphaCSR[ 74 ][ 51 ],
   alphaCSR[ 74 ][ 52 ],
   alphaCSR[ 74 ][ 53 ],
   alphaCSR[ 74 ][ 54 ],
   alphaCSR[ 74 ][ 55 ],
   alphaCSR[ 74 ][ 56 ],
   alphaCSR[ 74 ][ 57 ],
   alphaCSR[ 74 ][ 58 ],
   alphaCSR[ 74 ][ 59 ],
   alphaCSR[ 74 ][ 60 ],
   alphaCSR[ 74 ][ 61 ],
   alphaCSR[ 74 ][ 62 ],
   alphaCSR[ 74 ][ 63 ],
   alphaCSR[ 74 ][ 64 ],
   alphaCSR[ 74 ][ 65 ],
   alphaCSR[ 74 ][ 66 ],
   alphaCSR[ 74 ][ 67 ],
   alphaCSR[ 74 ][ 68 ],
   alphaCSR[ 74 ][ 69 ],
   alphaCSR[ 74 ][ 70 ],
   alphaCSR[ 74 ][ 71 ],
   alphaCSR[ 74 ][ 72 ],
   alphaCSR[ 74 ][ 73 ],
   alphaCSR[ 74 ][ 74 ],
   alphaCSR[ 74 ][ 75 ],
   alphaCSR[ 74 ][ 76 ],
   alphaCSR[ 74 ][ 77 ],
   alphaCSR[ 74 ][ 78 ],
   alphaCSR[ 74 ][ 79 ],
   alphaCSR[ 74 ][ 80 ],
   alphaCSR[ 74 ][ 81 ],
   alphaCSR[ 74 ][ 82 ],
   alphaCSR[ 74 ][ 83 ],
   alphaCSR[ 74 ][ 84 ],
   alphaCSR[ 74 ][ 85 ],
   alphaCSR[ 74 ][ 86 ],
   alphaCSR[ 74 ][ 87 ],
   alphaCSR[ 74 ][ 88 ],
   alphaCSR[ 74 ][ 89 ],
   alphaCSR[ 74 ][ 90 ],
   alphaCSR[ 74 ][ 91 ],
   alphaCSR[ 74 ][ 92 ],
   alphaCSR[ 74 ][ 93 ],
   alphaCSR[ 74 ][ 94 ],
   alphaCSR[ 74 ][ 95 ],
   alphaCSR[ 74 ][ 96 ],
   alphaCSR[ 74 ][ 97 ],
   alphaCSR[ 74 ][ 98 ],
   alphaCSR[ 74 ][ 99 ],
   alphaCSR[ 74 ][ 100 ],
   alphaCSR[ 74 ][ 101 ],
   alphaCSR[ 74 ][ 102 ],
   alphaCSR[ 74 ][ 103 ],
   alphaCSR[ 74 ][ 104 ],
   alphaCSR[ 74 ][ 105 ],
   alphaCSR[ 74 ][ 106 ],
   alphaCSR[ 74 ][ 107 ],
   alphaCSR[ 74 ][ 108 ],
   alphaCSR[ 74 ][ 109 ],
   alphaCSR[ 74 ][ 110 ],
   alphaCSR[ 74 ][ 111 ],
   alphaCSR[ 74 ][ 112 ],
   alphaCSR[ 74 ][ 113 ],
   alphaCSR[ 74 ][ 114 ],
   alphaCSR[ 74 ][ 115 ],
   alphaCSR[ 74 ][ 116 ],
   alphaCSR[ 74 ][ 117 ],
   alphaCSR[ 74 ][ 118 ],
   alphaCSR[ 74 ][ 119 ],
   alphaCSR[ 74 ][ 120 ],
   alphaCSR[ 74 ][ 121 ],
   alphaCSR[ 74 ][ 122 ],
   alphaCSR[ 74 ][ 123 ],
   alphaCSR[ 74 ][ 124 ],
   alphaCSR[ 74 ][ 125 ],
   alphaCSR[ 74 ][ 126 ],
   alphaCSR[ 74 ][ 127 ],
   alphaCSR[ 74 ][ 128 ],
   alphaCSR[ 74 ][ 129 ],
   alphaCSR[ 74 ][ 130 ],
   alphaCSR[ 74 ][ 131 ],
   alphaCSR[ 74 ][ 132 ],
   alphaCSR[ 74 ][ 133 ],
   alphaCSR[ 74 ][ 134 ],
   alphaCSR[ 74 ][ 135 ],
   alphaCSR[ 74 ][ 136 ],
   alphaCSR[ 74 ][ 137 ],
   alphaCSR[ 74 ][ 138 ],
   alphaCSR[ 74 ][ 139 ],
   alphaCSR[ 74 ][ 140 ],
   alphaCSR[ 74 ][ 141 ],
   alphaCSR[ 74 ][ 142 ],
   alphaCSR[ 74 ][ 143 ],
   alphaCSR[ 74 ][ 144 ],
   alphaCSR[ 74 ][ 145 ],
   alphaCSR[ 74 ][ 146 ],
   alphaCSR[ 74 ][ 147 ],
   alphaCSR[ 74 ][ 148 ],
   alphaCSR[ 74 ][ 149 ],
   alphaCSR[ 74 ][ 150 ],
   alphaCSR[ 74 ][ 151 ],
   alphaCSR[ 74 ][ 152 ],
   alphaCSR[ 74 ][ 153 ],
   alphaCSR[ 74 ][ 154 ],
   alphaCSR[ 74 ][ 155 ],
   alphaCSR[ 74 ][ 156 ],
   alphaCSR[ 74 ][ 157 ],
   alphaCSR[ 74 ][ 158 ],
   alphaCSR[ 74 ][ 159 ],
   alphaCSR[ 74 ][ 160 ],
   alphaCSR[ 74 ][ 161 ],
   alphaCSR[ 74 ][ 162 ],
   alphaCSR[ 74 ][ 163 ],
   alphaCSR[ 74 ][ 164 ],
   alphaCSR[ 74 ][ 165 ],
   alphaCSR[ 74 ][ 166 ],
   alphaCSR[ 74 ][ 167 ],
   alphaCSR[ 74 ][ 168 ],
   alphaCSR[ 74 ][ 169 ],
   alphaCSR[ 74 ][ 170 ],
   alphaCSR[ 74 ][ 171 ],
   alphaCSR[ 74 ][ 172 ],
   alphaCSR[ 74 ][ 173 ],
   alphaCSR[ 74 ][ 174 ],
   alphaCSR[ 74 ][ 175 ],
   alphaCSR[ 74 ][ 176 ],
   alphaCSR[ 74 ][ 177 ],
   alphaCSR[ 74 ][ 178 ],
   alphaCSR[ 74 ][ 179 ],
   alphaCSR[ 74 ][ 180 ],
   alphaCSR[ 74 ][ 181 ],
   alphaCSR[ 74 ][ 182 ],
   alphaCSR[ 74 ][ 183 ],
   alphaCSR[ 74 ][ 184 ],
   alphaCSR[ 74 ][ 185 ],
   alphaCSR[ 74 ][ 186 ],
   alphaCSR[ 74 ][ 187 ],
   alphaCSR[ 74 ][ 188 ],
   alphaCSR[ 74 ][ 189 ],
   alphaCSR[ 74 ][ 190 ],
   alphaCSR[ 74 ][ 191 ],
   alphaCSR[ 74 ][ 192 ],
   alphaCSR[ 74 ][ 193 ],
   alphaCSR[ 74 ][ 194 ],
   alphaCSR[ 74 ][ 195 ],
   alphaCSR[ 74 ][ 196 ],
   alphaCSR[ 74 ][ 197 ],
   alphaCSR[ 74 ][ 198 ],
   alphaCSR[ 74 ][ 199 ],
   alphaCSR[ 74 ][ 200 ],
   alphaCSR[ 74 ][ 201 ],
   alphaCSR[ 74 ][ 202 ],
   alphaCSR[ 74 ][ 203 ],
   alphaCSR[ 74 ][ 204 ],
   alphaCSR[ 74 ][ 205 ],
   alphaCSR[ 74 ][ 206 ],
   alphaCSR[ 74 ][ 207 ],
   alphaCSR[ 74 ][ 208 ],
   alphaCSR[ 74 ][ 209 ],
   alphaCSR[ 74 ][ 210 ],
   alphaCSR[ 74 ][ 211 ],
   alphaCSR[ 74 ][ 212 ],
   alphaCSR[ 74 ][ 213 ],
   alphaCSR[ 74 ][ 214 ],
   alphaCSR[ 74 ][ 215 ],
   alphaCSR[ 74 ][ 216 ],
   alphaCSR[ 74 ][ 217 ],
   alphaCSR[ 74 ][ 218 ],
   alphaCSR[ 74 ][ 219 ],
   alphaCSR[ 74 ][ 220 ],
   alphaCSR[ 74 ][ 221 ],
   alphaCSR[ 74 ][ 222 ],
   alphaCSR[ 74 ][ 223 ],
   alphaCSR[ 74 ][ 224 ],
   alphaCSR[ 74 ][ 225 ],
   alphaCSR[ 74 ][ 226 ],
   alphaCSR[ 74 ][ 227 ],
   alphaCSR[ 74 ][ 228 ],
   alphaCSR[ 74 ][ 229 ],
   alphaCSR[ 74 ][ 230 ],
   alphaCSR[ 74 ][ 231 ],
   alphaCSR[ 74 ][ 232 ],
   alphaCSR[ 74 ][ 233 ],
   alphaCSR[ 74 ][ 234 ],
   alphaCSR[ 74 ][ 235 ],
   alphaCSR[ 74 ][ 236 ],
   alphaCSR[ 74 ][ 237 ],
   alphaCSR[ 74 ][ 238 ],
   alphaCSR[ 74 ][ 239 ],
   alphaCSR[ 74 ][ 240 ],
   alphaCSR[ 74 ][ 241 ],
   alphaCSR[ 74 ][ 242 ],
   alphaCSR[ 74 ][ 243 ],
   alphaCSR[ 74 ][ 244 ],
   alphaCSR[ 74 ][ 245 ],
   alphaCSR[ 74 ][ 246 ],
   alphaCSR[ 74 ][ 247 ],
   alphaCSR[ 74 ][ 248 ],
   alphaCSR[ 74 ][ 249 ],
   alphaCSR[ 74 ][ 250 ],
   alphaCSR[ 74 ][ 251 ],
   alphaCSR[ 74 ][ 252 ],
   alphaCSR[ 74 ][ 253 ],
   alphaCSR[ 74 ][ 254 ],
   alphaCSR[ 74 ][ 255 ],
   alphaCSR[ 74 ][ 256 ],
   alphaCSR[ 74 ][ 257 ],
   alphaCSR[ 74 ][ 258 ],
   alphaCSR[ 74 ][ 259 ],
   alphaCSR[ 74 ][ 260 ],
   alphaCSR[ 74 ][ 261 ],
   alphaCSR[ 74 ][ 262 ],
   alphaCSR[ 74 ][ 263 ],
   alphaCSR[ 74 ][ 264 ],
   alphaCSR[ 74 ][ 265 ],
   alphaCSR[ 74 ][ 266 ],
   alphaCSR[ 74 ][ 267 ],
   alphaCSR[ 74 ][ 268 ],
   alphaCSR[ 74 ][ 269 ],
   alphaCSR[ 74 ][ 270 ],
   alphaCSR[ 74 ][ 271 ],
   alphaCSR[ 74 ][ 272 ],
   alphaCSR[ 74 ][ 273 ],
   alphaCSR[ 74 ][ 274 ],
   alphaCSR[ 74 ][ 275 ],
   alphaCSR[ 74 ][ 276 ],
   alphaCSR[ 74 ][ 277 ],
   alphaCSR[ 74 ][ 278 ],
   alphaCSR[ 74 ][ 279 ],
   alphaCSR[ 74 ][ 280 ],
   alphaCSR[ 74 ][ 281 ],
   alphaCSR[ 74 ][ 282 ],
   alphaCSR[ 74 ][ 283 ],
   alphaCSR[ 74 ][ 284 ],
   alphaCSR[ 74 ][ 285 ],
   alphaCSR[ 74 ][ 286 ],
   alphaCSR[ 74 ][ 287 ],
   alphaCSR[ 74 ][ 288 ],
   alphaCSR[ 74 ][ 289 ],
   alphaCSR[ 74 ][ 290 ],
   alphaCSR[ 74 ][ 291 ],
   alphaCSR[ 74 ][ 292 ],
   alphaCSR[ 74 ][ 293 ],
   alphaCSR[ 74 ][ 294 ],
   alphaCSR[ 74 ][ 295 ],
   alphaCSR[ 74 ][ 296 ],
   alphaCSR[ 74 ][ 297 ],
   alphaCSR[ 74 ][ 298 ],
   alphaCSR[ 74 ][ 299 ],
   alphaCSR[ 74 ][ 300 ],
   alphaCSR[ 74 ][ 301 ],
   alphaCSR[ 74 ][ 302 ],
   alphaCSR[ 74 ][ 303 ],
   alphaCSR[ 74 ][ 304 ],
   alphaCSR[ 74 ][ 305 ],
   alphaCSR[ 74 ][ 306 ],
   alphaCSR[ 74 ][ 307 ],
   alphaCSR[ 74 ][ 308 ],
   alphaCSR[ 74 ][ 309 ],
   alphaCSR[ 74 ][ 310 ],
   alphaCSR[ 74 ][ 311 ],
   alphaCSR[ 74 ][ 312 ],
   alphaCSR[ 74 ][ 313 ],
   alphaCSR[ 74 ][ 314 ],
   alphaCSR[ 74 ][ 315 ],
   alphaCSR[ 74 ][ 316 ],
   alphaCSR[ 74 ][ 317 ],
   alphaCSR[ 74 ][ 318 ],
   alphaCSR[ 74 ][ 319 ],
   alphaCSR[ 74 ][ 320 ],
   alphaCSR[ 74 ][ 321 ],
   alphaCSR[ 74 ][ 322 ],
   alphaCSR[ 74 ][ 323 ],
   alphaCSR[ 74 ][ 324 ],
   alphaCSR[ 74 ][ 325 ],
   alphaCSR[ 74 ][ 326 ],
   alphaCSR[ 74 ][ 327 ],
   alphaCSR[ 74 ][ 328 ],
   alphaCSR[ 74 ][ 329 ],
   alphaCSR[ 74 ][ 330 ],
   alphaCSR[ 74 ][ 331 ],
   alphaCSR[ 74 ][ 332 ],
   alphaCSR[ 74 ][ 333 ],
   alphaCSR[ 74 ][ 334 ],
   alphaCSR[ 74 ][ 335 ],
   alphaCSR[ 74 ][ 336 ],
   alphaCSR[ 74 ][ 337 ],
   alphaCSR[ 74 ][ 338 ],
   alphaCSR[ 74 ][ 339 ],
   alphaCSR[ 74 ][ 340 ],
   alphaCSR[ 74 ][ 341 ],
   alphaCSR[ 74 ][ 342 ],
   alphaCSR[ 74 ][ 343 ],
   alphaCSR[ 74 ][ 344 ],
   alphaCSR[ 74 ][ 345 ],
   alphaCSR[ 74 ][ 346 ],
   alphaCSR[ 74 ][ 347 ],
   alphaCSR[ 74 ][ 348 ],
   alphaCSR[ 74 ][ 349 ],
   alphaCSR[ 74 ][ 350 ],
   alphaCSR[ 74 ][ 351 ],
   alphaCSR[ 74 ][ 352 ],
   alphaCSR[ 74 ][ 353 ],
   alphaCSR[ 74 ][ 354 ],
   alphaCSR[ 74 ][ 355 ],
   alphaCSR[ 74 ][ 356 ],
   alphaCSR[ 74 ][ 357 ],
   alphaCSR[ 74 ][ 358 ],
   alphaCSR[ 74 ][ 359 ],
   alphaCSR[ 74 ][ 360 ],
   alphaCSR[ 74 ][ 361 ],
   alphaCSR[ 74 ][ 362 ],
   alphaCSR[ 74 ][ 363 ],
   alphaCSR[ 74 ][ 364 ],
   alphaCSR[ 74 ][ 365 ],
   alphaCSR[ 74 ][ 366 ],
   alphaCSR[ 74 ][ 367 ],
   alphaCSR[ 74 ][ 368 ],
   alphaCSR[ 74 ][ 369 ],
   alphaCSR[ 74 ][ 370 ],
   alphaCSR[ 74 ][ 371 ],
   alphaCSR[ 74 ][ 372 ],
   alphaCSR[ 74 ][ 373 ],
   alphaCSR[ 74 ][ 374 ],
   alphaCSR[ 74 ][ 375 ],
   alphaCSR[ 74 ][ 376 ],
   alphaCSR[ 74 ][ 377 ],
   alphaCSR[ 74 ][ 378 ],
   alphaCSR[ 74 ][ 379 ],
   alphaCSR[ 74 ][ 380 ],
   alphaCSR[ 74 ][ 381 ],
   alphaCSR[ 74 ][ 382 ],
   alphaCSR[ 74 ][ 383 ],
   alphaCSR[ 75 ][ 0 ],
   alphaCSR[ 75 ][ 1 ],
   alphaCSR[ 75 ][ 2 ],
   alphaCSR[ 75 ][ 3 ],
   alphaCSR[ 75 ][ 4 ],
   alphaCSR[ 75 ][ 5 ],
   alphaCSR[ 75 ][ 6 ],
   alphaCSR[ 75 ][ 7 ],
   alphaCSR[ 75 ][ 8 ],
   alphaCSR[ 75 ][ 9 ],
   alphaCSR[ 75 ][ 10 ],
   alphaCSR[ 75 ][ 11 ],
   alphaCSR[ 75 ][ 12 ],
   alphaCSR[ 75 ][ 13 ],
   alphaCSR[ 75 ][ 14 ],
   alphaCSR[ 75 ][ 15 ],
   alphaCSR[ 75 ][ 16 ],
   alphaCSR[ 75 ][ 17 ],
   alphaCSR[ 75 ][ 18 ],
   alphaCSR[ 75 ][ 19 ],
   alphaCSR[ 75 ][ 20 ],
   alphaCSR[ 75 ][ 21 ],
   alphaCSR[ 75 ][ 22 ],
   alphaCSR[ 75 ][ 23 ],
   alphaCSR[ 75 ][ 24 ],
   alphaCSR[ 75 ][ 25 ],
   alphaCSR[ 75 ][ 26 ],
   alphaCSR[ 75 ][ 27 ],
   alphaCSR[ 75 ][ 28 ],
   alphaCSR[ 75 ][ 29 ],
   alphaCSR[ 75 ][ 30 ],
   alphaCSR[ 75 ][ 31 ],
   alphaCSR[ 75 ][ 32 ],
   alphaCSR[ 75 ][ 33 ],
   alphaCSR[ 75 ][ 34 ],
   alphaCSR[ 75 ][ 35 ],
   alphaCSR[ 75 ][ 36 ],
   alphaCSR[ 75 ][ 37 ],
   alphaCSR[ 75 ][ 38 ],
   alphaCSR[ 75 ][ 39 ],
   alphaCSR[ 75 ][ 40 ],
   alphaCSR[ 75 ][ 41 ],
   alphaCSR[ 75 ][ 42 ],
   alphaCSR[ 75 ][ 43 ],
   alphaCSR[ 75 ][ 44 ],
   alphaCSR[ 75 ][ 45 ],
   alphaCSR[ 75 ][ 46 ],
   alphaCSR[ 75 ][ 47 ],
   alphaCSR[ 75 ][ 48 ],
   alphaCSR[ 75 ][ 49 ],
   alphaCSR[ 75 ][ 50 ],
   alphaCSR[ 75 ][ 51 ],
   alphaCSR[ 75 ][ 52 ],
   alphaCSR[ 75 ][ 53 ],
   alphaCSR[ 75 ][ 54 ],
   alphaCSR[ 75 ][ 55 ],
   alphaCSR[ 75 ][ 56 ],
   alphaCSR[ 75 ][ 57 ],
   alphaCSR[ 75 ][ 58 ],
   alphaCSR[ 75 ][ 59 ],
   alphaCSR[ 75 ][ 60 ],
   alphaCSR[ 75 ][ 61 ],
   alphaCSR[ 75 ][ 62 ],
   alphaCSR[ 75 ][ 63 ],
   alphaCSR[ 75 ][ 64 ],
   alphaCSR[ 75 ][ 65 ],
   alphaCSR[ 75 ][ 66 ],
   alphaCSR[ 75 ][ 67 ],
   alphaCSR[ 75 ][ 68 ],
   alphaCSR[ 75 ][ 69 ],
   alphaCSR[ 75 ][ 70 ],
   alphaCSR[ 75 ][ 71 ],
   alphaCSR[ 75 ][ 72 ],
   alphaCSR[ 75 ][ 73 ],
   alphaCSR[ 75 ][ 74 ],
   alphaCSR[ 75 ][ 75 ],
   alphaCSR[ 75 ][ 76 ],
   alphaCSR[ 75 ][ 77 ],
   alphaCSR[ 75 ][ 78 ],
   alphaCSR[ 75 ][ 79 ],
   alphaCSR[ 75 ][ 80 ],
   alphaCSR[ 75 ][ 81 ],
   alphaCSR[ 75 ][ 82 ],
   alphaCSR[ 75 ][ 83 ],
   alphaCSR[ 75 ][ 84 ],
   alphaCSR[ 75 ][ 85 ],
   alphaCSR[ 75 ][ 86 ],
   alphaCSR[ 75 ][ 87 ],
   alphaCSR[ 75 ][ 88 ],
   alphaCSR[ 75 ][ 89 ],
   alphaCSR[ 75 ][ 90 ],
   alphaCSR[ 75 ][ 91 ],
   alphaCSR[ 75 ][ 92 ],
   alphaCSR[ 75 ][ 93 ],
   alphaCSR[ 75 ][ 94 ],
   alphaCSR[ 75 ][ 95 ],
   alphaCSR[ 75 ][ 96 ],
   alphaCSR[ 75 ][ 97 ],
   alphaCSR[ 75 ][ 98 ],
   alphaCSR[ 75 ][ 99 ],
   alphaCSR[ 75 ][ 100 ],
   alphaCSR[ 75 ][ 101 ],
   alphaCSR[ 75 ][ 102 ],
   alphaCSR[ 75 ][ 103 ],
   alphaCSR[ 75 ][ 104 ],
   alphaCSR[ 75 ][ 105 ],
   alphaCSR[ 75 ][ 106 ],
   alphaCSR[ 75 ][ 107 ],
   alphaCSR[ 75 ][ 108 ],
   alphaCSR[ 75 ][ 109 ],
   alphaCSR[ 75 ][ 110 ],
   alphaCSR[ 75 ][ 111 ],
   alphaCSR[ 75 ][ 112 ],
   alphaCSR[ 75 ][ 113 ],
   alphaCSR[ 75 ][ 114 ],
   alphaCSR[ 75 ][ 115 ],
   alphaCSR[ 75 ][ 116 ],
   alphaCSR[ 75 ][ 117 ],
   alphaCSR[ 75 ][ 118 ],
   alphaCSR[ 75 ][ 119 ],
   alphaCSR[ 75 ][ 120 ],
   alphaCSR[ 75 ][ 121 ],
   alphaCSR[ 75 ][ 122 ],
   alphaCSR[ 75 ][ 123 ],
   alphaCSR[ 75 ][ 124 ],
   alphaCSR[ 75 ][ 125 ],
   alphaCSR[ 75 ][ 126 ],
   alphaCSR[ 75 ][ 127 ],
   alphaCSR[ 75 ][ 128 ],
   alphaCSR[ 75 ][ 129 ],
   alphaCSR[ 75 ][ 130 ],
   alphaCSR[ 75 ][ 131 ],
   alphaCSR[ 75 ][ 132 ],
   alphaCSR[ 75 ][ 133 ],
   alphaCSR[ 75 ][ 134 ],
   alphaCSR[ 75 ][ 135 ],
   alphaCSR[ 75 ][ 136 ],
   alphaCSR[ 75 ][ 137 ],
   alphaCSR[ 75 ][ 138 ],
   alphaCSR[ 75 ][ 139 ],
   alphaCSR[ 75 ][ 140 ],
   alphaCSR[ 75 ][ 141 ],
   alphaCSR[ 75 ][ 142 ],
   alphaCSR[ 75 ][ 143 ],
   alphaCSR[ 75 ][ 144 ],
   alphaCSR[ 75 ][ 145 ],
   alphaCSR[ 75 ][ 146 ],
   alphaCSR[ 75 ][ 147 ],
   alphaCSR[ 75 ][ 148 ],
   alphaCSR[ 75 ][ 149 ],
   alphaCSR[ 75 ][ 150 ],
   alphaCSR[ 75 ][ 151 ],
   alphaCSR[ 75 ][ 152 ],
   alphaCSR[ 75 ][ 153 ],
   alphaCSR[ 75 ][ 154 ],
   alphaCSR[ 75 ][ 155 ],
   alphaCSR[ 75 ][ 156 ],
   alphaCSR[ 75 ][ 157 ],
   alphaCSR[ 75 ][ 158 ],
   alphaCSR[ 75 ][ 159 ],
   alphaCSR[ 75 ][ 160 ],
   alphaCSR[ 75 ][ 161 ],
   alphaCSR[ 75 ][ 162 ],
   alphaCSR[ 75 ][ 163 ],
   alphaCSR[ 75 ][ 164 ],
   alphaCSR[ 75 ][ 165 ],
   alphaCSR[ 75 ][ 166 ],
   alphaCSR[ 75 ][ 167 ],
   alphaCSR[ 75 ][ 168 ],
   alphaCSR[ 75 ][ 169 ],
   alphaCSR[ 75 ][ 170 ],
   alphaCSR[ 75 ][ 171 ],
   alphaCSR[ 75 ][ 172 ],
   alphaCSR[ 75 ][ 173 ],
   alphaCSR[ 75 ][ 174 ],
   alphaCSR[ 75 ][ 175 ],
   alphaCSR[ 75 ][ 176 ],
   alphaCSR[ 75 ][ 177 ],
   alphaCSR[ 75 ][ 178 ],
   alphaCSR[ 75 ][ 179 ],
   alphaCSR[ 75 ][ 180 ],
   alphaCSR[ 75 ][ 181 ],
   alphaCSR[ 75 ][ 182 ],
   alphaCSR[ 75 ][ 183 ],
   alphaCSR[ 75 ][ 184 ],
   alphaCSR[ 75 ][ 185 ],
   alphaCSR[ 75 ][ 186 ],
   alphaCSR[ 75 ][ 187 ],
   alphaCSR[ 75 ][ 188 ],
   alphaCSR[ 75 ][ 189 ],
   alphaCSR[ 75 ][ 190 ],
   alphaCSR[ 75 ][ 191 ],
   alphaCSR[ 75 ][ 192 ],
   alphaCSR[ 75 ][ 193 ],
   alphaCSR[ 75 ][ 194 ],
   alphaCSR[ 75 ][ 195 ],
   alphaCSR[ 75 ][ 196 ],
   alphaCSR[ 75 ][ 197 ],
   alphaCSR[ 75 ][ 198 ],
   alphaCSR[ 75 ][ 199 ],
   alphaCSR[ 75 ][ 200 ],
   alphaCSR[ 75 ][ 201 ],
   alphaCSR[ 75 ][ 202 ],
   alphaCSR[ 75 ][ 203 ],
   alphaCSR[ 75 ][ 204 ],
   alphaCSR[ 75 ][ 205 ],
   alphaCSR[ 75 ][ 206 ],
   alphaCSR[ 75 ][ 207 ],
   alphaCSR[ 75 ][ 208 ],
   alphaCSR[ 75 ][ 209 ],
   alphaCSR[ 75 ][ 210 ],
   alphaCSR[ 75 ][ 211 ],
   alphaCSR[ 75 ][ 212 ],
   alphaCSR[ 75 ][ 213 ],
   alphaCSR[ 75 ][ 214 ],
   alphaCSR[ 75 ][ 215 ],
   alphaCSR[ 75 ][ 216 ],
   alphaCSR[ 75 ][ 217 ],
   alphaCSR[ 75 ][ 218 ],
   alphaCSR[ 75 ][ 219 ],
   alphaCSR[ 75 ][ 220 ],
   alphaCSR[ 75 ][ 221 ],
   alphaCSR[ 75 ][ 222 ],
   alphaCSR[ 75 ][ 223 ],
   alphaCSR[ 75 ][ 224 ],
   alphaCSR[ 75 ][ 225 ],
   alphaCSR[ 75 ][ 226 ],
   alphaCSR[ 75 ][ 227 ],
   alphaCSR[ 75 ][ 228 ],
   alphaCSR[ 75 ][ 229 ],
   alphaCSR[ 75 ][ 230 ],
   alphaCSR[ 75 ][ 231 ],
   alphaCSR[ 75 ][ 232 ],
   alphaCSR[ 75 ][ 233 ],
   alphaCSR[ 75 ][ 234 ],
   alphaCSR[ 75 ][ 235 ],
   alphaCSR[ 75 ][ 236 ],
   alphaCSR[ 75 ][ 237 ],
   alphaCSR[ 75 ][ 238 ],
   alphaCSR[ 75 ][ 239 ],
   alphaCSR[ 75 ][ 240 ],
   alphaCSR[ 75 ][ 241 ],
   alphaCSR[ 75 ][ 242 ],
   alphaCSR[ 75 ][ 243 ],
   alphaCSR[ 75 ][ 244 ],
   alphaCSR[ 75 ][ 245 ],
   alphaCSR[ 75 ][ 246 ],
   alphaCSR[ 75 ][ 247 ],
   alphaCSR[ 75 ][ 248 ],
   alphaCSR[ 75 ][ 249 ],
   alphaCSR[ 75 ][ 250 ],
   alphaCSR[ 75 ][ 251 ],
   alphaCSR[ 75 ][ 252 ],
   alphaCSR[ 75 ][ 253 ],
   alphaCSR[ 75 ][ 254 ],
   alphaCSR[ 75 ][ 255 ],
   alphaCSR[ 75 ][ 256 ],
   alphaCSR[ 75 ][ 257 ],
   alphaCSR[ 75 ][ 258 ],
   alphaCSR[ 75 ][ 259 ],
   alphaCSR[ 75 ][ 260 ],
   alphaCSR[ 75 ][ 261 ],
   alphaCSR[ 75 ][ 262 ],
   alphaCSR[ 75 ][ 263 ],
   alphaCSR[ 75 ][ 264 ],
   alphaCSR[ 75 ][ 265 ],
   alphaCSR[ 75 ][ 266 ],
   alphaCSR[ 75 ][ 267 ],
   alphaCSR[ 75 ][ 268 ],
   alphaCSR[ 75 ][ 269 ],
   alphaCSR[ 75 ][ 270 ],
   alphaCSR[ 75 ][ 271 ],
   alphaCSR[ 75 ][ 272 ],
   alphaCSR[ 75 ][ 273 ],
   alphaCSR[ 75 ][ 274 ],
   alphaCSR[ 75 ][ 275 ],
   alphaCSR[ 75 ][ 276 ],
   alphaCSR[ 75 ][ 277 ],
   alphaCSR[ 75 ][ 278 ],
   alphaCSR[ 75 ][ 279 ],
   alphaCSR[ 75 ][ 280 ],
   alphaCSR[ 75 ][ 281 ],
   alphaCSR[ 75 ][ 282 ],
   alphaCSR[ 75 ][ 283 ],
   alphaCSR[ 75 ][ 284 ],
   alphaCSR[ 75 ][ 285 ],
   alphaCSR[ 75 ][ 286 ],
   alphaCSR[ 75 ][ 287 ],
   alphaCSR[ 75 ][ 288 ],
   alphaCSR[ 75 ][ 289 ],
   alphaCSR[ 75 ][ 290 ],
   alphaCSR[ 75 ][ 291 ],
   alphaCSR[ 75 ][ 292 ],
   alphaCSR[ 75 ][ 293 ],
   alphaCSR[ 75 ][ 294 ],
   alphaCSR[ 75 ][ 295 ],
   alphaCSR[ 75 ][ 296 ],
   alphaCSR[ 75 ][ 297 ],
   alphaCSR[ 75 ][ 298 ],
   alphaCSR[ 75 ][ 299 ],
   alphaCSR[ 75 ][ 300 ],
   alphaCSR[ 75 ][ 301 ],
   alphaCSR[ 75 ][ 302 ],
   alphaCSR[ 75 ][ 303 ],
   alphaCSR[ 75 ][ 304 ],
   alphaCSR[ 75 ][ 305 ],
   alphaCSR[ 75 ][ 306 ],
   alphaCSR[ 75 ][ 307 ],
   alphaCSR[ 75 ][ 308 ],
   alphaCSR[ 75 ][ 309 ],
   alphaCSR[ 75 ][ 310 ],
   alphaCSR[ 75 ][ 311 ],
   alphaCSR[ 75 ][ 312 ],
   alphaCSR[ 75 ][ 313 ],
   alphaCSR[ 75 ][ 314 ],
   alphaCSR[ 75 ][ 315 ],
   alphaCSR[ 75 ][ 316 ],
   alphaCSR[ 75 ][ 317 ],
   alphaCSR[ 75 ][ 318 ],
   alphaCSR[ 75 ][ 319 ],
   alphaCSR[ 75 ][ 320 ],
   alphaCSR[ 75 ][ 321 ],
   alphaCSR[ 75 ][ 322 ],
   alphaCSR[ 75 ][ 323 ],
   alphaCSR[ 75 ][ 324 ],
   alphaCSR[ 75 ][ 325 ],
   alphaCSR[ 75 ][ 326 ],
   alphaCSR[ 75 ][ 327 ],
   alphaCSR[ 75 ][ 328 ],
   alphaCSR[ 75 ][ 329 ],
   alphaCSR[ 75 ][ 330 ],
   alphaCSR[ 75 ][ 331 ],
   alphaCSR[ 75 ][ 332 ],
   alphaCSR[ 75 ][ 333 ],
   alphaCSR[ 75 ][ 334 ],
   alphaCSR[ 75 ][ 335 ],
   alphaCSR[ 75 ][ 336 ],
   alphaCSR[ 75 ][ 337 ],
   alphaCSR[ 75 ][ 338 ],
   alphaCSR[ 75 ][ 339 ],
   alphaCSR[ 75 ][ 340 ],
   alphaCSR[ 75 ][ 341 ],
   alphaCSR[ 75 ][ 342 ],
   alphaCSR[ 75 ][ 343 ],
   alphaCSR[ 75 ][ 344 ],
   alphaCSR[ 75 ][ 345 ],
   alphaCSR[ 75 ][ 346 ],
   alphaCSR[ 75 ][ 347 ],
   alphaCSR[ 75 ][ 348 ],
   alphaCSR[ 75 ][ 349 ],
   alphaCSR[ 75 ][ 350 ],
   alphaCSR[ 75 ][ 351 ],
   alphaCSR[ 75 ][ 352 ],
   alphaCSR[ 75 ][ 353 ],
   alphaCSR[ 75 ][ 354 ],
   alphaCSR[ 75 ][ 355 ],
   alphaCSR[ 75 ][ 356 ],
   alphaCSR[ 75 ][ 357 ],
   alphaCSR[ 75 ][ 358 ],
   alphaCSR[ 75 ][ 359 ],
   alphaCSR[ 75 ][ 360 ],
   alphaCSR[ 75 ][ 361 ],
   alphaCSR[ 75 ][ 362 ],
   alphaCSR[ 75 ][ 363 ],
   alphaCSR[ 75 ][ 364 ],
   alphaCSR[ 75 ][ 365 ],
   alphaCSR[ 75 ][ 366 ],
   alphaCSR[ 75 ][ 367 ],
   alphaCSR[ 75 ][ 368 ],
   alphaCSR[ 75 ][ 369 ],
   alphaCSR[ 75 ][ 370 ],
   alphaCSR[ 75 ][ 371 ],
   alphaCSR[ 75 ][ 372 ],
   alphaCSR[ 75 ][ 373 ],
   alphaCSR[ 75 ][ 374 ],
   alphaCSR[ 75 ][ 375 ],
   alphaCSR[ 75 ][ 376 ],
   alphaCSR[ 75 ][ 377 ],
   alphaCSR[ 75 ][ 378 ],
   alphaCSR[ 75 ][ 379 ],
   alphaCSR[ 75 ][ 380 ],
   alphaCSR[ 75 ][ 381 ],
   alphaCSR[ 75 ][ 382 ],
   alphaCSR[ 75 ][ 383 ],
   alphaCSR[ 76 ][ 0 ],
   alphaCSR[ 76 ][ 1 ],
   alphaCSR[ 76 ][ 2 ],
   alphaCSR[ 76 ][ 3 ],
   alphaCSR[ 76 ][ 4 ],
   alphaCSR[ 76 ][ 5 ],
   alphaCSR[ 76 ][ 6 ],
   alphaCSR[ 76 ][ 7 ],
   alphaCSR[ 76 ][ 8 ],
   alphaCSR[ 76 ][ 9 ],
   alphaCSR[ 76 ][ 10 ],
   alphaCSR[ 76 ][ 11 ],
   alphaCSR[ 76 ][ 12 ],
   alphaCSR[ 76 ][ 13 ],
   alphaCSR[ 76 ][ 14 ],
   alphaCSR[ 76 ][ 15 ],
   alphaCSR[ 76 ][ 16 ],
   alphaCSR[ 76 ][ 17 ],
   alphaCSR[ 76 ][ 18 ],
   alphaCSR[ 76 ][ 19 ],
   alphaCSR[ 76 ][ 20 ],
   alphaCSR[ 76 ][ 21 ],
   alphaCSR[ 76 ][ 22 ],
   alphaCSR[ 76 ][ 23 ],
   alphaCSR[ 76 ][ 24 ],
   alphaCSR[ 76 ][ 25 ],
   alphaCSR[ 76 ][ 26 ],
   alphaCSR[ 76 ][ 27 ],
   alphaCSR[ 76 ][ 28 ],
   alphaCSR[ 76 ][ 29 ],
   alphaCSR[ 76 ][ 30 ],
   alphaCSR[ 76 ][ 31 ],
   alphaCSR[ 76 ][ 32 ],
   alphaCSR[ 76 ][ 33 ],
   alphaCSR[ 76 ][ 34 ],
   alphaCSR[ 76 ][ 35 ],
   alphaCSR[ 76 ][ 36 ],
   alphaCSR[ 76 ][ 37 ],
   alphaCSR[ 76 ][ 38 ],
   alphaCSR[ 76 ][ 39 ],
   alphaCSR[ 76 ][ 40 ],
   alphaCSR[ 76 ][ 41 ],
   alphaCSR[ 76 ][ 42 ],
   alphaCSR[ 76 ][ 43 ],
   alphaCSR[ 76 ][ 44 ],
   alphaCSR[ 76 ][ 45 ],
   alphaCSR[ 76 ][ 46 ],
   alphaCSR[ 76 ][ 47 ],
   alphaCSR[ 76 ][ 48 ],
   alphaCSR[ 76 ][ 49 ],
   alphaCSR[ 76 ][ 50 ],
   alphaCSR[ 76 ][ 51 ],
   alphaCSR[ 76 ][ 52 ],
   alphaCSR[ 76 ][ 53 ],
   alphaCSR[ 76 ][ 54 ],
   alphaCSR[ 76 ][ 55 ],
   alphaCSR[ 76 ][ 56 ],
   alphaCSR[ 76 ][ 57 ],
   alphaCSR[ 76 ][ 58 ],
   alphaCSR[ 76 ][ 59 ],
   alphaCSR[ 76 ][ 60 ],
   alphaCSR[ 76 ][ 61 ],
   alphaCSR[ 76 ][ 62 ],
   alphaCSR[ 76 ][ 63 ],
   alphaCSR[ 76 ][ 64 ],
   alphaCSR[ 76 ][ 65 ],
   alphaCSR[ 76 ][ 66 ],
   alphaCSR[ 76 ][ 67 ],
   alphaCSR[ 76 ][ 68 ],
   alphaCSR[ 76 ][ 69 ],
   alphaCSR[ 76 ][ 70 ],
   alphaCSR[ 76 ][ 71 ],
   alphaCSR[ 76 ][ 72 ],
   alphaCSR[ 76 ][ 73 ],
   alphaCSR[ 76 ][ 74 ],
   alphaCSR[ 76 ][ 75 ],
   alphaCSR[ 76 ][ 76 ],
   alphaCSR[ 76 ][ 77 ],
   alphaCSR[ 76 ][ 78 ],
   alphaCSR[ 76 ][ 79 ],
   alphaCSR[ 76 ][ 80 ],
   alphaCSR[ 76 ][ 81 ],
   alphaCSR[ 76 ][ 82 ],
   alphaCSR[ 76 ][ 83 ],
   alphaCSR[ 76 ][ 84 ],
   alphaCSR[ 76 ][ 85 ],
   alphaCSR[ 76 ][ 86 ],
   alphaCSR[ 76 ][ 87 ],
   alphaCSR[ 76 ][ 88 ],
   alphaCSR[ 76 ][ 89 ],
   alphaCSR[ 76 ][ 90 ],
   alphaCSR[ 76 ][ 91 ],
   alphaCSR[ 76 ][ 92 ],
   alphaCSR[ 76 ][ 93 ],
   alphaCSR[ 76 ][ 94 ],
   alphaCSR[ 76 ][ 95 ],
   alphaCSR[ 76 ][ 96 ],
   alphaCSR[ 76 ][ 97 ],
   alphaCSR[ 76 ][ 98 ],
   alphaCSR[ 76 ][ 99 ],
   alphaCSR[ 76 ][ 100 ],
   alphaCSR[ 76 ][ 101 ],
   alphaCSR[ 76 ][ 102 ],
   alphaCSR[ 76 ][ 103 ],
   alphaCSR[ 76 ][ 104 ],
   alphaCSR[ 76 ][ 105 ],
   alphaCSR[ 76 ][ 106 ],
   alphaCSR[ 76 ][ 107 ],
   alphaCSR[ 76 ][ 108 ],
   alphaCSR[ 76 ][ 109 ],
   alphaCSR[ 76 ][ 110 ],
   alphaCSR[ 76 ][ 111 ],
   alphaCSR[ 76 ][ 112 ],
   alphaCSR[ 76 ][ 113 ],
   alphaCSR[ 76 ][ 114 ],
   alphaCSR[ 76 ][ 115 ],
   alphaCSR[ 76 ][ 116 ],
   alphaCSR[ 76 ][ 117 ],
   alphaCSR[ 76 ][ 118 ],
   alphaCSR[ 76 ][ 119 ],
   alphaCSR[ 76 ][ 120 ],
   alphaCSR[ 76 ][ 121 ],
   alphaCSR[ 76 ][ 122 ],
   alphaCSR[ 76 ][ 123 ],
   alphaCSR[ 76 ][ 124 ],
   alphaCSR[ 76 ][ 125 ],
   alphaCSR[ 76 ][ 126 ],
   alphaCSR[ 76 ][ 127 ],
   alphaCSR[ 76 ][ 128 ],
   alphaCSR[ 76 ][ 129 ],
   alphaCSR[ 76 ][ 130 ],
   alphaCSR[ 76 ][ 131 ],
   alphaCSR[ 76 ][ 132 ],
   alphaCSR[ 76 ][ 133 ],
   alphaCSR[ 76 ][ 134 ],
   alphaCSR[ 76 ][ 135 ],
   alphaCSR[ 76 ][ 136 ],
   alphaCSR[ 76 ][ 137 ],
   alphaCSR[ 76 ][ 138 ],
   alphaCSR[ 76 ][ 139 ],
   alphaCSR[ 76 ][ 140 ],
   alphaCSR[ 76 ][ 141 ],
   alphaCSR[ 76 ][ 142 ],
   alphaCSR[ 76 ][ 143 ],
   alphaCSR[ 76 ][ 144 ],
   alphaCSR[ 76 ][ 145 ],
   alphaCSR[ 76 ][ 146 ],
   alphaCSR[ 76 ][ 147 ],
   alphaCSR[ 76 ][ 148 ],
   alphaCSR[ 76 ][ 149 ],
   alphaCSR[ 76 ][ 150 ],
   alphaCSR[ 76 ][ 151 ],
   alphaCSR[ 76 ][ 152 ],
   alphaCSR[ 76 ][ 153 ],
   alphaCSR[ 76 ][ 154 ],
   alphaCSR[ 76 ][ 155 ],
   alphaCSR[ 76 ][ 156 ],
   alphaCSR[ 76 ][ 157 ],
   alphaCSR[ 76 ][ 158 ],
   alphaCSR[ 76 ][ 159 ],
   alphaCSR[ 76 ][ 160 ],
   alphaCSR[ 76 ][ 161 ],
   alphaCSR[ 76 ][ 162 ],
   alphaCSR[ 76 ][ 163 ],
   alphaCSR[ 76 ][ 164 ],
   alphaCSR[ 76 ][ 165 ],
   alphaCSR[ 76 ][ 166 ],
   alphaCSR[ 76 ][ 167 ],
   alphaCSR[ 76 ][ 168 ],
   alphaCSR[ 76 ][ 169 ],
   alphaCSR[ 76 ][ 170 ],
   alphaCSR[ 76 ][ 171 ],
   alphaCSR[ 76 ][ 172 ],
   alphaCSR[ 76 ][ 173 ],
   alphaCSR[ 76 ][ 174 ],
   alphaCSR[ 76 ][ 175 ],
   alphaCSR[ 76 ][ 176 ],
   alphaCSR[ 76 ][ 177 ],
   alphaCSR[ 76 ][ 178 ],
   alphaCSR[ 76 ][ 179 ],
   alphaCSR[ 76 ][ 180 ],
   alphaCSR[ 76 ][ 181 ],
   alphaCSR[ 76 ][ 182 ],
   alphaCSR[ 76 ][ 183 ],
   alphaCSR[ 76 ][ 184 ],
   alphaCSR[ 76 ][ 185 ],
   alphaCSR[ 76 ][ 186 ],
   alphaCSR[ 76 ][ 187 ],
   alphaCSR[ 76 ][ 188 ],
   alphaCSR[ 76 ][ 189 ],
   alphaCSR[ 76 ][ 190 ],
   alphaCSR[ 76 ][ 191 ],
   alphaCSR[ 76 ][ 192 ],
   alphaCSR[ 76 ][ 193 ],
   alphaCSR[ 76 ][ 194 ],
   alphaCSR[ 76 ][ 195 ],
   alphaCSR[ 76 ][ 196 ],
   alphaCSR[ 76 ][ 197 ],
   alphaCSR[ 76 ][ 198 ],
   alphaCSR[ 76 ][ 199 ],
   alphaCSR[ 76 ][ 200 ],
   alphaCSR[ 76 ][ 201 ],
   alphaCSR[ 76 ][ 202 ],
   alphaCSR[ 76 ][ 203 ],
   alphaCSR[ 76 ][ 204 ],
   alphaCSR[ 76 ][ 205 ],
   alphaCSR[ 76 ][ 206 ],
   alphaCSR[ 76 ][ 207 ],
   alphaCSR[ 76 ][ 208 ],
   alphaCSR[ 76 ][ 209 ],
   alphaCSR[ 76 ][ 210 ],
   alphaCSR[ 76 ][ 211 ],
   alphaCSR[ 76 ][ 212 ],
   alphaCSR[ 76 ][ 213 ],
   alphaCSR[ 76 ][ 214 ],
   alphaCSR[ 76 ][ 215 ],
   alphaCSR[ 76 ][ 216 ],
   alphaCSR[ 76 ][ 217 ],
   alphaCSR[ 76 ][ 218 ],
   alphaCSR[ 76 ][ 219 ],
   alphaCSR[ 76 ][ 220 ],
   alphaCSR[ 76 ][ 221 ],
   alphaCSR[ 76 ][ 222 ],
   alphaCSR[ 76 ][ 223 ],
   alphaCSR[ 76 ][ 224 ],
   alphaCSR[ 76 ][ 225 ],
   alphaCSR[ 76 ][ 226 ],
   alphaCSR[ 76 ][ 227 ],
   alphaCSR[ 76 ][ 228 ],
   alphaCSR[ 76 ][ 229 ],
   alphaCSR[ 76 ][ 230 ],
   alphaCSR[ 76 ][ 231 ],
   alphaCSR[ 76 ][ 232 ],
   alphaCSR[ 76 ][ 233 ],
   alphaCSR[ 76 ][ 234 ],
   alphaCSR[ 76 ][ 235 ],
   alphaCSR[ 76 ][ 236 ],
   alphaCSR[ 76 ][ 237 ],
   alphaCSR[ 76 ][ 238 ],
   alphaCSR[ 76 ][ 239 ],
   alphaCSR[ 76 ][ 240 ],
   alphaCSR[ 76 ][ 241 ],
   alphaCSR[ 76 ][ 242 ],
   alphaCSR[ 76 ][ 243 ],
   alphaCSR[ 76 ][ 244 ],
   alphaCSR[ 76 ][ 245 ],
   alphaCSR[ 76 ][ 246 ],
   alphaCSR[ 76 ][ 247 ],
   alphaCSR[ 76 ][ 248 ],
   alphaCSR[ 76 ][ 249 ],
   alphaCSR[ 76 ][ 250 ],
   alphaCSR[ 76 ][ 251 ],
   alphaCSR[ 76 ][ 252 ],
   alphaCSR[ 76 ][ 253 ],
   alphaCSR[ 76 ][ 254 ],
   alphaCSR[ 76 ][ 255 ],
   alphaCSR[ 76 ][ 256 ],
   alphaCSR[ 76 ][ 257 ],
   alphaCSR[ 76 ][ 258 ],
   alphaCSR[ 76 ][ 259 ],
   alphaCSR[ 76 ][ 260 ],
   alphaCSR[ 76 ][ 261 ],
   alphaCSR[ 76 ][ 262 ],
   alphaCSR[ 76 ][ 263 ],
   alphaCSR[ 76 ][ 264 ],
   alphaCSR[ 76 ][ 265 ],
   alphaCSR[ 76 ][ 266 ],
   alphaCSR[ 76 ][ 267 ],
   alphaCSR[ 76 ][ 268 ],
   alphaCSR[ 76 ][ 269 ],
   alphaCSR[ 76 ][ 270 ],
   alphaCSR[ 76 ][ 271 ],
   alphaCSR[ 76 ][ 272 ],
   alphaCSR[ 76 ][ 273 ],
   alphaCSR[ 76 ][ 274 ],
   alphaCSR[ 76 ][ 275 ],
   alphaCSR[ 76 ][ 276 ],
   alphaCSR[ 76 ][ 277 ],
   alphaCSR[ 76 ][ 278 ],
   alphaCSR[ 76 ][ 279 ],
   alphaCSR[ 76 ][ 280 ],
   alphaCSR[ 76 ][ 281 ],
   alphaCSR[ 76 ][ 282 ],
   alphaCSR[ 76 ][ 283 ],
   alphaCSR[ 76 ][ 284 ],
   alphaCSR[ 76 ][ 285 ],
   alphaCSR[ 76 ][ 286 ],
   alphaCSR[ 76 ][ 287 ],
   alphaCSR[ 76 ][ 288 ],
   alphaCSR[ 76 ][ 289 ],
   alphaCSR[ 76 ][ 290 ],
   alphaCSR[ 76 ][ 291 ],
   alphaCSR[ 76 ][ 292 ],
   alphaCSR[ 76 ][ 293 ],
   alphaCSR[ 76 ][ 294 ],
   alphaCSR[ 76 ][ 295 ],
   alphaCSR[ 76 ][ 296 ],
   alphaCSR[ 76 ][ 297 ],
   alphaCSR[ 76 ][ 298 ],
   alphaCSR[ 76 ][ 299 ],
   alphaCSR[ 76 ][ 300 ],
   alphaCSR[ 76 ][ 301 ],
   alphaCSR[ 76 ][ 302 ],
   alphaCSR[ 76 ][ 303 ],
   alphaCSR[ 76 ][ 304 ],
   alphaCSR[ 76 ][ 305 ],
   alphaCSR[ 76 ][ 306 ],
   alphaCSR[ 76 ][ 307 ],
   alphaCSR[ 76 ][ 308 ],
   alphaCSR[ 76 ][ 309 ],
   alphaCSR[ 76 ][ 310 ],
   alphaCSR[ 76 ][ 311 ],
   alphaCSR[ 76 ][ 312 ],
   alphaCSR[ 76 ][ 313 ],
   alphaCSR[ 76 ][ 314 ],
   alphaCSR[ 76 ][ 315 ],
   alphaCSR[ 76 ][ 316 ],
   alphaCSR[ 76 ][ 317 ],
   alphaCSR[ 76 ][ 318 ],
   alphaCSR[ 76 ][ 319 ],
   alphaCSR[ 76 ][ 320 ],
   alphaCSR[ 76 ][ 321 ],
   alphaCSR[ 76 ][ 322 ],
   alphaCSR[ 76 ][ 323 ],
   alphaCSR[ 76 ][ 324 ],
   alphaCSR[ 76 ][ 325 ],
   alphaCSR[ 76 ][ 326 ],
   alphaCSR[ 76 ][ 327 ],
   alphaCSR[ 76 ][ 328 ],
   alphaCSR[ 76 ][ 329 ],
   alphaCSR[ 76 ][ 330 ],
   alphaCSR[ 76 ][ 331 ],
   alphaCSR[ 76 ][ 332 ],
   alphaCSR[ 76 ][ 333 ],
   alphaCSR[ 76 ][ 334 ],
   alphaCSR[ 76 ][ 335 ],
   alphaCSR[ 76 ][ 336 ],
   alphaCSR[ 76 ][ 337 ],
   alphaCSR[ 76 ][ 338 ],
   alphaCSR[ 76 ][ 339 ],
   alphaCSR[ 76 ][ 340 ],
   alphaCSR[ 76 ][ 341 ],
   alphaCSR[ 76 ][ 342 ],
   alphaCSR[ 76 ][ 343 ],
   alphaCSR[ 76 ][ 344 ],
   alphaCSR[ 76 ][ 345 ],
   alphaCSR[ 76 ][ 346 ],
   alphaCSR[ 76 ][ 347 ],
   alphaCSR[ 76 ][ 348 ],
   alphaCSR[ 76 ][ 349 ],
   alphaCSR[ 76 ][ 350 ],
   alphaCSR[ 76 ][ 351 ],
   alphaCSR[ 76 ][ 352 ],
   alphaCSR[ 76 ][ 353 ],
   alphaCSR[ 76 ][ 354 ],
   alphaCSR[ 76 ][ 355 ],
   alphaCSR[ 76 ][ 356 ],
   alphaCSR[ 76 ][ 357 ],
   alphaCSR[ 76 ][ 358 ],
   alphaCSR[ 76 ][ 359 ],
   alphaCSR[ 76 ][ 360 ],
   alphaCSR[ 76 ][ 361 ],
   alphaCSR[ 76 ][ 362 ],
   alphaCSR[ 76 ][ 363 ],
   alphaCSR[ 76 ][ 364 ],
   alphaCSR[ 76 ][ 365 ],
   alphaCSR[ 76 ][ 366 ],
   alphaCSR[ 76 ][ 367 ],
   alphaCSR[ 76 ][ 368 ],
   alphaCSR[ 76 ][ 369 ],
   alphaCSR[ 76 ][ 370 ],
   alphaCSR[ 76 ][ 371 ],
   alphaCSR[ 76 ][ 372 ],
   alphaCSR[ 76 ][ 373 ],
   alphaCSR[ 76 ][ 374 ],
   alphaCSR[ 76 ][ 375 ],
   alphaCSR[ 76 ][ 376 ],
   alphaCSR[ 76 ][ 377 ],
   alphaCSR[ 76 ][ 378 ],
   alphaCSR[ 76 ][ 379 ],
   alphaCSR[ 76 ][ 380 ],
   alphaCSR[ 76 ][ 381 ],
   alphaCSR[ 76 ][ 382 ],
   alphaCSR[ 76 ][ 383 ],
   alphaCSR[ 77 ][ 0 ],
   alphaCSR[ 77 ][ 1 ],
   alphaCSR[ 77 ][ 2 ],
   alphaCSR[ 77 ][ 3 ],
   alphaCSR[ 77 ][ 4 ],
   alphaCSR[ 77 ][ 5 ],
   alphaCSR[ 77 ][ 6 ],
   alphaCSR[ 77 ][ 7 ],
   alphaCSR[ 77 ][ 8 ],
   alphaCSR[ 77 ][ 9 ],
   alphaCSR[ 77 ][ 10 ],
   alphaCSR[ 77 ][ 11 ],
   alphaCSR[ 77 ][ 12 ],
   alphaCSR[ 77 ][ 13 ],
   alphaCSR[ 77 ][ 14 ],
   alphaCSR[ 77 ][ 15 ],
   alphaCSR[ 77 ][ 16 ],
   alphaCSR[ 77 ][ 17 ],
   alphaCSR[ 77 ][ 18 ],
   alphaCSR[ 77 ][ 19 ],
   alphaCSR[ 77 ][ 20 ],
   alphaCSR[ 77 ][ 21 ],
   alphaCSR[ 77 ][ 22 ],
   alphaCSR[ 77 ][ 23 ],
   alphaCSR[ 77 ][ 24 ],
   alphaCSR[ 77 ][ 25 ],
   alphaCSR[ 77 ][ 26 ],
   alphaCSR[ 77 ][ 27 ],
   alphaCSR[ 77 ][ 28 ],
   alphaCSR[ 77 ][ 29 ],
   alphaCSR[ 77 ][ 30 ],
   alphaCSR[ 77 ][ 31 ],
   alphaCSR[ 77 ][ 32 ],
   alphaCSR[ 77 ][ 33 ],
   alphaCSR[ 77 ][ 34 ],
   alphaCSR[ 77 ][ 35 ],
   alphaCSR[ 77 ][ 36 ],
   alphaCSR[ 77 ][ 37 ],
   alphaCSR[ 77 ][ 38 ],
   alphaCSR[ 77 ][ 39 ],
   alphaCSR[ 77 ][ 40 ],
   alphaCSR[ 77 ][ 41 ],
   alphaCSR[ 77 ][ 42 ],
   alphaCSR[ 77 ][ 43 ],
   alphaCSR[ 77 ][ 44 ],
   alphaCSR[ 77 ][ 45 ],
   alphaCSR[ 77 ][ 46 ],
   alphaCSR[ 77 ][ 47 ],
   alphaCSR[ 77 ][ 48 ],
   alphaCSR[ 77 ][ 49 ],
   alphaCSR[ 77 ][ 50 ],
   alphaCSR[ 77 ][ 51 ],
   alphaCSR[ 77 ][ 52 ],
   alphaCSR[ 77 ][ 53 ],
   alphaCSR[ 77 ][ 54 ],
   alphaCSR[ 77 ][ 55 ],
   alphaCSR[ 77 ][ 56 ],
   alphaCSR[ 77 ][ 57 ],
   alphaCSR[ 77 ][ 58 ],
   alphaCSR[ 77 ][ 59 ],
   alphaCSR[ 77 ][ 60 ],
   alphaCSR[ 77 ][ 61 ],
   alphaCSR[ 77 ][ 62 ],
   alphaCSR[ 77 ][ 63 ],
   alphaCSR[ 77 ][ 64 ],
   alphaCSR[ 77 ][ 65 ],
   alphaCSR[ 77 ][ 66 ],
   alphaCSR[ 77 ][ 67 ],
   alphaCSR[ 77 ][ 68 ],
   alphaCSR[ 77 ][ 69 ],
   alphaCSR[ 77 ][ 70 ],
   alphaCSR[ 77 ][ 71 ],
   alphaCSR[ 77 ][ 72 ],
   alphaCSR[ 77 ][ 73 ],
   alphaCSR[ 77 ][ 74 ],
   alphaCSR[ 77 ][ 75 ],
   alphaCSR[ 77 ][ 76 ],
   alphaCSR[ 77 ][ 77 ],
   alphaCSR[ 77 ][ 78 ],
   alphaCSR[ 77 ][ 79 ],
   alphaCSR[ 77 ][ 80 ],
   alphaCSR[ 77 ][ 81 ],
   alphaCSR[ 77 ][ 82 ],
   alphaCSR[ 77 ][ 83 ],
   alphaCSR[ 77 ][ 84 ],
   alphaCSR[ 77 ][ 85 ],
   alphaCSR[ 77 ][ 86 ],
   alphaCSR[ 77 ][ 87 ],
   alphaCSR[ 77 ][ 88 ],
   alphaCSR[ 77 ][ 89 ],
   alphaCSR[ 77 ][ 90 ],
   alphaCSR[ 77 ][ 91 ],
   alphaCSR[ 77 ][ 92 ],
   alphaCSR[ 77 ][ 93 ],
   alphaCSR[ 77 ][ 94 ],
   alphaCSR[ 77 ][ 95 ],
   alphaCSR[ 77 ][ 96 ],
   alphaCSR[ 77 ][ 97 ],
   alphaCSR[ 77 ][ 98 ],
   alphaCSR[ 77 ][ 99 ],
   alphaCSR[ 77 ][ 100 ],
   alphaCSR[ 77 ][ 101 ],
   alphaCSR[ 77 ][ 102 ],
   alphaCSR[ 77 ][ 103 ],
   alphaCSR[ 77 ][ 104 ],
   alphaCSR[ 77 ][ 105 ],
   alphaCSR[ 77 ][ 106 ],
   alphaCSR[ 77 ][ 107 ],
   alphaCSR[ 77 ][ 108 ],
   alphaCSR[ 77 ][ 109 ],
   alphaCSR[ 77 ][ 110 ],
   alphaCSR[ 77 ][ 111 ],
   alphaCSR[ 77 ][ 112 ],
   alphaCSR[ 77 ][ 113 ],
   alphaCSR[ 77 ][ 114 ],
   alphaCSR[ 77 ][ 115 ],
   alphaCSR[ 77 ][ 116 ],
   alphaCSR[ 77 ][ 117 ],
   alphaCSR[ 77 ][ 118 ],
   alphaCSR[ 77 ][ 119 ],
   alphaCSR[ 77 ][ 120 ],
   alphaCSR[ 77 ][ 121 ],
   alphaCSR[ 77 ][ 122 ],
   alphaCSR[ 77 ][ 123 ],
   alphaCSR[ 77 ][ 124 ],
   alphaCSR[ 77 ][ 125 ],
   alphaCSR[ 77 ][ 126 ],
   alphaCSR[ 77 ][ 127 ],
   alphaCSR[ 77 ][ 128 ],
   alphaCSR[ 77 ][ 129 ],
   alphaCSR[ 77 ][ 130 ],
   alphaCSR[ 77 ][ 131 ],
   alphaCSR[ 77 ][ 132 ],
   alphaCSR[ 77 ][ 133 ],
   alphaCSR[ 77 ][ 134 ],
   alphaCSR[ 77 ][ 135 ],
   alphaCSR[ 77 ][ 136 ],
   alphaCSR[ 77 ][ 137 ],
   alphaCSR[ 77 ][ 138 ],
   alphaCSR[ 77 ][ 139 ],
   alphaCSR[ 77 ][ 140 ],
   alphaCSR[ 77 ][ 141 ],
   alphaCSR[ 77 ][ 142 ],
   alphaCSR[ 77 ][ 143 ],
   alphaCSR[ 77 ][ 144 ],
   alphaCSR[ 77 ][ 145 ],
   alphaCSR[ 77 ][ 146 ],
   alphaCSR[ 77 ][ 147 ],
   alphaCSR[ 77 ][ 148 ],
   alphaCSR[ 77 ][ 149 ],
   alphaCSR[ 77 ][ 150 ],
   alphaCSR[ 77 ][ 151 ],
   alphaCSR[ 77 ][ 152 ],
   alphaCSR[ 77 ][ 153 ],
   alphaCSR[ 77 ][ 154 ],
   alphaCSR[ 77 ][ 155 ],
   alphaCSR[ 77 ][ 156 ],
   alphaCSR[ 77 ][ 157 ],
   alphaCSR[ 77 ][ 158 ],
   alphaCSR[ 77 ][ 159 ],
   alphaCSR[ 77 ][ 160 ],
   alphaCSR[ 77 ][ 161 ],
   alphaCSR[ 77 ][ 162 ],
   alphaCSR[ 77 ][ 163 ],
   alphaCSR[ 77 ][ 164 ],
   alphaCSR[ 77 ][ 165 ],
   alphaCSR[ 77 ][ 166 ],
   alphaCSR[ 77 ][ 167 ],
   alphaCSR[ 77 ][ 168 ],
   alphaCSR[ 77 ][ 169 ],
   alphaCSR[ 77 ][ 170 ],
   alphaCSR[ 77 ][ 171 ],
   alphaCSR[ 77 ][ 172 ],
   alphaCSR[ 77 ][ 173 ],
   alphaCSR[ 77 ][ 174 ],
   alphaCSR[ 77 ][ 175 ],
   alphaCSR[ 77 ][ 176 ],
   alphaCSR[ 77 ][ 177 ],
   alphaCSR[ 77 ][ 178 ],
   alphaCSR[ 77 ][ 179 ],
   alphaCSR[ 77 ][ 180 ],
   alphaCSR[ 77 ][ 181 ],
   alphaCSR[ 77 ][ 182 ],
   alphaCSR[ 77 ][ 183 ],
   alphaCSR[ 77 ][ 184 ],
   alphaCSR[ 77 ][ 185 ],
   alphaCSR[ 77 ][ 186 ],
   alphaCSR[ 77 ][ 187 ],
   alphaCSR[ 77 ][ 188 ],
   alphaCSR[ 77 ][ 189 ],
   alphaCSR[ 77 ][ 190 ],
   alphaCSR[ 77 ][ 191 ],
   alphaCSR[ 77 ][ 192 ],
   alphaCSR[ 77 ][ 193 ],
   alphaCSR[ 77 ][ 194 ],
   alphaCSR[ 77 ][ 195 ],
   alphaCSR[ 77 ][ 196 ],
   alphaCSR[ 77 ][ 197 ],
   alphaCSR[ 77 ][ 198 ],
   alphaCSR[ 77 ][ 199 ],
   alphaCSR[ 77 ][ 200 ],
   alphaCSR[ 77 ][ 201 ],
   alphaCSR[ 77 ][ 202 ],
   alphaCSR[ 77 ][ 203 ],
   alphaCSR[ 77 ][ 204 ],
   alphaCSR[ 77 ][ 205 ],
   alphaCSR[ 77 ][ 206 ],
   alphaCSR[ 77 ][ 207 ],
   alphaCSR[ 77 ][ 208 ],
   alphaCSR[ 77 ][ 209 ],
   alphaCSR[ 77 ][ 210 ],
   alphaCSR[ 77 ][ 211 ],
   alphaCSR[ 77 ][ 212 ],
   alphaCSR[ 77 ][ 213 ],
   alphaCSR[ 77 ][ 214 ],
   alphaCSR[ 77 ][ 215 ],
   alphaCSR[ 77 ][ 216 ],
   alphaCSR[ 77 ][ 217 ],
   alphaCSR[ 77 ][ 218 ],
   alphaCSR[ 77 ][ 219 ],
   alphaCSR[ 77 ][ 220 ],
   alphaCSR[ 77 ][ 221 ],
   alphaCSR[ 77 ][ 222 ],
   alphaCSR[ 77 ][ 223 ],
   alphaCSR[ 77 ][ 224 ],
   alphaCSR[ 77 ][ 225 ],
   alphaCSR[ 77 ][ 226 ],
   alphaCSR[ 77 ][ 227 ],
   alphaCSR[ 77 ][ 228 ],
   alphaCSR[ 77 ][ 229 ],
   alphaCSR[ 77 ][ 230 ],
   alphaCSR[ 77 ][ 231 ],
   alphaCSR[ 77 ][ 232 ],
   alphaCSR[ 77 ][ 233 ],
   alphaCSR[ 77 ][ 234 ],
   alphaCSR[ 77 ][ 235 ],
   alphaCSR[ 77 ][ 236 ],
   alphaCSR[ 77 ][ 237 ],
   alphaCSR[ 77 ][ 238 ],
   alphaCSR[ 77 ][ 239 ],
   alphaCSR[ 77 ][ 240 ],
   alphaCSR[ 77 ][ 241 ],
   alphaCSR[ 77 ][ 242 ],
   alphaCSR[ 77 ][ 243 ],
   alphaCSR[ 77 ][ 244 ],
   alphaCSR[ 77 ][ 245 ],
   alphaCSR[ 77 ][ 246 ],
   alphaCSR[ 77 ][ 247 ],
   alphaCSR[ 77 ][ 248 ],
   alphaCSR[ 77 ][ 249 ],
   alphaCSR[ 77 ][ 250 ],
   alphaCSR[ 77 ][ 251 ],
   alphaCSR[ 77 ][ 252 ],
   alphaCSR[ 77 ][ 253 ],
   alphaCSR[ 77 ][ 254 ],
   alphaCSR[ 77 ][ 255 ],
   alphaCSR[ 77 ][ 256 ],
   alphaCSR[ 77 ][ 257 ],
   alphaCSR[ 77 ][ 258 ],
   alphaCSR[ 77 ][ 259 ],
   alphaCSR[ 77 ][ 260 ],
   alphaCSR[ 77 ][ 261 ],
   alphaCSR[ 77 ][ 262 ],
   alphaCSR[ 77 ][ 263 ],
   alphaCSR[ 77 ][ 264 ],
   alphaCSR[ 77 ][ 265 ],
   alphaCSR[ 77 ][ 266 ],
   alphaCSR[ 77 ][ 267 ],
   alphaCSR[ 77 ][ 268 ],
   alphaCSR[ 77 ][ 269 ],
   alphaCSR[ 77 ][ 270 ],
   alphaCSR[ 77 ][ 271 ],
   alphaCSR[ 77 ][ 272 ],
   alphaCSR[ 77 ][ 273 ],
   alphaCSR[ 77 ][ 274 ],
   alphaCSR[ 77 ][ 275 ],
   alphaCSR[ 77 ][ 276 ],
   alphaCSR[ 77 ][ 277 ],
   alphaCSR[ 77 ][ 278 ],
   alphaCSR[ 77 ][ 279 ],
   alphaCSR[ 77 ][ 280 ],
   alphaCSR[ 77 ][ 281 ],
   alphaCSR[ 77 ][ 282 ],
   alphaCSR[ 77 ][ 283 ],
   alphaCSR[ 77 ][ 284 ],
   alphaCSR[ 77 ][ 285 ],
   alphaCSR[ 77 ][ 286 ],
   alphaCSR[ 77 ][ 287 ],
   alphaCSR[ 77 ][ 288 ],
   alphaCSR[ 77 ][ 289 ],
   alphaCSR[ 77 ][ 290 ],
   alphaCSR[ 77 ][ 291 ],
   alphaCSR[ 77 ][ 292 ],
   alphaCSR[ 77 ][ 293 ],
   alphaCSR[ 77 ][ 294 ],
   alphaCSR[ 77 ][ 295 ],
   alphaCSR[ 77 ][ 296 ],
   alphaCSR[ 77 ][ 297 ],
   alphaCSR[ 77 ][ 298 ],
   alphaCSR[ 77 ][ 299 ],
   alphaCSR[ 77 ][ 300 ],
   alphaCSR[ 77 ][ 301 ],
   alphaCSR[ 77 ][ 302 ],
   alphaCSR[ 77 ][ 303 ],
   alphaCSR[ 77 ][ 304 ],
   alphaCSR[ 77 ][ 305 ],
   alphaCSR[ 77 ][ 306 ],
   alphaCSR[ 77 ][ 307 ],
   alphaCSR[ 77 ][ 308 ],
   alphaCSR[ 77 ][ 309 ],
   alphaCSR[ 77 ][ 310 ],
   alphaCSR[ 77 ][ 311 ],
   alphaCSR[ 77 ][ 312 ],
   alphaCSR[ 77 ][ 313 ],
   alphaCSR[ 77 ][ 314 ],
   alphaCSR[ 77 ][ 315 ],
   alphaCSR[ 77 ][ 316 ],
   alphaCSR[ 77 ][ 317 ],
   alphaCSR[ 77 ][ 318 ],
   alphaCSR[ 77 ][ 319 ],
   alphaCSR[ 77 ][ 320 ],
   alphaCSR[ 77 ][ 321 ],
   alphaCSR[ 77 ][ 322 ],
   alphaCSR[ 77 ][ 323 ],
   alphaCSR[ 77 ][ 324 ],
   alphaCSR[ 77 ][ 325 ],
   alphaCSR[ 77 ][ 326 ],
   alphaCSR[ 77 ][ 327 ],
   alphaCSR[ 77 ][ 328 ],
   alphaCSR[ 77 ][ 329 ],
   alphaCSR[ 77 ][ 330 ],
   alphaCSR[ 77 ][ 331 ],
   alphaCSR[ 77 ][ 332 ],
   alphaCSR[ 77 ][ 333 ],
   alphaCSR[ 77 ][ 334 ],
   alphaCSR[ 77 ][ 335 ],
   alphaCSR[ 77 ][ 336 ],
   alphaCSR[ 77 ][ 337 ],
   alphaCSR[ 77 ][ 338 ],
   alphaCSR[ 77 ][ 339 ],
   alphaCSR[ 77 ][ 340 ],
   alphaCSR[ 77 ][ 341 ],
   alphaCSR[ 77 ][ 342 ],
   alphaCSR[ 77 ][ 343 ],
   alphaCSR[ 77 ][ 344 ],
   alphaCSR[ 77 ][ 345 ],
   alphaCSR[ 77 ][ 346 ],
   alphaCSR[ 77 ][ 347 ],
   alphaCSR[ 77 ][ 348 ],
   alphaCSR[ 77 ][ 349 ],
   alphaCSR[ 77 ][ 350 ],
   alphaCSR[ 77 ][ 351 ],
   alphaCSR[ 77 ][ 352 ],
   alphaCSR[ 77 ][ 353 ],
   alphaCSR[ 77 ][ 354 ],
   alphaCSR[ 77 ][ 355 ],
   alphaCSR[ 77 ][ 356 ],
   alphaCSR[ 77 ][ 357 ],
   alphaCSR[ 77 ][ 358 ],
   alphaCSR[ 77 ][ 359 ],
   alphaCSR[ 77 ][ 360 ],
   alphaCSR[ 77 ][ 361 ],
   alphaCSR[ 77 ][ 362 ],
   alphaCSR[ 77 ][ 363 ],
   alphaCSR[ 77 ][ 364 ],
   alphaCSR[ 77 ][ 365 ],
   alphaCSR[ 77 ][ 366 ],
   alphaCSR[ 77 ][ 367 ],
   alphaCSR[ 77 ][ 368 ],
   alphaCSR[ 77 ][ 369 ],
   alphaCSR[ 77 ][ 370 ],
   alphaCSR[ 77 ][ 371 ],
   alphaCSR[ 77 ][ 372 ],
   alphaCSR[ 77 ][ 373 ],
   alphaCSR[ 77 ][ 374 ],
   alphaCSR[ 77 ][ 375 ],
   alphaCSR[ 77 ][ 376 ],
   alphaCSR[ 77 ][ 377 ],
   alphaCSR[ 77 ][ 378 ],
   alphaCSR[ 77 ][ 379 ],
   alphaCSR[ 77 ][ 380 ],
   alphaCSR[ 77 ][ 381 ],
   alphaCSR[ 77 ][ 382 ],
   alphaCSR[ 77 ][ 383 ],
   alphaCSR[ 78 ][ 0 ],
   alphaCSR[ 78 ][ 1 ],
   alphaCSR[ 78 ][ 2 ],
   alphaCSR[ 78 ][ 3 ],
   alphaCSR[ 78 ][ 4 ],
   alphaCSR[ 78 ][ 5 ],
   alphaCSR[ 78 ][ 6 ],
   alphaCSR[ 78 ][ 7 ],
   alphaCSR[ 78 ][ 8 ],
   alphaCSR[ 78 ][ 9 ],
   alphaCSR[ 78 ][ 10 ],
   alphaCSR[ 78 ][ 11 ],
   alphaCSR[ 78 ][ 12 ],
   alphaCSR[ 78 ][ 13 ],
   alphaCSR[ 78 ][ 14 ],
   alphaCSR[ 78 ][ 15 ],
   alphaCSR[ 78 ][ 16 ],
   alphaCSR[ 78 ][ 17 ],
   alphaCSR[ 78 ][ 18 ],
   alphaCSR[ 78 ][ 19 ],
   alphaCSR[ 78 ][ 20 ],
   alphaCSR[ 78 ][ 21 ],
   alphaCSR[ 78 ][ 22 ],
   alphaCSR[ 78 ][ 23 ],
   alphaCSR[ 78 ][ 24 ],
   alphaCSR[ 78 ][ 25 ],
   alphaCSR[ 78 ][ 26 ],
   alphaCSR[ 78 ][ 27 ],
   alphaCSR[ 78 ][ 28 ],
   alphaCSR[ 78 ][ 29 ],
   alphaCSR[ 78 ][ 30 ],
   alphaCSR[ 78 ][ 31 ],
   alphaCSR[ 78 ][ 32 ],
   alphaCSR[ 78 ][ 33 ],
   alphaCSR[ 78 ][ 34 ],
   alphaCSR[ 78 ][ 35 ],
   alphaCSR[ 78 ][ 36 ],
   alphaCSR[ 78 ][ 37 ],
   alphaCSR[ 78 ][ 38 ],
   alphaCSR[ 78 ][ 39 ],
   alphaCSR[ 78 ][ 40 ],
   alphaCSR[ 78 ][ 41 ],
   alphaCSR[ 78 ][ 42 ],
   alphaCSR[ 78 ][ 43 ],
   alphaCSR[ 78 ][ 44 ],
   alphaCSR[ 78 ][ 45 ],
   alphaCSR[ 78 ][ 46 ],
   alphaCSR[ 78 ][ 47 ],
   alphaCSR[ 78 ][ 48 ],
   alphaCSR[ 78 ][ 49 ],
   alphaCSR[ 78 ][ 50 ],
   alphaCSR[ 78 ][ 51 ],
   alphaCSR[ 78 ][ 52 ],
   alphaCSR[ 78 ][ 53 ],
   alphaCSR[ 78 ][ 54 ],
   alphaCSR[ 78 ][ 55 ],
   alphaCSR[ 78 ][ 56 ],
   alphaCSR[ 78 ][ 57 ],
   alphaCSR[ 78 ][ 58 ],
   alphaCSR[ 78 ][ 59 ],
   alphaCSR[ 78 ][ 60 ],
   alphaCSR[ 78 ][ 61 ],
   alphaCSR[ 78 ][ 62 ],
   alphaCSR[ 78 ][ 63 ],
   alphaCSR[ 78 ][ 64 ],
   alphaCSR[ 78 ][ 65 ],
   alphaCSR[ 78 ][ 66 ],
   alphaCSR[ 78 ][ 67 ],
   alphaCSR[ 78 ][ 68 ],
   alphaCSR[ 78 ][ 69 ],
   alphaCSR[ 78 ][ 70 ],
   alphaCSR[ 78 ][ 71 ],
   alphaCSR[ 78 ][ 72 ],
   alphaCSR[ 78 ][ 73 ],
   alphaCSR[ 78 ][ 74 ],
   alphaCSR[ 78 ][ 75 ],
   alphaCSR[ 78 ][ 76 ],
   alphaCSR[ 78 ][ 77 ],
   alphaCSR[ 78 ][ 78 ],
   alphaCSR[ 78 ][ 79 ],
   alphaCSR[ 78 ][ 80 ],
   alphaCSR[ 78 ][ 81 ],
   alphaCSR[ 78 ][ 82 ],
   alphaCSR[ 78 ][ 83 ],
   alphaCSR[ 78 ][ 84 ],
   alphaCSR[ 78 ][ 85 ],
   alphaCSR[ 78 ][ 86 ],
   alphaCSR[ 78 ][ 87 ],
   alphaCSR[ 78 ][ 88 ],
   alphaCSR[ 78 ][ 89 ],
   alphaCSR[ 78 ][ 90 ],
   alphaCSR[ 78 ][ 91 ],
   alphaCSR[ 78 ][ 92 ],
   alphaCSR[ 78 ][ 93 ],
   alphaCSR[ 78 ][ 94 ],
   alphaCSR[ 78 ][ 95 ],
   alphaCSR[ 78 ][ 96 ],
   alphaCSR[ 78 ][ 97 ],
   alphaCSR[ 78 ][ 98 ],
   alphaCSR[ 78 ][ 99 ],
   alphaCSR[ 78 ][ 100 ],
   alphaCSR[ 78 ][ 101 ],
   alphaCSR[ 78 ][ 102 ],
   alphaCSR[ 78 ][ 103 ],
   alphaCSR[ 78 ][ 104 ],
   alphaCSR[ 78 ][ 105 ],
   alphaCSR[ 78 ][ 106 ],
   alphaCSR[ 78 ][ 107 ],
   alphaCSR[ 78 ][ 108 ],
   alphaCSR[ 78 ][ 109 ],
   alphaCSR[ 78 ][ 110 ],
   alphaCSR[ 78 ][ 111 ],
   alphaCSR[ 78 ][ 112 ],
   alphaCSR[ 78 ][ 113 ],
   alphaCSR[ 78 ][ 114 ],
   alphaCSR[ 78 ][ 115 ],
   alphaCSR[ 78 ][ 116 ],
   alphaCSR[ 78 ][ 117 ],
   alphaCSR[ 78 ][ 118 ],
   alphaCSR[ 78 ][ 119 ],
   alphaCSR[ 78 ][ 120 ],
   alphaCSR[ 78 ][ 121 ],
   alphaCSR[ 78 ][ 122 ],
   alphaCSR[ 78 ][ 123 ],
   alphaCSR[ 78 ][ 124 ],
   alphaCSR[ 78 ][ 125 ],
   alphaCSR[ 78 ][ 126 ],
   alphaCSR[ 78 ][ 127 ],
   alphaCSR[ 78 ][ 128 ],
   alphaCSR[ 78 ][ 129 ],
   alphaCSR[ 78 ][ 130 ],
   alphaCSR[ 78 ][ 131 ],
   alphaCSR[ 78 ][ 132 ],
   alphaCSR[ 78 ][ 133 ],
   alphaCSR[ 78 ][ 134 ],
   alphaCSR[ 78 ][ 135 ],
   alphaCSR[ 78 ][ 136 ],
   alphaCSR[ 78 ][ 137 ],
   alphaCSR[ 78 ][ 138 ],
   alphaCSR[ 78 ][ 139 ],
   alphaCSR[ 78 ][ 140 ],
   alphaCSR[ 78 ][ 141 ],
   alphaCSR[ 78 ][ 142 ],
   alphaCSR[ 78 ][ 143 ],
   alphaCSR[ 78 ][ 144 ],
   alphaCSR[ 78 ][ 145 ],
   alphaCSR[ 78 ][ 146 ],
   alphaCSR[ 78 ][ 147 ],
   alphaCSR[ 78 ][ 148 ],
   alphaCSR[ 78 ][ 149 ],
   alphaCSR[ 78 ][ 150 ],
   alphaCSR[ 78 ][ 151 ],
   alphaCSR[ 78 ][ 152 ],
   alphaCSR[ 78 ][ 153 ],
   alphaCSR[ 78 ][ 154 ],
   alphaCSR[ 78 ][ 155 ],
   alphaCSR[ 78 ][ 156 ],
   alphaCSR[ 78 ][ 157 ],
   alphaCSR[ 78 ][ 158 ],
   alphaCSR[ 78 ][ 159 ],
   alphaCSR[ 78 ][ 160 ],
   alphaCSR[ 78 ][ 161 ],
   alphaCSR[ 78 ][ 162 ],
   alphaCSR[ 78 ][ 163 ],
   alphaCSR[ 78 ][ 164 ],
   alphaCSR[ 78 ][ 165 ],
   alphaCSR[ 78 ][ 166 ],
   alphaCSR[ 78 ][ 167 ],
   alphaCSR[ 78 ][ 168 ],
   alphaCSR[ 78 ][ 169 ],
   alphaCSR[ 78 ][ 170 ],
   alphaCSR[ 78 ][ 171 ],
   alphaCSR[ 78 ][ 172 ],
   alphaCSR[ 78 ][ 173 ],
   alphaCSR[ 78 ][ 174 ],
   alphaCSR[ 78 ][ 175 ],
   alphaCSR[ 78 ][ 176 ],
   alphaCSR[ 78 ][ 177 ],
   alphaCSR[ 78 ][ 178 ],
   alphaCSR[ 78 ][ 179 ],
   alphaCSR[ 78 ][ 180 ],
   alphaCSR[ 78 ][ 181 ],
   alphaCSR[ 78 ][ 182 ],
   alphaCSR[ 78 ][ 183 ],
   alphaCSR[ 78 ][ 184 ],
   alphaCSR[ 78 ][ 185 ],
   alphaCSR[ 78 ][ 186 ],
   alphaCSR[ 78 ][ 187 ],
   alphaCSR[ 78 ][ 188 ],
   alphaCSR[ 78 ][ 189 ],
   alphaCSR[ 78 ][ 190 ],
   alphaCSR[ 78 ][ 191 ],
   alphaCSR[ 78 ][ 192 ],
   alphaCSR[ 78 ][ 193 ],
   alphaCSR[ 78 ][ 194 ],
   alphaCSR[ 78 ][ 195 ],
   alphaCSR[ 78 ][ 196 ],
   alphaCSR[ 78 ][ 197 ],
   alphaCSR[ 78 ][ 198 ],
   alphaCSR[ 78 ][ 199 ],
   alphaCSR[ 78 ][ 200 ],
   alphaCSR[ 78 ][ 201 ],
   alphaCSR[ 78 ][ 202 ],
   alphaCSR[ 78 ][ 203 ],
   alphaCSR[ 78 ][ 204 ],
   alphaCSR[ 78 ][ 205 ],
   alphaCSR[ 78 ][ 206 ],
   alphaCSR[ 78 ][ 207 ],
   alphaCSR[ 78 ][ 208 ],
   alphaCSR[ 78 ][ 209 ],
   alphaCSR[ 78 ][ 210 ],
   alphaCSR[ 78 ][ 211 ],
   alphaCSR[ 78 ][ 212 ],
   alphaCSR[ 78 ][ 213 ],
   alphaCSR[ 78 ][ 214 ],
   alphaCSR[ 78 ][ 215 ],
   alphaCSR[ 78 ][ 216 ],
   alphaCSR[ 78 ][ 217 ],
   alphaCSR[ 78 ][ 218 ],
   alphaCSR[ 78 ][ 219 ],
   alphaCSR[ 78 ][ 220 ],
   alphaCSR[ 78 ][ 221 ],
   alphaCSR[ 78 ][ 222 ],
   alphaCSR[ 78 ][ 223 ],
   alphaCSR[ 78 ][ 224 ],
   alphaCSR[ 78 ][ 225 ],
   alphaCSR[ 78 ][ 226 ],
   alphaCSR[ 78 ][ 227 ],
   alphaCSR[ 78 ][ 228 ],
   alphaCSR[ 78 ][ 229 ],
   alphaCSR[ 78 ][ 230 ],
   alphaCSR[ 78 ][ 231 ],
   alphaCSR[ 78 ][ 232 ],
   alphaCSR[ 78 ][ 233 ],
   alphaCSR[ 78 ][ 234 ],
   alphaCSR[ 78 ][ 235 ],
   alphaCSR[ 78 ][ 236 ],
   alphaCSR[ 78 ][ 237 ],
   alphaCSR[ 78 ][ 238 ],
   alphaCSR[ 78 ][ 239 ],
   alphaCSR[ 78 ][ 240 ],
   alphaCSR[ 78 ][ 241 ],
   alphaCSR[ 78 ][ 242 ],
   alphaCSR[ 78 ][ 243 ],
   alphaCSR[ 78 ][ 244 ],
   alphaCSR[ 78 ][ 245 ],
   alphaCSR[ 78 ][ 246 ],
   alphaCSR[ 78 ][ 247 ],
   alphaCSR[ 78 ][ 248 ],
   alphaCSR[ 78 ][ 249 ],
   alphaCSR[ 78 ][ 250 ],
   alphaCSR[ 78 ][ 251 ],
   alphaCSR[ 78 ][ 252 ],
   alphaCSR[ 78 ][ 253 ],
   alphaCSR[ 78 ][ 254 ],
   alphaCSR[ 78 ][ 255 ],
   alphaCSR[ 78 ][ 256 ],
   alphaCSR[ 78 ][ 257 ],
   alphaCSR[ 78 ][ 258 ],
   alphaCSR[ 78 ][ 259 ],
   alphaCSR[ 78 ][ 260 ],
   alphaCSR[ 78 ][ 261 ],
   alphaCSR[ 78 ][ 262 ],
   alphaCSR[ 78 ][ 263 ],
   alphaCSR[ 78 ][ 264 ],
   alphaCSR[ 78 ][ 265 ],
   alphaCSR[ 78 ][ 266 ],
   alphaCSR[ 78 ][ 267 ],
   alphaCSR[ 78 ][ 268 ],
   alphaCSR[ 78 ][ 269 ],
   alphaCSR[ 78 ][ 270 ],
   alphaCSR[ 78 ][ 271 ],
   alphaCSR[ 78 ][ 272 ],
   alphaCSR[ 78 ][ 273 ],
   alphaCSR[ 78 ][ 274 ],
   alphaCSR[ 78 ][ 275 ],
   alphaCSR[ 78 ][ 276 ],
   alphaCSR[ 78 ][ 277 ],
   alphaCSR[ 78 ][ 278 ],
   alphaCSR[ 78 ][ 279 ],
   alphaCSR[ 78 ][ 280 ],
   alphaCSR[ 78 ][ 281 ],
   alphaCSR[ 78 ][ 282 ],
   alphaCSR[ 78 ][ 283 ],
   alphaCSR[ 78 ][ 284 ],
   alphaCSR[ 78 ][ 285 ],
   alphaCSR[ 78 ][ 286 ],
   alphaCSR[ 78 ][ 287 ],
   alphaCSR[ 78 ][ 288 ],
   alphaCSR[ 78 ][ 289 ],
   alphaCSR[ 78 ][ 290 ],
   alphaCSR[ 78 ][ 291 ],
   alphaCSR[ 78 ][ 292 ],
   alphaCSR[ 78 ][ 293 ],
   alphaCSR[ 78 ][ 294 ],
   alphaCSR[ 78 ][ 295 ],
   alphaCSR[ 78 ][ 296 ],
   alphaCSR[ 78 ][ 297 ],
   alphaCSR[ 78 ][ 298 ],
   alphaCSR[ 78 ][ 299 ],
   alphaCSR[ 78 ][ 300 ],
   alphaCSR[ 78 ][ 301 ],
   alphaCSR[ 78 ][ 302 ],
   alphaCSR[ 78 ][ 303 ],
   alphaCSR[ 78 ][ 304 ],
   alphaCSR[ 78 ][ 305 ],
   alphaCSR[ 78 ][ 306 ],
   alphaCSR[ 78 ][ 307 ],
   alphaCSR[ 78 ][ 308 ],
   alphaCSR[ 78 ][ 309 ],
   alphaCSR[ 78 ][ 310 ],
   alphaCSR[ 78 ][ 311 ],
   alphaCSR[ 78 ][ 312 ],
   alphaCSR[ 78 ][ 313 ],
   alphaCSR[ 78 ][ 314 ],
   alphaCSR[ 78 ][ 315 ],
   alphaCSR[ 78 ][ 316 ],
   alphaCSR[ 78 ][ 317 ],
   alphaCSR[ 78 ][ 318 ],
   alphaCSR[ 78 ][ 319 ],
   alphaCSR[ 78 ][ 320 ],
   alphaCSR[ 78 ][ 321 ],
   alphaCSR[ 78 ][ 322 ],
   alphaCSR[ 78 ][ 323 ],
   alphaCSR[ 78 ][ 324 ],
   alphaCSR[ 78 ][ 325 ],
   alphaCSR[ 78 ][ 326 ],
   alphaCSR[ 78 ][ 327 ],
   alphaCSR[ 78 ][ 328 ],
   alphaCSR[ 78 ][ 329 ],
   alphaCSR[ 78 ][ 330 ],
   alphaCSR[ 78 ][ 331 ],
   alphaCSR[ 78 ][ 332 ],
   alphaCSR[ 78 ][ 333 ],
   alphaCSR[ 78 ][ 334 ],
   alphaCSR[ 78 ][ 335 ],
   alphaCSR[ 78 ][ 336 ],
   alphaCSR[ 78 ][ 337 ],
   alphaCSR[ 78 ][ 338 ],
   alphaCSR[ 78 ][ 339 ],
   alphaCSR[ 78 ][ 340 ],
   alphaCSR[ 78 ][ 341 ],
   alphaCSR[ 78 ][ 342 ],
   alphaCSR[ 78 ][ 343 ],
   alphaCSR[ 78 ][ 344 ],
   alphaCSR[ 78 ][ 345 ],
   alphaCSR[ 78 ][ 346 ],
   alphaCSR[ 78 ][ 347 ],
   alphaCSR[ 78 ][ 348 ],
   alphaCSR[ 78 ][ 349 ],
   alphaCSR[ 78 ][ 350 ],
   alphaCSR[ 78 ][ 351 ],
   alphaCSR[ 78 ][ 352 ],
   alphaCSR[ 78 ][ 353 ],
   alphaCSR[ 78 ][ 354 ],
   alphaCSR[ 78 ][ 355 ],
   alphaCSR[ 78 ][ 356 ],
   alphaCSR[ 78 ][ 357 ],
   alphaCSR[ 78 ][ 358 ],
   alphaCSR[ 78 ][ 359 ],
   alphaCSR[ 78 ][ 360 ],
   alphaCSR[ 78 ][ 361 ],
   alphaCSR[ 78 ][ 362 ],
   alphaCSR[ 78 ][ 363 ],
   alphaCSR[ 78 ][ 364 ],
   alphaCSR[ 78 ][ 365 ],
   alphaCSR[ 78 ][ 366 ],
   alphaCSR[ 78 ][ 367 ],
   alphaCSR[ 78 ][ 368 ],
   alphaCSR[ 78 ][ 369 ],
   alphaCSR[ 78 ][ 370 ],
   alphaCSR[ 78 ][ 371 ],
   alphaCSR[ 78 ][ 372 ],
   alphaCSR[ 78 ][ 373 ],
   alphaCSR[ 78 ][ 374 ],
   alphaCSR[ 78 ][ 375 ],
   alphaCSR[ 78 ][ 376 ],
   alphaCSR[ 78 ][ 377 ],
   alphaCSR[ 78 ][ 378 ],
   alphaCSR[ 78 ][ 379 ],
   alphaCSR[ 78 ][ 380 ],
   alphaCSR[ 78 ][ 381 ],
   alphaCSR[ 78 ][ 382 ],
   alphaCSR[ 78 ][ 383 ],
   alphaCSR[ 79 ][ 0 ],
   alphaCSR[ 79 ][ 1 ],
   alphaCSR[ 79 ][ 2 ],
   alphaCSR[ 79 ][ 3 ],
   alphaCSR[ 79 ][ 4 ],
   alphaCSR[ 79 ][ 5 ],
   alphaCSR[ 79 ][ 6 ],
   alphaCSR[ 79 ][ 7 ],
   alphaCSR[ 79 ][ 8 ],
   alphaCSR[ 79 ][ 9 ],
   alphaCSR[ 79 ][ 10 ],
   alphaCSR[ 79 ][ 11 ],
   alphaCSR[ 79 ][ 12 ],
   alphaCSR[ 79 ][ 13 ],
   alphaCSR[ 79 ][ 14 ],
   alphaCSR[ 79 ][ 15 ],
   alphaCSR[ 79 ][ 16 ],
   alphaCSR[ 79 ][ 17 ],
   alphaCSR[ 79 ][ 18 ],
   alphaCSR[ 79 ][ 19 ],
   alphaCSR[ 79 ][ 20 ],
   alphaCSR[ 79 ][ 21 ],
   alphaCSR[ 79 ][ 22 ],
   alphaCSR[ 79 ][ 23 ],
   alphaCSR[ 79 ][ 24 ],
   alphaCSR[ 79 ][ 25 ],
   alphaCSR[ 79 ][ 26 ],
   alphaCSR[ 79 ][ 27 ],
   alphaCSR[ 79 ][ 28 ],
   alphaCSR[ 79 ][ 29 ],
   alphaCSR[ 79 ][ 30 ],
   alphaCSR[ 79 ][ 31 ],
   alphaCSR[ 79 ][ 32 ],
   alphaCSR[ 79 ][ 33 ],
   alphaCSR[ 79 ][ 34 ],
   alphaCSR[ 79 ][ 35 ],
   alphaCSR[ 79 ][ 36 ],
   alphaCSR[ 79 ][ 37 ],
   alphaCSR[ 79 ][ 38 ],
   alphaCSR[ 79 ][ 39 ],
   alphaCSR[ 79 ][ 40 ],
   alphaCSR[ 79 ][ 41 ],
   alphaCSR[ 79 ][ 42 ],
   alphaCSR[ 79 ][ 43 ],
   alphaCSR[ 79 ][ 44 ],
   alphaCSR[ 79 ][ 45 ],
   alphaCSR[ 79 ][ 46 ],
   alphaCSR[ 79 ][ 47 ],
   alphaCSR[ 79 ][ 48 ],
   alphaCSR[ 79 ][ 49 ],
   alphaCSR[ 79 ][ 50 ],
   alphaCSR[ 79 ][ 51 ],
   alphaCSR[ 79 ][ 52 ],
   alphaCSR[ 79 ][ 53 ],
   alphaCSR[ 79 ][ 54 ],
   alphaCSR[ 79 ][ 55 ],
   alphaCSR[ 79 ][ 56 ],
   alphaCSR[ 79 ][ 57 ],
   alphaCSR[ 79 ][ 58 ],
   alphaCSR[ 79 ][ 59 ],
   alphaCSR[ 79 ][ 60 ],
   alphaCSR[ 79 ][ 61 ],
   alphaCSR[ 79 ][ 62 ],
   alphaCSR[ 79 ][ 63 ],
   alphaCSR[ 79 ][ 64 ],
   alphaCSR[ 79 ][ 65 ],
   alphaCSR[ 79 ][ 66 ],
   alphaCSR[ 79 ][ 67 ],
   alphaCSR[ 79 ][ 68 ],
   alphaCSR[ 79 ][ 69 ],
   alphaCSR[ 79 ][ 70 ],
   alphaCSR[ 79 ][ 71 ],
   alphaCSR[ 79 ][ 72 ],
   alphaCSR[ 79 ][ 73 ],
   alphaCSR[ 79 ][ 74 ],
   alphaCSR[ 79 ][ 75 ],
   alphaCSR[ 79 ][ 76 ],
   alphaCSR[ 79 ][ 77 ],
   alphaCSR[ 79 ][ 78 ],
   alphaCSR[ 79 ][ 79 ],
   alphaCSR[ 79 ][ 80 ],
   alphaCSR[ 79 ][ 81 ],
   alphaCSR[ 79 ][ 82 ],
   alphaCSR[ 79 ][ 83 ],
   alphaCSR[ 79 ][ 84 ],
   alphaCSR[ 79 ][ 85 ],
   alphaCSR[ 79 ][ 86 ],
   alphaCSR[ 79 ][ 87 ],
   alphaCSR[ 79 ][ 88 ],
   alphaCSR[ 79 ][ 89 ],
   alphaCSR[ 79 ][ 90 ],
   alphaCSR[ 79 ][ 91 ],
   alphaCSR[ 79 ][ 92 ],
   alphaCSR[ 79 ][ 93 ],
   alphaCSR[ 79 ][ 94 ],
   alphaCSR[ 79 ][ 95 ],
   alphaCSR[ 79 ][ 96 ],
   alphaCSR[ 79 ][ 97 ],
   alphaCSR[ 79 ][ 98 ],
   alphaCSR[ 79 ][ 99 ],
   alphaCSR[ 79 ][ 100 ],
   alphaCSR[ 79 ][ 101 ],
   alphaCSR[ 79 ][ 102 ],
   alphaCSR[ 79 ][ 103 ],
   alphaCSR[ 79 ][ 104 ],
   alphaCSR[ 79 ][ 105 ],
   alphaCSR[ 79 ][ 106 ],
   alphaCSR[ 79 ][ 107 ],
   alphaCSR[ 79 ][ 108 ],
   alphaCSR[ 79 ][ 109 ],
   alphaCSR[ 79 ][ 110 ],
   alphaCSR[ 79 ][ 111 ],
   alphaCSR[ 79 ][ 112 ],
   alphaCSR[ 79 ][ 113 ],
   alphaCSR[ 79 ][ 114 ],
   alphaCSR[ 79 ][ 115 ],
   alphaCSR[ 79 ][ 116 ],
   alphaCSR[ 79 ][ 117 ],
   alphaCSR[ 79 ][ 118 ],
   alphaCSR[ 79 ][ 119 ],
   alphaCSR[ 79 ][ 120 ],
   alphaCSR[ 79 ][ 121 ],
   alphaCSR[ 79 ][ 122 ],
   alphaCSR[ 79 ][ 123 ],
   alphaCSR[ 79 ][ 124 ],
   alphaCSR[ 79 ][ 125 ],
   alphaCSR[ 79 ][ 126 ],
   alphaCSR[ 79 ][ 127 ],
   alphaCSR[ 79 ][ 128 ],
   alphaCSR[ 79 ][ 129 ],
   alphaCSR[ 79 ][ 130 ],
   alphaCSR[ 79 ][ 131 ],
   alphaCSR[ 79 ][ 132 ],
   alphaCSR[ 79 ][ 133 ],
   alphaCSR[ 79 ][ 134 ],
   alphaCSR[ 79 ][ 135 ],
   alphaCSR[ 79 ][ 136 ],
   alphaCSR[ 79 ][ 137 ],
   alphaCSR[ 79 ][ 138 ],
   alphaCSR[ 79 ][ 139 ],
   alphaCSR[ 79 ][ 140 ],
   alphaCSR[ 79 ][ 141 ],
   alphaCSR[ 79 ][ 142 ],
   alphaCSR[ 79 ][ 143 ],
   alphaCSR[ 79 ][ 144 ],
   alphaCSR[ 79 ][ 145 ],
   alphaCSR[ 79 ][ 146 ],
   alphaCSR[ 79 ][ 147 ],
   alphaCSR[ 79 ][ 148 ],
   alphaCSR[ 79 ][ 149 ],
   alphaCSR[ 79 ][ 150 ],
   alphaCSR[ 79 ][ 151 ],
   alphaCSR[ 79 ][ 152 ],
   alphaCSR[ 79 ][ 153 ],
   alphaCSR[ 79 ][ 154 ],
   alphaCSR[ 79 ][ 155 ],
   alphaCSR[ 79 ][ 156 ],
   alphaCSR[ 79 ][ 157 ],
   alphaCSR[ 79 ][ 158 ],
   alphaCSR[ 79 ][ 159 ],
   alphaCSR[ 79 ][ 160 ],
   alphaCSR[ 79 ][ 161 ],
   alphaCSR[ 79 ][ 162 ],
   alphaCSR[ 79 ][ 163 ],
   alphaCSR[ 79 ][ 164 ],
   alphaCSR[ 79 ][ 165 ],
   alphaCSR[ 79 ][ 166 ],
   alphaCSR[ 79 ][ 167 ],
   alphaCSR[ 79 ][ 168 ],
   alphaCSR[ 79 ][ 169 ],
   alphaCSR[ 79 ][ 170 ],
   alphaCSR[ 79 ][ 171 ],
   alphaCSR[ 79 ][ 172 ],
   alphaCSR[ 79 ][ 173 ],
   alphaCSR[ 79 ][ 174 ],
   alphaCSR[ 79 ][ 175 ],
   alphaCSR[ 79 ][ 176 ],
   alphaCSR[ 79 ][ 177 ],
   alphaCSR[ 79 ][ 178 ],
   alphaCSR[ 79 ][ 179 ],
   alphaCSR[ 79 ][ 180 ],
   alphaCSR[ 79 ][ 181 ],
   alphaCSR[ 79 ][ 182 ],
   alphaCSR[ 79 ][ 183 ],
   alphaCSR[ 79 ][ 184 ],
   alphaCSR[ 79 ][ 185 ],
   alphaCSR[ 79 ][ 186 ],
   alphaCSR[ 79 ][ 187 ],
   alphaCSR[ 79 ][ 188 ],
   alphaCSR[ 79 ][ 189 ],
   alphaCSR[ 79 ][ 190 ],
   alphaCSR[ 79 ][ 191 ],
   alphaCSR[ 79 ][ 192 ],
   alphaCSR[ 79 ][ 193 ],
   alphaCSR[ 79 ][ 194 ],
   alphaCSR[ 79 ][ 195 ],
   alphaCSR[ 79 ][ 196 ],
   alphaCSR[ 79 ][ 197 ],
   alphaCSR[ 79 ][ 198 ],
   alphaCSR[ 79 ][ 199 ],
   alphaCSR[ 79 ][ 200 ],
   alphaCSR[ 79 ][ 201 ],
   alphaCSR[ 79 ][ 202 ],
   alphaCSR[ 79 ][ 203 ],
   alphaCSR[ 79 ][ 204 ],
   alphaCSR[ 79 ][ 205 ],
   alphaCSR[ 79 ][ 206 ],
   alphaCSR[ 79 ][ 207 ],
   alphaCSR[ 79 ][ 208 ],
   alphaCSR[ 79 ][ 209 ],
   alphaCSR[ 79 ][ 210 ],
   alphaCSR[ 79 ][ 211 ],
   alphaCSR[ 79 ][ 212 ],
   alphaCSR[ 79 ][ 213 ],
   alphaCSR[ 79 ][ 214 ],
   alphaCSR[ 79 ][ 215 ],
   alphaCSR[ 79 ][ 216 ],
   alphaCSR[ 79 ][ 217 ],
   alphaCSR[ 79 ][ 218 ],
   alphaCSR[ 79 ][ 219 ],
   alphaCSR[ 79 ][ 220 ],
   alphaCSR[ 79 ][ 221 ],
   alphaCSR[ 79 ][ 222 ],
   alphaCSR[ 79 ][ 223 ],
   alphaCSR[ 79 ][ 224 ],
   alphaCSR[ 79 ][ 225 ],
   alphaCSR[ 79 ][ 226 ],
   alphaCSR[ 79 ][ 227 ],
   alphaCSR[ 79 ][ 228 ],
   alphaCSR[ 79 ][ 229 ],
   alphaCSR[ 79 ][ 230 ],
   alphaCSR[ 79 ][ 231 ],
   alphaCSR[ 79 ][ 232 ],
   alphaCSR[ 79 ][ 233 ],
   alphaCSR[ 79 ][ 234 ],
   alphaCSR[ 79 ][ 235 ],
   alphaCSR[ 79 ][ 236 ],
   alphaCSR[ 79 ][ 237 ],
   alphaCSR[ 79 ][ 238 ],
   alphaCSR[ 79 ][ 239 ],
   alphaCSR[ 79 ][ 240 ],
   alphaCSR[ 79 ][ 241 ],
   alphaCSR[ 79 ][ 242 ],
   alphaCSR[ 79 ][ 243 ],
   alphaCSR[ 79 ][ 244 ],
   alphaCSR[ 79 ][ 245 ],
   alphaCSR[ 79 ][ 246 ],
   alphaCSR[ 79 ][ 247 ],
   alphaCSR[ 79 ][ 248 ],
   alphaCSR[ 79 ][ 249 ],
   alphaCSR[ 79 ][ 250 ],
   alphaCSR[ 79 ][ 251 ],
   alphaCSR[ 79 ][ 252 ],
   alphaCSR[ 79 ][ 253 ],
   alphaCSR[ 79 ][ 254 ],
   alphaCSR[ 79 ][ 255 ],
   alphaCSR[ 79 ][ 256 ],
   alphaCSR[ 79 ][ 257 ],
   alphaCSR[ 79 ][ 258 ],
   alphaCSR[ 79 ][ 259 ],
   alphaCSR[ 79 ][ 260 ],
   alphaCSR[ 79 ][ 261 ],
   alphaCSR[ 79 ][ 262 ],
   alphaCSR[ 79 ][ 263 ],
   alphaCSR[ 79 ][ 264 ],
   alphaCSR[ 79 ][ 265 ],
   alphaCSR[ 79 ][ 266 ],
   alphaCSR[ 79 ][ 267 ],
   alphaCSR[ 79 ][ 268 ],
   alphaCSR[ 79 ][ 269 ],
   alphaCSR[ 79 ][ 270 ],
   alphaCSR[ 79 ][ 271 ],
   alphaCSR[ 79 ][ 272 ],
   alphaCSR[ 79 ][ 273 ],
   alphaCSR[ 79 ][ 274 ],
   alphaCSR[ 79 ][ 275 ],
   alphaCSR[ 79 ][ 276 ],
   alphaCSR[ 79 ][ 277 ],
   alphaCSR[ 79 ][ 278 ],
   alphaCSR[ 79 ][ 279 ],
   alphaCSR[ 79 ][ 280 ],
   alphaCSR[ 79 ][ 281 ],
   alphaCSR[ 79 ][ 282 ],
   alphaCSR[ 79 ][ 283 ],
   alphaCSR[ 79 ][ 284 ],
   alphaCSR[ 79 ][ 285 ],
   alphaCSR[ 79 ][ 286 ],
   alphaCSR[ 79 ][ 287 ],
   alphaCSR[ 79 ][ 288 ],
   alphaCSR[ 79 ][ 289 ],
   alphaCSR[ 79 ][ 290 ],
   alphaCSR[ 79 ][ 291 ],
   alphaCSR[ 79 ][ 292 ],
   alphaCSR[ 79 ][ 293 ],
   alphaCSR[ 79 ][ 294 ],
   alphaCSR[ 79 ][ 295 ],
   alphaCSR[ 79 ][ 296 ],
   alphaCSR[ 79 ][ 297 ],
   alphaCSR[ 79 ][ 298 ],
   alphaCSR[ 79 ][ 299 ],
   alphaCSR[ 79 ][ 300 ],
   alphaCSR[ 79 ][ 301 ],
   alphaCSR[ 79 ][ 302 ],
   alphaCSR[ 79 ][ 303 ],
   alphaCSR[ 79 ][ 304 ],
   alphaCSR[ 79 ][ 305 ],
   alphaCSR[ 79 ][ 306 ],
   alphaCSR[ 79 ][ 307 ],
   alphaCSR[ 79 ][ 308 ],
   alphaCSR[ 79 ][ 309 ],
   alphaCSR[ 79 ][ 310 ],
   alphaCSR[ 79 ][ 311 ],
   alphaCSR[ 79 ][ 312 ],
   alphaCSR[ 79 ][ 313 ],
   alphaCSR[ 79 ][ 314 ],
   alphaCSR[ 79 ][ 315 ],
   alphaCSR[ 79 ][ 316 ],
   alphaCSR[ 79 ][ 317 ],
   alphaCSR[ 79 ][ 318 ],
   alphaCSR[ 79 ][ 319 ],
   alphaCSR[ 79 ][ 320 ],
   alphaCSR[ 79 ][ 321 ],
   alphaCSR[ 79 ][ 322 ],
   alphaCSR[ 79 ][ 323 ],
   alphaCSR[ 79 ][ 324 ],
   alphaCSR[ 79 ][ 325 ],
   alphaCSR[ 79 ][ 326 ],
   alphaCSR[ 79 ][ 327 ],
   alphaCSR[ 79 ][ 328 ],
   alphaCSR[ 79 ][ 329 ],
   alphaCSR[ 79 ][ 330 ],
   alphaCSR[ 79 ][ 331 ],
   alphaCSR[ 79 ][ 332 ],
   alphaCSR[ 79 ][ 333 ],
   alphaCSR[ 79 ][ 334 ],
   alphaCSR[ 79 ][ 335 ],
   alphaCSR[ 79 ][ 336 ],
   alphaCSR[ 79 ][ 337 ],
   alphaCSR[ 79 ][ 338 ],
   alphaCSR[ 79 ][ 339 ],
   alphaCSR[ 79 ][ 340 ],
   alphaCSR[ 79 ][ 341 ],
   alphaCSR[ 79 ][ 342 ],
   alphaCSR[ 79 ][ 343 ],
   alphaCSR[ 79 ][ 344 ],
   alphaCSR[ 79 ][ 345 ],
   alphaCSR[ 79 ][ 346 ],
   alphaCSR[ 79 ][ 347 ],
   alphaCSR[ 79 ][ 348 ],
   alphaCSR[ 79 ][ 349 ],
   alphaCSR[ 79 ][ 350 ],
   alphaCSR[ 79 ][ 351 ],
   alphaCSR[ 79 ][ 352 ],
   alphaCSR[ 79 ][ 353 ],
   alphaCSR[ 79 ][ 354 ],
   alphaCSR[ 79 ][ 355 ],
   alphaCSR[ 79 ][ 356 ],
   alphaCSR[ 79 ][ 357 ],
   alphaCSR[ 79 ][ 358 ],
   alphaCSR[ 79 ][ 359 ],
   alphaCSR[ 79 ][ 360 ],
   alphaCSR[ 79 ][ 361 ],
   alphaCSR[ 79 ][ 362 ],
   alphaCSR[ 79 ][ 363 ],
   alphaCSR[ 79 ][ 364 ],
   alphaCSR[ 79 ][ 365 ],
   alphaCSR[ 79 ][ 366 ],
   alphaCSR[ 79 ][ 367 ],
   alphaCSR[ 79 ][ 368 ],
   alphaCSR[ 79 ][ 369 ],
   alphaCSR[ 79 ][ 370 ],
   alphaCSR[ 79 ][ 371 ],
   alphaCSR[ 79 ][ 372 ],
   alphaCSR[ 79 ][ 373 ],
   alphaCSR[ 79 ][ 374 ],
   alphaCSR[ 79 ][ 375 ],
   alphaCSR[ 79 ][ 376 ],
   alphaCSR[ 79 ][ 377 ],
   alphaCSR[ 79 ][ 378 ],
   alphaCSR[ 79 ][ 379 ],
   alphaCSR[ 79 ][ 380 ],
   alphaCSR[ 79 ][ 381 ],
   alphaCSR[ 79 ][ 382 ],
   alphaCSR[ 79 ][ 383 ],
   alphaCSR[ 80 ][ 0 ],
   alphaCSR[ 80 ][ 1 ],
   alphaCSR[ 80 ][ 2 ],
   alphaCSR[ 80 ][ 3 ],
   alphaCSR[ 80 ][ 4 ],
   alphaCSR[ 80 ][ 5 ],
   alphaCSR[ 80 ][ 6 ],
   alphaCSR[ 80 ][ 7 ],
   alphaCSR[ 80 ][ 8 ],
   alphaCSR[ 80 ][ 9 ],
   alphaCSR[ 80 ][ 10 ],
   alphaCSR[ 80 ][ 11 ],
   alphaCSR[ 80 ][ 12 ],
   alphaCSR[ 80 ][ 13 ],
   alphaCSR[ 80 ][ 14 ],
   alphaCSR[ 80 ][ 15 ],
   alphaCSR[ 80 ][ 16 ],
   alphaCSR[ 80 ][ 17 ],
   alphaCSR[ 80 ][ 18 ],
   alphaCSR[ 80 ][ 19 ],
   alphaCSR[ 80 ][ 20 ],
   alphaCSR[ 80 ][ 21 ],
   alphaCSR[ 80 ][ 22 ],
   alphaCSR[ 80 ][ 23 ],
   alphaCSR[ 80 ][ 24 ],
   alphaCSR[ 80 ][ 25 ],
   alphaCSR[ 80 ][ 26 ],
   alphaCSR[ 80 ][ 27 ],
   alphaCSR[ 80 ][ 28 ],
   alphaCSR[ 80 ][ 29 ],
   alphaCSR[ 80 ][ 30 ],
   alphaCSR[ 80 ][ 31 ],
   alphaCSR[ 80 ][ 32 ],
   alphaCSR[ 80 ][ 33 ],
   alphaCSR[ 80 ][ 34 ],
   alphaCSR[ 80 ][ 35 ],
   alphaCSR[ 80 ][ 36 ],
   alphaCSR[ 80 ][ 37 ],
   alphaCSR[ 80 ][ 38 ],
   alphaCSR[ 80 ][ 39 ],
   alphaCSR[ 80 ][ 40 ],
   alphaCSR[ 80 ][ 41 ],
   alphaCSR[ 80 ][ 42 ],
   alphaCSR[ 80 ][ 43 ],
   alphaCSR[ 80 ][ 44 ],
   alphaCSR[ 80 ][ 45 ],
   alphaCSR[ 80 ][ 46 ],
   alphaCSR[ 80 ][ 47 ],
   alphaCSR[ 80 ][ 48 ],
   alphaCSR[ 80 ][ 49 ],
   alphaCSR[ 80 ][ 50 ],
   alphaCSR[ 80 ][ 51 ],
   alphaCSR[ 80 ][ 52 ],
   alphaCSR[ 80 ][ 53 ],
   alphaCSR[ 80 ][ 54 ],
   alphaCSR[ 80 ][ 55 ],
   alphaCSR[ 80 ][ 56 ],
   alphaCSR[ 80 ][ 57 ],
   alphaCSR[ 80 ][ 58 ],
   alphaCSR[ 80 ][ 59 ],
   alphaCSR[ 80 ][ 60 ],
   alphaCSR[ 80 ][ 61 ],
   alphaCSR[ 80 ][ 62 ],
   alphaCSR[ 80 ][ 63 ],
   alphaCSR[ 80 ][ 64 ],
   alphaCSR[ 80 ][ 65 ],
   alphaCSR[ 80 ][ 66 ],
   alphaCSR[ 80 ][ 67 ],
   alphaCSR[ 80 ][ 68 ],
   alphaCSR[ 80 ][ 69 ],
   alphaCSR[ 80 ][ 70 ],
   alphaCSR[ 80 ][ 71 ],
   alphaCSR[ 80 ][ 72 ],
   alphaCSR[ 80 ][ 73 ],
   alphaCSR[ 80 ][ 74 ],
   alphaCSR[ 80 ][ 75 ],
   alphaCSR[ 80 ][ 76 ],
   alphaCSR[ 80 ][ 77 ],
   alphaCSR[ 80 ][ 78 ],
   alphaCSR[ 80 ][ 79 ],
   alphaCSR[ 80 ][ 80 ],
   alphaCSR[ 80 ][ 81 ],
   alphaCSR[ 80 ][ 82 ],
   alphaCSR[ 80 ][ 83 ],
   alphaCSR[ 80 ][ 84 ],
   alphaCSR[ 80 ][ 85 ],
   alphaCSR[ 80 ][ 86 ],
   alphaCSR[ 80 ][ 87 ],
   alphaCSR[ 80 ][ 88 ],
   alphaCSR[ 80 ][ 89 ],
   alphaCSR[ 80 ][ 90 ],
   alphaCSR[ 80 ][ 91 ],
   alphaCSR[ 80 ][ 92 ],
   alphaCSR[ 80 ][ 93 ],
   alphaCSR[ 80 ][ 94 ],
   alphaCSR[ 80 ][ 95 ],
   alphaCSR[ 80 ][ 96 ],
   alphaCSR[ 80 ][ 97 ],
   alphaCSR[ 80 ][ 98 ],
   alphaCSR[ 80 ][ 99 ],
   alphaCSR[ 80 ][ 100 ],
   alphaCSR[ 80 ][ 101 ],
   alphaCSR[ 80 ][ 102 ],
   alphaCSR[ 80 ][ 103 ],
   alphaCSR[ 80 ][ 104 ],
   alphaCSR[ 80 ][ 105 ],
   alphaCSR[ 80 ][ 106 ],
   alphaCSR[ 80 ][ 107 ],
   alphaCSR[ 80 ][ 108 ],
   alphaCSR[ 80 ][ 109 ],
   alphaCSR[ 80 ][ 110 ],
   alphaCSR[ 80 ][ 111 ],
   alphaCSR[ 80 ][ 112 ],
   alphaCSR[ 80 ][ 113 ],
   alphaCSR[ 80 ][ 114 ],
   alphaCSR[ 80 ][ 115 ],
   alphaCSR[ 80 ][ 116 ],
   alphaCSR[ 80 ][ 117 ],
   alphaCSR[ 80 ][ 118 ],
   alphaCSR[ 80 ][ 119 ],
   alphaCSR[ 80 ][ 120 ],
   alphaCSR[ 80 ][ 121 ],
   alphaCSR[ 80 ][ 122 ],
   alphaCSR[ 80 ][ 123 ],
   alphaCSR[ 80 ][ 124 ],
   alphaCSR[ 80 ][ 125 ],
   alphaCSR[ 80 ][ 126 ],
   alphaCSR[ 80 ][ 127 ],
   alphaCSR[ 80 ][ 128 ],
   alphaCSR[ 80 ][ 129 ],
   alphaCSR[ 80 ][ 130 ],
   alphaCSR[ 80 ][ 131 ],
   alphaCSR[ 80 ][ 132 ],
   alphaCSR[ 80 ][ 133 ],
   alphaCSR[ 80 ][ 134 ],
   alphaCSR[ 80 ][ 135 ],
   alphaCSR[ 80 ][ 136 ],
   alphaCSR[ 80 ][ 137 ],
   alphaCSR[ 80 ][ 138 ],
   alphaCSR[ 80 ][ 139 ],
   alphaCSR[ 80 ][ 140 ],
   alphaCSR[ 80 ][ 141 ],
   alphaCSR[ 80 ][ 142 ],
   alphaCSR[ 80 ][ 143 ],
   alphaCSR[ 80 ][ 144 ],
   alphaCSR[ 80 ][ 145 ],
   alphaCSR[ 80 ][ 146 ],
   alphaCSR[ 80 ][ 147 ],
   alphaCSR[ 80 ][ 148 ],
   alphaCSR[ 80 ][ 149 ],
   alphaCSR[ 80 ][ 150 ],
   alphaCSR[ 80 ][ 151 ],
   alphaCSR[ 80 ][ 152 ],
   alphaCSR[ 80 ][ 153 ],
   alphaCSR[ 80 ][ 154 ],
   alphaCSR[ 80 ][ 155 ],
   alphaCSR[ 80 ][ 156 ],
   alphaCSR[ 80 ][ 157 ],
   alphaCSR[ 80 ][ 158 ],
   alphaCSR[ 80 ][ 159 ],
   alphaCSR[ 80 ][ 160 ],
   alphaCSR[ 80 ][ 161 ],
   alphaCSR[ 80 ][ 162 ],
   alphaCSR[ 80 ][ 163 ],
   alphaCSR[ 80 ][ 164 ],
   alphaCSR[ 80 ][ 165 ],
   alphaCSR[ 80 ][ 166 ],
   alphaCSR[ 80 ][ 167 ],
   alphaCSR[ 80 ][ 168 ],
   alphaCSR[ 80 ][ 169 ],
   alphaCSR[ 80 ][ 170 ],
   alphaCSR[ 80 ][ 171 ],
   alphaCSR[ 80 ][ 172 ],
   alphaCSR[ 80 ][ 173 ],
   alphaCSR[ 80 ][ 174 ],
   alphaCSR[ 80 ][ 175 ],
   alphaCSR[ 80 ][ 176 ],
   alphaCSR[ 80 ][ 177 ],
   alphaCSR[ 80 ][ 178 ],
   alphaCSR[ 80 ][ 179 ],
   alphaCSR[ 80 ][ 180 ],
   alphaCSR[ 80 ][ 181 ],
   alphaCSR[ 80 ][ 182 ],
   alphaCSR[ 80 ][ 183 ],
   alphaCSR[ 80 ][ 184 ],
   alphaCSR[ 80 ][ 185 ],
   alphaCSR[ 80 ][ 186 ],
   alphaCSR[ 80 ][ 187 ],
   alphaCSR[ 80 ][ 188 ],
   alphaCSR[ 80 ][ 189 ],
   alphaCSR[ 80 ][ 190 ],
   alphaCSR[ 80 ][ 191 ],
   alphaCSR[ 80 ][ 192 ],
   alphaCSR[ 80 ][ 193 ],
   alphaCSR[ 80 ][ 194 ],
   alphaCSR[ 80 ][ 195 ],
   alphaCSR[ 80 ][ 196 ],
   alphaCSR[ 80 ][ 197 ],
   alphaCSR[ 80 ][ 198 ],
   alphaCSR[ 80 ][ 199 ],
   alphaCSR[ 80 ][ 200 ],
   alphaCSR[ 80 ][ 201 ],
   alphaCSR[ 80 ][ 202 ],
   alphaCSR[ 80 ][ 203 ],
   alphaCSR[ 80 ][ 204 ],
   alphaCSR[ 80 ][ 205 ],
   alphaCSR[ 80 ][ 206 ],
   alphaCSR[ 80 ][ 207 ],
   alphaCSR[ 80 ][ 208 ],
   alphaCSR[ 80 ][ 209 ],
   alphaCSR[ 80 ][ 210 ],
   alphaCSR[ 80 ][ 211 ],
   alphaCSR[ 80 ][ 212 ],
   alphaCSR[ 80 ][ 213 ],
   alphaCSR[ 80 ][ 214 ],
   alphaCSR[ 80 ][ 215 ],
   alphaCSR[ 80 ][ 216 ],
   alphaCSR[ 80 ][ 217 ],
   alphaCSR[ 80 ][ 218 ],
   alphaCSR[ 80 ][ 219 ],
   alphaCSR[ 80 ][ 220 ],
   alphaCSR[ 80 ][ 221 ],
   alphaCSR[ 80 ][ 222 ],
   alphaCSR[ 80 ][ 223 ],
   alphaCSR[ 80 ][ 224 ],
   alphaCSR[ 80 ][ 225 ],
   alphaCSR[ 80 ][ 226 ],
   alphaCSR[ 80 ][ 227 ],
   alphaCSR[ 80 ][ 228 ],
   alphaCSR[ 80 ][ 229 ],
   alphaCSR[ 80 ][ 230 ],
   alphaCSR[ 80 ][ 231 ],
   alphaCSR[ 80 ][ 232 ],
   alphaCSR[ 80 ][ 233 ],
   alphaCSR[ 80 ][ 234 ],
   alphaCSR[ 80 ][ 235 ],
   alphaCSR[ 80 ][ 236 ],
   alphaCSR[ 80 ][ 237 ],
   alphaCSR[ 80 ][ 238 ],
   alphaCSR[ 80 ][ 239 ],
   alphaCSR[ 80 ][ 240 ],
   alphaCSR[ 80 ][ 241 ],
   alphaCSR[ 80 ][ 242 ],
   alphaCSR[ 80 ][ 243 ],
   alphaCSR[ 80 ][ 244 ],
   alphaCSR[ 80 ][ 245 ],
   alphaCSR[ 80 ][ 246 ],
   alphaCSR[ 80 ][ 247 ],
   alphaCSR[ 80 ][ 248 ],
   alphaCSR[ 80 ][ 249 ],
   alphaCSR[ 80 ][ 250 ],
   alphaCSR[ 80 ][ 251 ],
   alphaCSR[ 80 ][ 252 ],
   alphaCSR[ 80 ][ 253 ],
   alphaCSR[ 80 ][ 254 ],
   alphaCSR[ 80 ][ 255 ],
   alphaCSR[ 80 ][ 256 ],
   alphaCSR[ 80 ][ 257 ],
   alphaCSR[ 80 ][ 258 ],
   alphaCSR[ 80 ][ 259 ],
   alphaCSR[ 80 ][ 260 ],
   alphaCSR[ 80 ][ 261 ],
   alphaCSR[ 80 ][ 262 ],
   alphaCSR[ 80 ][ 263 ],
   alphaCSR[ 80 ][ 264 ],
   alphaCSR[ 80 ][ 265 ],
   alphaCSR[ 80 ][ 266 ],
   alphaCSR[ 80 ][ 267 ],
   alphaCSR[ 80 ][ 268 ],
   alphaCSR[ 80 ][ 269 ],
   alphaCSR[ 80 ][ 270 ],
   alphaCSR[ 80 ][ 271 ],
   alphaCSR[ 80 ][ 272 ],
   alphaCSR[ 80 ][ 273 ],
   alphaCSR[ 80 ][ 274 ],
   alphaCSR[ 80 ][ 275 ],
   alphaCSR[ 80 ][ 276 ],
   alphaCSR[ 80 ][ 277 ],
   alphaCSR[ 80 ][ 278 ],
   alphaCSR[ 80 ][ 279 ],
   alphaCSR[ 80 ][ 280 ],
   alphaCSR[ 80 ][ 281 ],
   alphaCSR[ 80 ][ 282 ],
   alphaCSR[ 80 ][ 283 ],
   alphaCSR[ 80 ][ 284 ],
   alphaCSR[ 80 ][ 285 ],
   alphaCSR[ 80 ][ 286 ],
   alphaCSR[ 80 ][ 287 ],
   alphaCSR[ 80 ][ 288 ],
   alphaCSR[ 80 ][ 289 ],
   alphaCSR[ 80 ][ 290 ],
   alphaCSR[ 80 ][ 291 ],
   alphaCSR[ 80 ][ 292 ],
   alphaCSR[ 80 ][ 293 ],
   alphaCSR[ 80 ][ 294 ],
   alphaCSR[ 80 ][ 295 ],
   alphaCSR[ 80 ][ 296 ],
   alphaCSR[ 80 ][ 297 ],
   alphaCSR[ 80 ][ 298 ],
   alphaCSR[ 80 ][ 299 ],
   alphaCSR[ 80 ][ 300 ],
   alphaCSR[ 80 ][ 301 ],
   alphaCSR[ 80 ][ 302 ],
   alphaCSR[ 80 ][ 303 ],
   alphaCSR[ 80 ][ 304 ],
   alphaCSR[ 80 ][ 305 ],
   alphaCSR[ 80 ][ 306 ],
   alphaCSR[ 80 ][ 307 ],
   alphaCSR[ 80 ][ 308 ],
   alphaCSR[ 80 ][ 309 ],
   alphaCSR[ 80 ][ 310 ],
   alphaCSR[ 80 ][ 311 ],
   alphaCSR[ 80 ][ 312 ],
   alphaCSR[ 80 ][ 313 ],
   alphaCSR[ 80 ][ 314 ],
   alphaCSR[ 80 ][ 315 ],
   alphaCSR[ 80 ][ 316 ],
   alphaCSR[ 80 ][ 317 ],
   alphaCSR[ 80 ][ 318 ],
   alphaCSR[ 80 ][ 319 ],
   alphaCSR[ 80 ][ 320 ],
   alphaCSR[ 80 ][ 321 ],
   alphaCSR[ 80 ][ 322 ],
   alphaCSR[ 80 ][ 323 ],
   alphaCSR[ 80 ][ 324 ],
   alphaCSR[ 80 ][ 325 ],
   alphaCSR[ 80 ][ 326 ],
   alphaCSR[ 80 ][ 327 ],
   alphaCSR[ 80 ][ 328 ],
   alphaCSR[ 80 ][ 329 ],
   alphaCSR[ 80 ][ 330 ],
   alphaCSR[ 80 ][ 331 ],
   alphaCSR[ 80 ][ 332 ],
   alphaCSR[ 80 ][ 333 ],
   alphaCSR[ 80 ][ 334 ],
   alphaCSR[ 80 ][ 335 ],
   alphaCSR[ 80 ][ 336 ],
   alphaCSR[ 80 ][ 337 ],
   alphaCSR[ 80 ][ 338 ],
   alphaCSR[ 80 ][ 339 ],
   alphaCSR[ 80 ][ 340 ],
   alphaCSR[ 80 ][ 341 ],
   alphaCSR[ 80 ][ 342 ],
   alphaCSR[ 80 ][ 343 ],
   alphaCSR[ 80 ][ 344 ],
   alphaCSR[ 80 ][ 345 ],
   alphaCSR[ 80 ][ 346 ],
   alphaCSR[ 80 ][ 347 ],
   alphaCSR[ 80 ][ 348 ],
   alphaCSR[ 80 ][ 349 ],
   alphaCSR[ 80 ][ 350 ],
   alphaCSR[ 80 ][ 351 ],
   alphaCSR[ 80 ][ 352 ],
   alphaCSR[ 80 ][ 353 ],
   alphaCSR[ 80 ][ 354 ],
   alphaCSR[ 80 ][ 355 ],
   alphaCSR[ 80 ][ 356 ],
   alphaCSR[ 80 ][ 357 ],
   alphaCSR[ 80 ][ 358 ],
   alphaCSR[ 80 ][ 359 ],
   alphaCSR[ 80 ][ 360 ],
   alphaCSR[ 80 ][ 361 ],
   alphaCSR[ 80 ][ 362 ],
   alphaCSR[ 80 ][ 363 ],
   alphaCSR[ 80 ][ 364 ],
   alphaCSR[ 80 ][ 365 ],
   alphaCSR[ 80 ][ 366 ],
   alphaCSR[ 80 ][ 367 ],
   alphaCSR[ 80 ][ 368 ],
   alphaCSR[ 80 ][ 369 ],
   alphaCSR[ 80 ][ 370 ],
   alphaCSR[ 80 ][ 371 ],
   alphaCSR[ 80 ][ 372 ],
   alphaCSR[ 80 ][ 373 ],
   alphaCSR[ 80 ][ 374 ],
   alphaCSR[ 80 ][ 375 ],
   alphaCSR[ 80 ][ 376 ],
   alphaCSR[ 80 ][ 377 ],
   alphaCSR[ 80 ][ 378 ],
   alphaCSR[ 80 ][ 379 ],
   alphaCSR[ 80 ][ 380 ],
   alphaCSR[ 80 ][ 381 ],
   alphaCSR[ 80 ][ 382 ],
   alphaCSR[ 80 ][ 383 ],
   alphaCSR[ 81 ][ 0 ],
   alphaCSR[ 81 ][ 1 ],
   alphaCSR[ 81 ][ 2 ],
   alphaCSR[ 81 ][ 3 ],
   alphaCSR[ 81 ][ 4 ],
   alphaCSR[ 81 ][ 5 ],
   alphaCSR[ 81 ][ 6 ],
   alphaCSR[ 81 ][ 7 ],
   alphaCSR[ 81 ][ 8 ],
   alphaCSR[ 81 ][ 9 ],
   alphaCSR[ 81 ][ 10 ],
   alphaCSR[ 81 ][ 11 ],
   alphaCSR[ 81 ][ 12 ],
   alphaCSR[ 81 ][ 13 ],
   alphaCSR[ 81 ][ 14 ],
   alphaCSR[ 81 ][ 15 ],
   alphaCSR[ 81 ][ 16 ],
   alphaCSR[ 81 ][ 17 ],
   alphaCSR[ 81 ][ 18 ],
   alphaCSR[ 81 ][ 19 ],
   alphaCSR[ 81 ][ 20 ],
   alphaCSR[ 81 ][ 21 ],
   alphaCSR[ 81 ][ 22 ],
   alphaCSR[ 81 ][ 23 ],
   alphaCSR[ 81 ][ 24 ],
   alphaCSR[ 81 ][ 25 ],
   alphaCSR[ 81 ][ 26 ],
   alphaCSR[ 81 ][ 27 ],
   alphaCSR[ 81 ][ 28 ],
   alphaCSR[ 81 ][ 29 ],
   alphaCSR[ 81 ][ 30 ],
   alphaCSR[ 81 ][ 31 ],
   alphaCSR[ 81 ][ 32 ],
   alphaCSR[ 81 ][ 33 ],
   alphaCSR[ 81 ][ 34 ],
   alphaCSR[ 81 ][ 35 ],
   alphaCSR[ 81 ][ 36 ],
   alphaCSR[ 81 ][ 37 ],
   alphaCSR[ 81 ][ 38 ],
   alphaCSR[ 81 ][ 39 ],
   alphaCSR[ 81 ][ 40 ],
   alphaCSR[ 81 ][ 41 ],
   alphaCSR[ 81 ][ 42 ],
   alphaCSR[ 81 ][ 43 ],
   alphaCSR[ 81 ][ 44 ],
   alphaCSR[ 81 ][ 45 ],
   alphaCSR[ 81 ][ 46 ],
   alphaCSR[ 81 ][ 47 ],
   alphaCSR[ 81 ][ 48 ],
   alphaCSR[ 81 ][ 49 ],
   alphaCSR[ 81 ][ 50 ],
   alphaCSR[ 81 ][ 51 ],
   alphaCSR[ 81 ][ 52 ],
   alphaCSR[ 81 ][ 53 ],
   alphaCSR[ 81 ][ 54 ],
   alphaCSR[ 81 ][ 55 ],
   alphaCSR[ 81 ][ 56 ],
   alphaCSR[ 81 ][ 57 ],
   alphaCSR[ 81 ][ 58 ],
   alphaCSR[ 81 ][ 59 ],
   alphaCSR[ 81 ][ 60 ],
   alphaCSR[ 81 ][ 61 ],
   alphaCSR[ 81 ][ 62 ],
   alphaCSR[ 81 ][ 63 ],
   alphaCSR[ 81 ][ 64 ],
   alphaCSR[ 81 ][ 65 ],
   alphaCSR[ 81 ][ 66 ],
   alphaCSR[ 81 ][ 67 ],
   alphaCSR[ 81 ][ 68 ],
   alphaCSR[ 81 ][ 69 ],
   alphaCSR[ 81 ][ 70 ],
   alphaCSR[ 81 ][ 71 ],
   alphaCSR[ 81 ][ 72 ],
   alphaCSR[ 81 ][ 73 ],
   alphaCSR[ 81 ][ 74 ],
   alphaCSR[ 81 ][ 75 ],
   alphaCSR[ 81 ][ 76 ],
   alphaCSR[ 81 ][ 77 ],
   alphaCSR[ 81 ][ 78 ],
   alphaCSR[ 81 ][ 79 ],
   alphaCSR[ 81 ][ 80 ],
   alphaCSR[ 81 ][ 81 ],
   alphaCSR[ 81 ][ 82 ],
   alphaCSR[ 81 ][ 83 ],
   alphaCSR[ 81 ][ 84 ],
   alphaCSR[ 81 ][ 85 ],
   alphaCSR[ 81 ][ 86 ],
   alphaCSR[ 81 ][ 87 ],
   alphaCSR[ 81 ][ 88 ],
   alphaCSR[ 81 ][ 89 ],
   alphaCSR[ 81 ][ 90 ],
   alphaCSR[ 81 ][ 91 ],
   alphaCSR[ 81 ][ 92 ],
   alphaCSR[ 81 ][ 93 ],
   alphaCSR[ 81 ][ 94 ],
   alphaCSR[ 81 ][ 95 ],
   alphaCSR[ 81 ][ 96 ],
   alphaCSR[ 81 ][ 97 ],
   alphaCSR[ 81 ][ 98 ],
   alphaCSR[ 81 ][ 99 ],
   alphaCSR[ 81 ][ 100 ],
   alphaCSR[ 81 ][ 101 ],
   alphaCSR[ 81 ][ 102 ],
   alphaCSR[ 81 ][ 103 ],
   alphaCSR[ 81 ][ 104 ],
   alphaCSR[ 81 ][ 105 ],
   alphaCSR[ 81 ][ 106 ],
   alphaCSR[ 81 ][ 107 ],
   alphaCSR[ 81 ][ 108 ],
   alphaCSR[ 81 ][ 109 ],
   alphaCSR[ 81 ][ 110 ],
   alphaCSR[ 81 ][ 111 ],
   alphaCSR[ 81 ][ 112 ],
   alphaCSR[ 81 ][ 113 ],
   alphaCSR[ 81 ][ 114 ],
   alphaCSR[ 81 ][ 115 ],
   alphaCSR[ 81 ][ 116 ],
   alphaCSR[ 81 ][ 117 ],
   alphaCSR[ 81 ][ 118 ],
   alphaCSR[ 81 ][ 119 ],
   alphaCSR[ 81 ][ 120 ],
   alphaCSR[ 81 ][ 121 ],
   alphaCSR[ 81 ][ 122 ],
   alphaCSR[ 81 ][ 123 ],
   alphaCSR[ 81 ][ 124 ],
   alphaCSR[ 81 ][ 125 ],
   alphaCSR[ 81 ][ 126 ],
   alphaCSR[ 81 ][ 127 ],
   alphaCSR[ 81 ][ 128 ],
   alphaCSR[ 81 ][ 129 ],
   alphaCSR[ 81 ][ 130 ],
   alphaCSR[ 81 ][ 131 ],
   alphaCSR[ 81 ][ 132 ],
   alphaCSR[ 81 ][ 133 ],
   alphaCSR[ 81 ][ 134 ],
   alphaCSR[ 81 ][ 135 ],
   alphaCSR[ 81 ][ 136 ],
   alphaCSR[ 81 ][ 137 ],
   alphaCSR[ 81 ][ 138 ],
   alphaCSR[ 81 ][ 139 ],
   alphaCSR[ 81 ][ 140 ],
   alphaCSR[ 81 ][ 141 ],
   alphaCSR[ 81 ][ 142 ],
   alphaCSR[ 81 ][ 143 ],
   alphaCSR[ 81 ][ 144 ],
   alphaCSR[ 81 ][ 145 ],
   alphaCSR[ 81 ][ 146 ],
   alphaCSR[ 81 ][ 147 ],
   alphaCSR[ 81 ][ 148 ],
   alphaCSR[ 81 ][ 149 ],
   alphaCSR[ 81 ][ 150 ],
   alphaCSR[ 81 ][ 151 ],
   alphaCSR[ 81 ][ 152 ],
   alphaCSR[ 81 ][ 153 ],
   alphaCSR[ 81 ][ 154 ],
   alphaCSR[ 81 ][ 155 ],
   alphaCSR[ 81 ][ 156 ],
   alphaCSR[ 81 ][ 157 ],
   alphaCSR[ 81 ][ 158 ],
   alphaCSR[ 81 ][ 159 ],
   alphaCSR[ 81 ][ 160 ],
   alphaCSR[ 81 ][ 161 ],
   alphaCSR[ 81 ][ 162 ],
   alphaCSR[ 81 ][ 163 ],
   alphaCSR[ 81 ][ 164 ],
   alphaCSR[ 81 ][ 165 ],
   alphaCSR[ 81 ][ 166 ],
   alphaCSR[ 81 ][ 167 ],
   alphaCSR[ 81 ][ 168 ],
   alphaCSR[ 81 ][ 169 ],
   alphaCSR[ 81 ][ 170 ],
   alphaCSR[ 81 ][ 171 ],
   alphaCSR[ 81 ][ 172 ],
   alphaCSR[ 81 ][ 173 ],
   alphaCSR[ 81 ][ 174 ],
   alphaCSR[ 81 ][ 175 ],
   alphaCSR[ 81 ][ 176 ],
   alphaCSR[ 81 ][ 177 ],
   alphaCSR[ 81 ][ 178 ],
   alphaCSR[ 81 ][ 179 ],
   alphaCSR[ 81 ][ 180 ],
   alphaCSR[ 81 ][ 181 ],
   alphaCSR[ 81 ][ 182 ],
   alphaCSR[ 81 ][ 183 ],
   alphaCSR[ 81 ][ 184 ],
   alphaCSR[ 81 ][ 185 ],
   alphaCSR[ 81 ][ 186 ],
   alphaCSR[ 81 ][ 187 ],
   alphaCSR[ 81 ][ 188 ],
   alphaCSR[ 81 ][ 189 ],
   alphaCSR[ 81 ][ 190 ],
   alphaCSR[ 81 ][ 191 ],
   alphaCSR[ 81 ][ 192 ],
   alphaCSR[ 81 ][ 193 ],
   alphaCSR[ 81 ][ 194 ],
   alphaCSR[ 81 ][ 195 ],
   alphaCSR[ 81 ][ 196 ],
   alphaCSR[ 81 ][ 197 ],
   alphaCSR[ 81 ][ 198 ],
   alphaCSR[ 81 ][ 199 ],
   alphaCSR[ 81 ][ 200 ],
   alphaCSR[ 81 ][ 201 ],
   alphaCSR[ 81 ][ 202 ],
   alphaCSR[ 81 ][ 203 ],
   alphaCSR[ 81 ][ 204 ],
   alphaCSR[ 81 ][ 205 ],
   alphaCSR[ 81 ][ 206 ],
   alphaCSR[ 81 ][ 207 ],
   alphaCSR[ 81 ][ 208 ],
   alphaCSR[ 81 ][ 209 ],
   alphaCSR[ 81 ][ 210 ],
   alphaCSR[ 81 ][ 211 ],
   alphaCSR[ 81 ][ 212 ],
   alphaCSR[ 81 ][ 213 ],
   alphaCSR[ 81 ][ 214 ],
   alphaCSR[ 81 ][ 215 ],
   alphaCSR[ 81 ][ 216 ],
   alphaCSR[ 81 ][ 217 ],
   alphaCSR[ 81 ][ 218 ],
   alphaCSR[ 81 ][ 219 ],
   alphaCSR[ 81 ][ 220 ],
   alphaCSR[ 81 ][ 221 ],
   alphaCSR[ 81 ][ 222 ],
   alphaCSR[ 81 ][ 223 ],
   alphaCSR[ 81 ][ 224 ],
   alphaCSR[ 81 ][ 225 ],
   alphaCSR[ 81 ][ 226 ],
   alphaCSR[ 81 ][ 227 ],
   alphaCSR[ 81 ][ 228 ],
   alphaCSR[ 81 ][ 229 ],
   alphaCSR[ 81 ][ 230 ],
   alphaCSR[ 81 ][ 231 ],
   alphaCSR[ 81 ][ 232 ],
   alphaCSR[ 81 ][ 233 ],
   alphaCSR[ 81 ][ 234 ],
   alphaCSR[ 81 ][ 235 ],
   alphaCSR[ 81 ][ 236 ],
   alphaCSR[ 81 ][ 237 ],
   alphaCSR[ 81 ][ 238 ],
   alphaCSR[ 81 ][ 239 ],
   alphaCSR[ 81 ][ 240 ],
   alphaCSR[ 81 ][ 241 ],
   alphaCSR[ 81 ][ 242 ],
   alphaCSR[ 81 ][ 243 ],
   alphaCSR[ 81 ][ 244 ],
   alphaCSR[ 81 ][ 245 ],
   alphaCSR[ 81 ][ 246 ],
   alphaCSR[ 81 ][ 247 ],
   alphaCSR[ 81 ][ 248 ],
   alphaCSR[ 81 ][ 249 ],
   alphaCSR[ 81 ][ 250 ],
   alphaCSR[ 81 ][ 251 ],
   alphaCSR[ 81 ][ 252 ],
   alphaCSR[ 81 ][ 253 ],
   alphaCSR[ 81 ][ 254 ],
   alphaCSR[ 81 ][ 255 ],
   alphaCSR[ 81 ][ 256 ],
   alphaCSR[ 81 ][ 257 ],
   alphaCSR[ 81 ][ 258 ],
   alphaCSR[ 81 ][ 259 ],
   alphaCSR[ 81 ][ 260 ],
   alphaCSR[ 81 ][ 261 ],
   alphaCSR[ 81 ][ 262 ],
   alphaCSR[ 81 ][ 263 ],
   alphaCSR[ 81 ][ 264 ],
   alphaCSR[ 81 ][ 265 ],
   alphaCSR[ 81 ][ 266 ],
   alphaCSR[ 81 ][ 267 ],
   alphaCSR[ 81 ][ 268 ],
   alphaCSR[ 81 ][ 269 ],
   alphaCSR[ 81 ][ 270 ],
   alphaCSR[ 81 ][ 271 ],
   alphaCSR[ 81 ][ 272 ],
   alphaCSR[ 81 ][ 273 ],
   alphaCSR[ 81 ][ 274 ],
   alphaCSR[ 81 ][ 275 ],
   alphaCSR[ 81 ][ 276 ],
   alphaCSR[ 81 ][ 277 ],
   alphaCSR[ 81 ][ 278 ],
   alphaCSR[ 81 ][ 279 ],
   alphaCSR[ 81 ][ 280 ],
   alphaCSR[ 81 ][ 281 ],
   alphaCSR[ 81 ][ 282 ],
   alphaCSR[ 81 ][ 283 ],
   alphaCSR[ 81 ][ 284 ],
   alphaCSR[ 81 ][ 285 ],
   alphaCSR[ 81 ][ 286 ],
   alphaCSR[ 81 ][ 287 ],
   alphaCSR[ 81 ][ 288 ],
   alphaCSR[ 81 ][ 289 ],
   alphaCSR[ 81 ][ 290 ],
   alphaCSR[ 81 ][ 291 ],
   alphaCSR[ 81 ][ 292 ],
   alphaCSR[ 81 ][ 293 ],
   alphaCSR[ 81 ][ 294 ],
   alphaCSR[ 81 ][ 295 ],
   alphaCSR[ 81 ][ 296 ],
   alphaCSR[ 81 ][ 297 ],
   alphaCSR[ 81 ][ 298 ],
   alphaCSR[ 81 ][ 299 ],
   alphaCSR[ 81 ][ 300 ],
   alphaCSR[ 81 ][ 301 ],
   alphaCSR[ 81 ][ 302 ],
   alphaCSR[ 81 ][ 303 ],
   alphaCSR[ 81 ][ 304 ],
   alphaCSR[ 81 ][ 305 ],
   alphaCSR[ 81 ][ 306 ],
   alphaCSR[ 81 ][ 307 ],
   alphaCSR[ 81 ][ 308 ],
   alphaCSR[ 81 ][ 309 ],
   alphaCSR[ 81 ][ 310 ],
   alphaCSR[ 81 ][ 311 ],
   alphaCSR[ 81 ][ 312 ],
   alphaCSR[ 81 ][ 313 ],
   alphaCSR[ 81 ][ 314 ],
   alphaCSR[ 81 ][ 315 ],
   alphaCSR[ 81 ][ 316 ],
   alphaCSR[ 81 ][ 317 ],
   alphaCSR[ 81 ][ 318 ],
   alphaCSR[ 81 ][ 319 ],
   alphaCSR[ 81 ][ 320 ],
   alphaCSR[ 81 ][ 321 ],
   alphaCSR[ 81 ][ 322 ],
   alphaCSR[ 81 ][ 323 ],
   alphaCSR[ 81 ][ 324 ],
   alphaCSR[ 81 ][ 325 ],
   alphaCSR[ 81 ][ 326 ],
   alphaCSR[ 81 ][ 327 ],
   alphaCSR[ 81 ][ 328 ],
   alphaCSR[ 81 ][ 329 ],
   alphaCSR[ 81 ][ 330 ],
   alphaCSR[ 81 ][ 331 ],
   alphaCSR[ 81 ][ 332 ],
   alphaCSR[ 81 ][ 333 ],
   alphaCSR[ 81 ][ 334 ],
   alphaCSR[ 81 ][ 335 ],
   alphaCSR[ 81 ][ 336 ],
   alphaCSR[ 81 ][ 337 ],
   alphaCSR[ 81 ][ 338 ],
   alphaCSR[ 81 ][ 339 ],
   alphaCSR[ 81 ][ 340 ],
   alphaCSR[ 81 ][ 341 ],
   alphaCSR[ 81 ][ 342 ],
   alphaCSR[ 81 ][ 343 ],
   alphaCSR[ 81 ][ 344 ],
   alphaCSR[ 81 ][ 345 ],
   alphaCSR[ 81 ][ 346 ],
   alphaCSR[ 81 ][ 347 ],
   alphaCSR[ 81 ][ 348 ],
   alphaCSR[ 81 ][ 349 ],
   alphaCSR[ 81 ][ 350 ],
   alphaCSR[ 81 ][ 351 ],
   alphaCSR[ 81 ][ 352 ],
   alphaCSR[ 81 ][ 353 ],
   alphaCSR[ 81 ][ 354 ],
   alphaCSR[ 81 ][ 355 ],
   alphaCSR[ 81 ][ 356 ],
   alphaCSR[ 81 ][ 357 ],
   alphaCSR[ 81 ][ 358 ],
   alphaCSR[ 81 ][ 359 ],
   alphaCSR[ 81 ][ 360 ],
   alphaCSR[ 81 ][ 361 ],
   alphaCSR[ 81 ][ 362 ],
   alphaCSR[ 81 ][ 363 ],
   alphaCSR[ 81 ][ 364 ],
   alphaCSR[ 81 ][ 365 ],
   alphaCSR[ 81 ][ 366 ],
   alphaCSR[ 81 ][ 367 ],
   alphaCSR[ 81 ][ 368 ],
   alphaCSR[ 81 ][ 369 ],
   alphaCSR[ 81 ][ 370 ],
   alphaCSR[ 81 ][ 371 ],
   alphaCSR[ 81 ][ 372 ],
   alphaCSR[ 81 ][ 373 ],
   alphaCSR[ 81 ][ 374 ],
   alphaCSR[ 81 ][ 375 ],
   alphaCSR[ 81 ][ 376 ],
   alphaCSR[ 81 ][ 377 ],
   alphaCSR[ 81 ][ 378 ],
   alphaCSR[ 81 ][ 379 ],
   alphaCSR[ 81 ][ 380 ],
   alphaCSR[ 81 ][ 381 ],
   alphaCSR[ 81 ][ 382 ],
   alphaCSR[ 81 ][ 383 ],
   alphaCSR[ 82 ][ 0 ],
   alphaCSR[ 82 ][ 1 ],
   alphaCSR[ 82 ][ 2 ],
   alphaCSR[ 82 ][ 3 ],
   alphaCSR[ 82 ][ 4 ],
   alphaCSR[ 82 ][ 5 ],
   alphaCSR[ 82 ][ 6 ],
   alphaCSR[ 82 ][ 7 ],
   alphaCSR[ 82 ][ 8 ],
   alphaCSR[ 82 ][ 9 ],
   alphaCSR[ 82 ][ 10 ],
   alphaCSR[ 82 ][ 11 ],
   alphaCSR[ 82 ][ 12 ],
   alphaCSR[ 82 ][ 13 ],
   alphaCSR[ 82 ][ 14 ],
   alphaCSR[ 82 ][ 15 ],
   alphaCSR[ 82 ][ 16 ],
   alphaCSR[ 82 ][ 17 ],
   alphaCSR[ 82 ][ 18 ],
   alphaCSR[ 82 ][ 19 ],
   alphaCSR[ 82 ][ 20 ],
   alphaCSR[ 82 ][ 21 ],
   alphaCSR[ 82 ][ 22 ],
   alphaCSR[ 82 ][ 23 ],
   alphaCSR[ 82 ][ 24 ],
   alphaCSR[ 82 ][ 25 ],
   alphaCSR[ 82 ][ 26 ],
   alphaCSR[ 82 ][ 27 ],
   alphaCSR[ 82 ][ 28 ],
   alphaCSR[ 82 ][ 29 ],
   alphaCSR[ 82 ][ 30 ],
   alphaCSR[ 82 ][ 31 ],
   alphaCSR[ 82 ][ 32 ],
   alphaCSR[ 82 ][ 33 ],
   alphaCSR[ 82 ][ 34 ],
   alphaCSR[ 82 ][ 35 ],
   alphaCSR[ 82 ][ 36 ],
   alphaCSR[ 82 ][ 37 ],
   alphaCSR[ 82 ][ 38 ],
   alphaCSR[ 82 ][ 39 ],
   alphaCSR[ 82 ][ 40 ],
   alphaCSR[ 82 ][ 41 ],
   alphaCSR[ 82 ][ 42 ],
   alphaCSR[ 82 ][ 43 ],
   alphaCSR[ 82 ][ 44 ],
   alphaCSR[ 82 ][ 45 ],
   alphaCSR[ 82 ][ 46 ],
   alphaCSR[ 82 ][ 47 ],
   alphaCSR[ 82 ][ 48 ],
   alphaCSR[ 82 ][ 49 ],
   alphaCSR[ 82 ][ 50 ],
   alphaCSR[ 82 ][ 51 ],
   alphaCSR[ 82 ][ 52 ],
   alphaCSR[ 82 ][ 53 ],
   alphaCSR[ 82 ][ 54 ],
   alphaCSR[ 82 ][ 55 ],
   alphaCSR[ 82 ][ 56 ],
   alphaCSR[ 82 ][ 57 ],
   alphaCSR[ 82 ][ 58 ],
   alphaCSR[ 82 ][ 59 ],
   alphaCSR[ 82 ][ 60 ],
   alphaCSR[ 82 ][ 61 ],
   alphaCSR[ 82 ][ 62 ],
   alphaCSR[ 82 ][ 63 ],
   alphaCSR[ 82 ][ 64 ],
   alphaCSR[ 82 ][ 65 ],
   alphaCSR[ 82 ][ 66 ],
   alphaCSR[ 82 ][ 67 ],
   alphaCSR[ 82 ][ 68 ],
   alphaCSR[ 82 ][ 69 ],
   alphaCSR[ 82 ][ 70 ],
   alphaCSR[ 82 ][ 71 ],
   alphaCSR[ 82 ][ 72 ],
   alphaCSR[ 82 ][ 73 ],
   alphaCSR[ 82 ][ 74 ],
   alphaCSR[ 82 ][ 75 ],
   alphaCSR[ 82 ][ 76 ],
   alphaCSR[ 82 ][ 77 ],
   alphaCSR[ 82 ][ 78 ],
   alphaCSR[ 82 ][ 79 ],
   alphaCSR[ 82 ][ 80 ],
   alphaCSR[ 82 ][ 81 ],
   alphaCSR[ 82 ][ 82 ],
   alphaCSR[ 82 ][ 83 ],
   alphaCSR[ 82 ][ 84 ],
   alphaCSR[ 82 ][ 85 ],
   alphaCSR[ 82 ][ 86 ],
   alphaCSR[ 82 ][ 87 ],
   alphaCSR[ 82 ][ 88 ],
   alphaCSR[ 82 ][ 89 ],
   alphaCSR[ 82 ][ 90 ],
   alphaCSR[ 82 ][ 91 ],
   alphaCSR[ 82 ][ 92 ],
   alphaCSR[ 82 ][ 93 ],
   alphaCSR[ 82 ][ 94 ],
   alphaCSR[ 82 ][ 95 ],
   alphaCSR[ 82 ][ 96 ],
   alphaCSR[ 82 ][ 97 ],
   alphaCSR[ 82 ][ 98 ],
   alphaCSR[ 82 ][ 99 ],
   alphaCSR[ 82 ][ 100 ],
   alphaCSR[ 82 ][ 101 ],
   alphaCSR[ 82 ][ 102 ],
   alphaCSR[ 82 ][ 103 ],
   alphaCSR[ 82 ][ 104 ],
   alphaCSR[ 82 ][ 105 ],
   alphaCSR[ 82 ][ 106 ],
   alphaCSR[ 82 ][ 107 ],
   alphaCSR[ 82 ][ 108 ],
   alphaCSR[ 82 ][ 109 ],
   alphaCSR[ 82 ][ 110 ],
   alphaCSR[ 82 ][ 111 ],
   alphaCSR[ 82 ][ 112 ],
   alphaCSR[ 82 ][ 113 ],
   alphaCSR[ 82 ][ 114 ],
   alphaCSR[ 82 ][ 115 ],
   alphaCSR[ 82 ][ 116 ],
   alphaCSR[ 82 ][ 117 ],
   alphaCSR[ 82 ][ 118 ],
   alphaCSR[ 82 ][ 119 ],
   alphaCSR[ 82 ][ 120 ],
   alphaCSR[ 82 ][ 121 ],
   alphaCSR[ 82 ][ 122 ],
   alphaCSR[ 82 ][ 123 ],
   alphaCSR[ 82 ][ 124 ],
   alphaCSR[ 82 ][ 125 ],
   alphaCSR[ 82 ][ 126 ],
   alphaCSR[ 82 ][ 127 ],
   alphaCSR[ 82 ][ 128 ],
   alphaCSR[ 82 ][ 129 ],
   alphaCSR[ 82 ][ 130 ],
   alphaCSR[ 82 ][ 131 ],
   alphaCSR[ 82 ][ 132 ],
   alphaCSR[ 82 ][ 133 ],
   alphaCSR[ 82 ][ 134 ],
   alphaCSR[ 82 ][ 135 ],
   alphaCSR[ 82 ][ 136 ],
   alphaCSR[ 82 ][ 137 ],
   alphaCSR[ 82 ][ 138 ],
   alphaCSR[ 82 ][ 139 ],
   alphaCSR[ 82 ][ 140 ],
   alphaCSR[ 82 ][ 141 ],
   alphaCSR[ 82 ][ 142 ],
   alphaCSR[ 82 ][ 143 ],
   alphaCSR[ 82 ][ 144 ],
   alphaCSR[ 82 ][ 145 ],
   alphaCSR[ 82 ][ 146 ],
   alphaCSR[ 82 ][ 147 ],
   alphaCSR[ 82 ][ 148 ],
   alphaCSR[ 82 ][ 149 ],
   alphaCSR[ 82 ][ 150 ],
   alphaCSR[ 82 ][ 151 ],
   alphaCSR[ 82 ][ 152 ],
   alphaCSR[ 82 ][ 153 ],
   alphaCSR[ 82 ][ 154 ],
   alphaCSR[ 82 ][ 155 ],
   alphaCSR[ 82 ][ 156 ],
   alphaCSR[ 82 ][ 157 ],
   alphaCSR[ 82 ][ 158 ],
   alphaCSR[ 82 ][ 159 ],
   alphaCSR[ 82 ][ 160 ],
   alphaCSR[ 82 ][ 161 ],
   alphaCSR[ 82 ][ 162 ],
   alphaCSR[ 82 ][ 163 ],
   alphaCSR[ 82 ][ 164 ],
   alphaCSR[ 82 ][ 165 ],
   alphaCSR[ 82 ][ 166 ],
   alphaCSR[ 82 ][ 167 ],
   alphaCSR[ 82 ][ 168 ],
   alphaCSR[ 82 ][ 169 ],
   alphaCSR[ 82 ][ 170 ],
   alphaCSR[ 82 ][ 171 ],
   alphaCSR[ 82 ][ 172 ],
   alphaCSR[ 82 ][ 173 ],
   alphaCSR[ 82 ][ 174 ],
   alphaCSR[ 82 ][ 175 ],
   alphaCSR[ 82 ][ 176 ],
   alphaCSR[ 82 ][ 177 ],
   alphaCSR[ 82 ][ 178 ],
   alphaCSR[ 82 ][ 179 ],
   alphaCSR[ 82 ][ 180 ],
   alphaCSR[ 82 ][ 181 ],
   alphaCSR[ 82 ][ 182 ],
   alphaCSR[ 82 ][ 183 ],
   alphaCSR[ 82 ][ 184 ],
   alphaCSR[ 82 ][ 185 ],
   alphaCSR[ 82 ][ 186 ],
   alphaCSR[ 82 ][ 187 ],
   alphaCSR[ 82 ][ 188 ],
   alphaCSR[ 82 ][ 189 ],
   alphaCSR[ 82 ][ 190 ],
   alphaCSR[ 82 ][ 191 ],
   alphaCSR[ 82 ][ 192 ],
   alphaCSR[ 82 ][ 193 ],
   alphaCSR[ 82 ][ 194 ],
   alphaCSR[ 82 ][ 195 ],
   alphaCSR[ 82 ][ 196 ],
   alphaCSR[ 82 ][ 197 ],
   alphaCSR[ 82 ][ 198 ],
   alphaCSR[ 82 ][ 199 ],
   alphaCSR[ 82 ][ 200 ],
   alphaCSR[ 82 ][ 201 ],
   alphaCSR[ 82 ][ 202 ],
   alphaCSR[ 82 ][ 203 ],
   alphaCSR[ 82 ][ 204 ],
   alphaCSR[ 82 ][ 205 ],
   alphaCSR[ 82 ][ 206 ],
   alphaCSR[ 82 ][ 207 ],
   alphaCSR[ 82 ][ 208 ],
   alphaCSR[ 82 ][ 209 ],
   alphaCSR[ 82 ][ 210 ],
   alphaCSR[ 82 ][ 211 ],
   alphaCSR[ 82 ][ 212 ],
   alphaCSR[ 82 ][ 213 ],
   alphaCSR[ 82 ][ 214 ],
   alphaCSR[ 82 ][ 215 ],
   alphaCSR[ 82 ][ 216 ],
   alphaCSR[ 82 ][ 217 ],
   alphaCSR[ 82 ][ 218 ],
   alphaCSR[ 82 ][ 219 ],
   alphaCSR[ 82 ][ 220 ],
   alphaCSR[ 82 ][ 221 ],
   alphaCSR[ 82 ][ 222 ],
   alphaCSR[ 82 ][ 223 ],
   alphaCSR[ 82 ][ 224 ],
   alphaCSR[ 82 ][ 225 ],
   alphaCSR[ 82 ][ 226 ],
   alphaCSR[ 82 ][ 227 ],
   alphaCSR[ 82 ][ 228 ],
   alphaCSR[ 82 ][ 229 ],
   alphaCSR[ 82 ][ 230 ],
   alphaCSR[ 82 ][ 231 ],
   alphaCSR[ 82 ][ 232 ],
   alphaCSR[ 82 ][ 233 ],
   alphaCSR[ 82 ][ 234 ],
   alphaCSR[ 82 ][ 235 ],
   alphaCSR[ 82 ][ 236 ],
   alphaCSR[ 82 ][ 237 ],
   alphaCSR[ 82 ][ 238 ],
   alphaCSR[ 82 ][ 239 ],
   alphaCSR[ 82 ][ 240 ],
   alphaCSR[ 82 ][ 241 ],
   alphaCSR[ 82 ][ 242 ],
   alphaCSR[ 82 ][ 243 ],
   alphaCSR[ 82 ][ 244 ],
   alphaCSR[ 82 ][ 245 ],
   alphaCSR[ 82 ][ 246 ],
   alphaCSR[ 82 ][ 247 ],
   alphaCSR[ 82 ][ 248 ],
   alphaCSR[ 82 ][ 249 ],
   alphaCSR[ 82 ][ 250 ],
   alphaCSR[ 82 ][ 251 ],
   alphaCSR[ 82 ][ 252 ],
   alphaCSR[ 82 ][ 253 ],
   alphaCSR[ 82 ][ 254 ],
   alphaCSR[ 82 ][ 255 ],
   alphaCSR[ 82 ][ 256 ],
   alphaCSR[ 82 ][ 257 ],
   alphaCSR[ 82 ][ 258 ],
   alphaCSR[ 82 ][ 259 ],
   alphaCSR[ 82 ][ 260 ],
   alphaCSR[ 82 ][ 261 ],
   alphaCSR[ 82 ][ 262 ],
   alphaCSR[ 82 ][ 263 ],
   alphaCSR[ 82 ][ 264 ],
   alphaCSR[ 82 ][ 265 ],
   alphaCSR[ 82 ][ 266 ],
   alphaCSR[ 82 ][ 267 ],
   alphaCSR[ 82 ][ 268 ],
   alphaCSR[ 82 ][ 269 ],
   alphaCSR[ 82 ][ 270 ],
   alphaCSR[ 82 ][ 271 ],
   alphaCSR[ 82 ][ 272 ],
   alphaCSR[ 82 ][ 273 ],
   alphaCSR[ 82 ][ 274 ],
   alphaCSR[ 82 ][ 275 ],
   alphaCSR[ 82 ][ 276 ],
   alphaCSR[ 82 ][ 277 ],
   alphaCSR[ 82 ][ 278 ],
   alphaCSR[ 82 ][ 279 ],
   alphaCSR[ 82 ][ 280 ],
   alphaCSR[ 82 ][ 281 ],
   alphaCSR[ 82 ][ 282 ],
   alphaCSR[ 82 ][ 283 ],
   alphaCSR[ 82 ][ 284 ],
   alphaCSR[ 82 ][ 285 ],
   alphaCSR[ 82 ][ 286 ],
   alphaCSR[ 82 ][ 287 ],
   alphaCSR[ 82 ][ 288 ],
   alphaCSR[ 82 ][ 289 ],
   alphaCSR[ 82 ][ 290 ],
   alphaCSR[ 82 ][ 291 ],
   alphaCSR[ 82 ][ 292 ],
   alphaCSR[ 82 ][ 293 ],
   alphaCSR[ 82 ][ 294 ],
   alphaCSR[ 82 ][ 295 ],
   alphaCSR[ 82 ][ 296 ],
   alphaCSR[ 82 ][ 297 ],
   alphaCSR[ 82 ][ 298 ],
   alphaCSR[ 82 ][ 299 ],
   alphaCSR[ 82 ][ 300 ],
   alphaCSR[ 82 ][ 301 ],
   alphaCSR[ 82 ][ 302 ],
   alphaCSR[ 82 ][ 303 ],
   alphaCSR[ 82 ][ 304 ],
   alphaCSR[ 82 ][ 305 ],
   alphaCSR[ 82 ][ 306 ],
   alphaCSR[ 82 ][ 307 ],
   alphaCSR[ 82 ][ 308 ],
   alphaCSR[ 82 ][ 309 ],
   alphaCSR[ 82 ][ 310 ],
   alphaCSR[ 82 ][ 311 ],
   alphaCSR[ 82 ][ 312 ],
   alphaCSR[ 82 ][ 313 ],
   alphaCSR[ 82 ][ 314 ],
   alphaCSR[ 82 ][ 315 ],
   alphaCSR[ 82 ][ 316 ],
   alphaCSR[ 82 ][ 317 ],
   alphaCSR[ 82 ][ 318 ],
   alphaCSR[ 82 ][ 319 ],
   alphaCSR[ 82 ][ 320 ],
   alphaCSR[ 82 ][ 321 ],
   alphaCSR[ 82 ][ 322 ],
   alphaCSR[ 82 ][ 323 ],
   alphaCSR[ 82 ][ 324 ],
   alphaCSR[ 82 ][ 325 ],
   alphaCSR[ 82 ][ 326 ],
   alphaCSR[ 82 ][ 327 ],
   alphaCSR[ 82 ][ 328 ],
   alphaCSR[ 82 ][ 329 ],
   alphaCSR[ 82 ][ 330 ],
   alphaCSR[ 82 ][ 331 ],
   alphaCSR[ 82 ][ 332 ],
   alphaCSR[ 82 ][ 333 ],
   alphaCSR[ 82 ][ 334 ],
   alphaCSR[ 82 ][ 335 ],
   alphaCSR[ 82 ][ 336 ],
   alphaCSR[ 82 ][ 337 ],
   alphaCSR[ 82 ][ 338 ],
   alphaCSR[ 82 ][ 339 ],
   alphaCSR[ 82 ][ 340 ],
   alphaCSR[ 82 ][ 341 ],
   alphaCSR[ 82 ][ 342 ],
   alphaCSR[ 82 ][ 343 ],
   alphaCSR[ 82 ][ 344 ],
   alphaCSR[ 82 ][ 345 ],
   alphaCSR[ 82 ][ 346 ],
   alphaCSR[ 82 ][ 347 ],
   alphaCSR[ 82 ][ 348 ],
   alphaCSR[ 82 ][ 349 ],
   alphaCSR[ 82 ][ 350 ],
   alphaCSR[ 82 ][ 351 ],
   alphaCSR[ 82 ][ 352 ],
   alphaCSR[ 82 ][ 353 ],
   alphaCSR[ 82 ][ 354 ],
   alphaCSR[ 82 ][ 355 ],
   alphaCSR[ 82 ][ 356 ],
   alphaCSR[ 82 ][ 357 ],
   alphaCSR[ 82 ][ 358 ],
   alphaCSR[ 82 ][ 359 ],
   alphaCSR[ 82 ][ 360 ],
   alphaCSR[ 82 ][ 361 ],
   alphaCSR[ 82 ][ 362 ],
   alphaCSR[ 82 ][ 363 ],
   alphaCSR[ 82 ][ 364 ],
   alphaCSR[ 82 ][ 365 ],
   alphaCSR[ 82 ][ 366 ],
   alphaCSR[ 82 ][ 367 ],
   alphaCSR[ 82 ][ 368 ],
   alphaCSR[ 82 ][ 369 ],
   alphaCSR[ 82 ][ 370 ],
   alphaCSR[ 82 ][ 371 ],
   alphaCSR[ 82 ][ 372 ],
   alphaCSR[ 82 ][ 373 ],
   alphaCSR[ 82 ][ 374 ],
   alphaCSR[ 82 ][ 375 ],
   alphaCSR[ 82 ][ 376 ],
   alphaCSR[ 82 ][ 377 ],
   alphaCSR[ 82 ][ 378 ],
   alphaCSR[ 82 ][ 379 ],
   alphaCSR[ 82 ][ 380 ],
   alphaCSR[ 82 ][ 381 ],
   alphaCSR[ 82 ][ 382 ],
   alphaCSR[ 82 ][ 383 ],
   alphaCSR[ 83 ][ 0 ],
   alphaCSR[ 83 ][ 1 ],
   alphaCSR[ 83 ][ 2 ],
   alphaCSR[ 83 ][ 3 ],
   alphaCSR[ 83 ][ 4 ],
   alphaCSR[ 83 ][ 5 ],
   alphaCSR[ 83 ][ 6 ],
   alphaCSR[ 83 ][ 7 ],
   alphaCSR[ 83 ][ 8 ],
   alphaCSR[ 83 ][ 9 ],
   alphaCSR[ 83 ][ 10 ],
   alphaCSR[ 83 ][ 11 ],
   alphaCSR[ 83 ][ 12 ],
   alphaCSR[ 83 ][ 13 ],
   alphaCSR[ 83 ][ 14 ],
   alphaCSR[ 83 ][ 15 ],
   alphaCSR[ 83 ][ 16 ],
   alphaCSR[ 83 ][ 17 ],
   alphaCSR[ 83 ][ 18 ],
   alphaCSR[ 83 ][ 19 ],
   alphaCSR[ 83 ][ 20 ],
   alphaCSR[ 83 ][ 21 ],
   alphaCSR[ 83 ][ 22 ],
   alphaCSR[ 83 ][ 23 ],
   alphaCSR[ 83 ][ 24 ],
   alphaCSR[ 83 ][ 25 ],
   alphaCSR[ 83 ][ 26 ],
   alphaCSR[ 83 ][ 27 ],
   alphaCSR[ 83 ][ 28 ],
   alphaCSR[ 83 ][ 29 ],
   alphaCSR[ 83 ][ 30 ],
   alphaCSR[ 83 ][ 31 ],
   alphaCSR[ 83 ][ 32 ],
   alphaCSR[ 83 ][ 33 ],
   alphaCSR[ 83 ][ 34 ],
   alphaCSR[ 83 ][ 35 ],
   alphaCSR[ 83 ][ 36 ],
   alphaCSR[ 83 ][ 37 ],
   alphaCSR[ 83 ][ 38 ],
   alphaCSR[ 83 ][ 39 ],
   alphaCSR[ 83 ][ 40 ],
   alphaCSR[ 83 ][ 41 ],
   alphaCSR[ 83 ][ 42 ],
   alphaCSR[ 83 ][ 43 ],
   alphaCSR[ 83 ][ 44 ],
   alphaCSR[ 83 ][ 45 ],
   alphaCSR[ 83 ][ 46 ],
   alphaCSR[ 83 ][ 47 ],
   alphaCSR[ 83 ][ 48 ],
   alphaCSR[ 83 ][ 49 ],
   alphaCSR[ 83 ][ 50 ],
   alphaCSR[ 83 ][ 51 ],
   alphaCSR[ 83 ][ 52 ],
   alphaCSR[ 83 ][ 53 ],
   alphaCSR[ 83 ][ 54 ],
   alphaCSR[ 83 ][ 55 ],
   alphaCSR[ 83 ][ 56 ],
   alphaCSR[ 83 ][ 57 ],
   alphaCSR[ 83 ][ 58 ],
   alphaCSR[ 83 ][ 59 ],
   alphaCSR[ 83 ][ 60 ],
   alphaCSR[ 83 ][ 61 ],
   alphaCSR[ 83 ][ 62 ],
   alphaCSR[ 83 ][ 63 ],
   alphaCSR[ 83 ][ 64 ],
   alphaCSR[ 83 ][ 65 ],
   alphaCSR[ 83 ][ 66 ],
   alphaCSR[ 83 ][ 67 ],
   alphaCSR[ 83 ][ 68 ],
   alphaCSR[ 83 ][ 69 ],
   alphaCSR[ 83 ][ 70 ],
   alphaCSR[ 83 ][ 71 ],
   alphaCSR[ 83 ][ 72 ],
   alphaCSR[ 83 ][ 73 ],
   alphaCSR[ 83 ][ 74 ],
   alphaCSR[ 83 ][ 75 ],
   alphaCSR[ 83 ][ 76 ],
   alphaCSR[ 83 ][ 77 ],
   alphaCSR[ 83 ][ 78 ],
   alphaCSR[ 83 ][ 79 ],
   alphaCSR[ 83 ][ 80 ],
   alphaCSR[ 83 ][ 81 ],
   alphaCSR[ 83 ][ 82 ],
   alphaCSR[ 83 ][ 83 ],
   alphaCSR[ 83 ][ 84 ],
   alphaCSR[ 83 ][ 85 ],
   alphaCSR[ 83 ][ 86 ],
   alphaCSR[ 83 ][ 87 ],
   alphaCSR[ 83 ][ 88 ],
   alphaCSR[ 83 ][ 89 ],
   alphaCSR[ 83 ][ 90 ],
   alphaCSR[ 83 ][ 91 ],
   alphaCSR[ 83 ][ 92 ],
   alphaCSR[ 83 ][ 93 ],
   alphaCSR[ 83 ][ 94 ],
   alphaCSR[ 83 ][ 95 ],
   alphaCSR[ 83 ][ 96 ],
   alphaCSR[ 83 ][ 97 ],
   alphaCSR[ 83 ][ 98 ],
   alphaCSR[ 83 ][ 99 ],
   alphaCSR[ 83 ][ 100 ],
   alphaCSR[ 83 ][ 101 ],
   alphaCSR[ 83 ][ 102 ],
   alphaCSR[ 83 ][ 103 ],
   alphaCSR[ 83 ][ 104 ],
   alphaCSR[ 83 ][ 105 ],
   alphaCSR[ 83 ][ 106 ],
   alphaCSR[ 83 ][ 107 ],
   alphaCSR[ 83 ][ 108 ],
   alphaCSR[ 83 ][ 109 ],
   alphaCSR[ 83 ][ 110 ],
   alphaCSR[ 83 ][ 111 ],
   alphaCSR[ 83 ][ 112 ],
   alphaCSR[ 83 ][ 113 ],
   alphaCSR[ 83 ][ 114 ],
   alphaCSR[ 83 ][ 115 ],
   alphaCSR[ 83 ][ 116 ],
   alphaCSR[ 83 ][ 117 ],
   alphaCSR[ 83 ][ 118 ],
   alphaCSR[ 83 ][ 119 ],
   alphaCSR[ 83 ][ 120 ],
   alphaCSR[ 83 ][ 121 ],
   alphaCSR[ 83 ][ 122 ],
   alphaCSR[ 83 ][ 123 ],
   alphaCSR[ 83 ][ 124 ],
   alphaCSR[ 83 ][ 125 ],
   alphaCSR[ 83 ][ 126 ],
   alphaCSR[ 83 ][ 127 ],
   alphaCSR[ 83 ][ 128 ],
   alphaCSR[ 83 ][ 129 ],
   alphaCSR[ 83 ][ 130 ],
   alphaCSR[ 83 ][ 131 ],
   alphaCSR[ 83 ][ 132 ],
   alphaCSR[ 83 ][ 133 ],
   alphaCSR[ 83 ][ 134 ],
   alphaCSR[ 83 ][ 135 ],
   alphaCSR[ 83 ][ 136 ],
   alphaCSR[ 83 ][ 137 ],
   alphaCSR[ 83 ][ 138 ],
   alphaCSR[ 83 ][ 139 ],
   alphaCSR[ 83 ][ 140 ],
   alphaCSR[ 83 ][ 141 ],
   alphaCSR[ 83 ][ 142 ],
   alphaCSR[ 83 ][ 143 ],
   alphaCSR[ 83 ][ 144 ],
   alphaCSR[ 83 ][ 145 ],
   alphaCSR[ 83 ][ 146 ],
   alphaCSR[ 83 ][ 147 ],
   alphaCSR[ 83 ][ 148 ],
   alphaCSR[ 83 ][ 149 ],
   alphaCSR[ 83 ][ 150 ],
   alphaCSR[ 83 ][ 151 ],
   alphaCSR[ 83 ][ 152 ],
   alphaCSR[ 83 ][ 153 ],
   alphaCSR[ 83 ][ 154 ],
   alphaCSR[ 83 ][ 155 ],
   alphaCSR[ 83 ][ 156 ],
   alphaCSR[ 83 ][ 157 ],
   alphaCSR[ 83 ][ 158 ],
   alphaCSR[ 83 ][ 159 ],
   alphaCSR[ 83 ][ 160 ],
   alphaCSR[ 83 ][ 161 ],
   alphaCSR[ 83 ][ 162 ],
   alphaCSR[ 83 ][ 163 ],
   alphaCSR[ 83 ][ 164 ],
   alphaCSR[ 83 ][ 165 ],
   alphaCSR[ 83 ][ 166 ],
   alphaCSR[ 83 ][ 167 ],
   alphaCSR[ 83 ][ 168 ],
   alphaCSR[ 83 ][ 169 ],
   alphaCSR[ 83 ][ 170 ],
   alphaCSR[ 83 ][ 171 ],
   alphaCSR[ 83 ][ 172 ],
   alphaCSR[ 83 ][ 173 ],
   alphaCSR[ 83 ][ 174 ],
   alphaCSR[ 83 ][ 175 ],
   alphaCSR[ 83 ][ 176 ],
   alphaCSR[ 83 ][ 177 ],
   alphaCSR[ 83 ][ 178 ],
   alphaCSR[ 83 ][ 179 ],
   alphaCSR[ 83 ][ 180 ],
   alphaCSR[ 83 ][ 181 ],
   alphaCSR[ 83 ][ 182 ],
   alphaCSR[ 83 ][ 183 ],
   alphaCSR[ 83 ][ 184 ],
   alphaCSR[ 83 ][ 185 ],
   alphaCSR[ 83 ][ 186 ],
   alphaCSR[ 83 ][ 187 ],
   alphaCSR[ 83 ][ 188 ],
   alphaCSR[ 83 ][ 189 ],
   alphaCSR[ 83 ][ 190 ],
   alphaCSR[ 83 ][ 191 ],
   alphaCSR[ 83 ][ 192 ],
   alphaCSR[ 83 ][ 193 ],
   alphaCSR[ 83 ][ 194 ],
   alphaCSR[ 83 ][ 195 ],
   alphaCSR[ 83 ][ 196 ],
   alphaCSR[ 83 ][ 197 ],
   alphaCSR[ 83 ][ 198 ],
   alphaCSR[ 83 ][ 199 ],
   alphaCSR[ 83 ][ 200 ],
   alphaCSR[ 83 ][ 201 ],
   alphaCSR[ 83 ][ 202 ],
   alphaCSR[ 83 ][ 203 ],
   alphaCSR[ 83 ][ 204 ],
   alphaCSR[ 83 ][ 205 ],
   alphaCSR[ 83 ][ 206 ],
   alphaCSR[ 83 ][ 207 ],
   alphaCSR[ 83 ][ 208 ],
   alphaCSR[ 83 ][ 209 ],
   alphaCSR[ 83 ][ 210 ],
   alphaCSR[ 83 ][ 211 ],
   alphaCSR[ 83 ][ 212 ],
   alphaCSR[ 83 ][ 213 ],
   alphaCSR[ 83 ][ 214 ],
   alphaCSR[ 83 ][ 215 ],
   alphaCSR[ 83 ][ 216 ],
   alphaCSR[ 83 ][ 217 ],
   alphaCSR[ 83 ][ 218 ],
   alphaCSR[ 83 ][ 219 ],
   alphaCSR[ 83 ][ 220 ],
   alphaCSR[ 83 ][ 221 ],
   alphaCSR[ 83 ][ 222 ],
   alphaCSR[ 83 ][ 223 ],
   alphaCSR[ 83 ][ 224 ],
   alphaCSR[ 83 ][ 225 ],
   alphaCSR[ 83 ][ 226 ],
   alphaCSR[ 83 ][ 227 ],
   alphaCSR[ 83 ][ 228 ],
   alphaCSR[ 83 ][ 229 ],
   alphaCSR[ 83 ][ 230 ],
   alphaCSR[ 83 ][ 231 ],
   alphaCSR[ 83 ][ 232 ],
   alphaCSR[ 83 ][ 233 ],
   alphaCSR[ 83 ][ 234 ],
   alphaCSR[ 83 ][ 235 ],
   alphaCSR[ 83 ][ 236 ],
   alphaCSR[ 83 ][ 237 ],
   alphaCSR[ 83 ][ 238 ],
   alphaCSR[ 83 ][ 239 ],
   alphaCSR[ 83 ][ 240 ],
   alphaCSR[ 83 ][ 241 ],
   alphaCSR[ 83 ][ 242 ],
   alphaCSR[ 83 ][ 243 ],
   alphaCSR[ 83 ][ 244 ],
   alphaCSR[ 83 ][ 245 ],
   alphaCSR[ 83 ][ 246 ],
   alphaCSR[ 83 ][ 247 ],
   alphaCSR[ 83 ][ 248 ],
   alphaCSR[ 83 ][ 249 ],
   alphaCSR[ 83 ][ 250 ],
   alphaCSR[ 83 ][ 251 ],
   alphaCSR[ 83 ][ 252 ],
   alphaCSR[ 83 ][ 253 ],
   alphaCSR[ 83 ][ 254 ],
   alphaCSR[ 83 ][ 255 ],
   alphaCSR[ 83 ][ 256 ],
   alphaCSR[ 83 ][ 257 ],
   alphaCSR[ 83 ][ 258 ],
   alphaCSR[ 83 ][ 259 ],
   alphaCSR[ 83 ][ 260 ],
   alphaCSR[ 83 ][ 261 ],
   alphaCSR[ 83 ][ 262 ],
   alphaCSR[ 83 ][ 263 ],
   alphaCSR[ 83 ][ 264 ],
   alphaCSR[ 83 ][ 265 ],
   alphaCSR[ 83 ][ 266 ],
   alphaCSR[ 83 ][ 267 ],
   alphaCSR[ 83 ][ 268 ],
   alphaCSR[ 83 ][ 269 ],
   alphaCSR[ 83 ][ 270 ],
   alphaCSR[ 83 ][ 271 ],
   alphaCSR[ 83 ][ 272 ],
   alphaCSR[ 83 ][ 273 ],
   alphaCSR[ 83 ][ 274 ],
   alphaCSR[ 83 ][ 275 ],
   alphaCSR[ 83 ][ 276 ],
   alphaCSR[ 83 ][ 277 ],
   alphaCSR[ 83 ][ 278 ],
   alphaCSR[ 83 ][ 279 ],
   alphaCSR[ 83 ][ 280 ],
   alphaCSR[ 83 ][ 281 ],
   alphaCSR[ 83 ][ 282 ],
   alphaCSR[ 83 ][ 283 ],
   alphaCSR[ 83 ][ 284 ],
   alphaCSR[ 83 ][ 285 ],
   alphaCSR[ 83 ][ 286 ],
   alphaCSR[ 83 ][ 287 ],
   alphaCSR[ 83 ][ 288 ],
   alphaCSR[ 83 ][ 289 ],
   alphaCSR[ 83 ][ 290 ],
   alphaCSR[ 83 ][ 291 ],
   alphaCSR[ 83 ][ 292 ],
   alphaCSR[ 83 ][ 293 ],
   alphaCSR[ 83 ][ 294 ],
   alphaCSR[ 83 ][ 295 ],
   alphaCSR[ 83 ][ 296 ],
   alphaCSR[ 83 ][ 297 ],
   alphaCSR[ 83 ][ 298 ],
   alphaCSR[ 83 ][ 299 ],
   alphaCSR[ 83 ][ 300 ],
   alphaCSR[ 83 ][ 301 ],
   alphaCSR[ 83 ][ 302 ],
   alphaCSR[ 83 ][ 303 ],
   alphaCSR[ 83 ][ 304 ],
   alphaCSR[ 83 ][ 305 ],
   alphaCSR[ 83 ][ 306 ],
   alphaCSR[ 83 ][ 307 ],
   alphaCSR[ 83 ][ 308 ],
   alphaCSR[ 83 ][ 309 ],
   alphaCSR[ 83 ][ 310 ],
   alphaCSR[ 83 ][ 311 ],
   alphaCSR[ 83 ][ 312 ],
   alphaCSR[ 83 ][ 313 ],
   alphaCSR[ 83 ][ 314 ],
   alphaCSR[ 83 ][ 315 ],
   alphaCSR[ 83 ][ 316 ],
   alphaCSR[ 83 ][ 317 ],
   alphaCSR[ 83 ][ 318 ],
   alphaCSR[ 83 ][ 319 ],
   alphaCSR[ 83 ][ 320 ],
   alphaCSR[ 83 ][ 321 ],
   alphaCSR[ 83 ][ 322 ],
   alphaCSR[ 83 ][ 323 ],
   alphaCSR[ 83 ][ 324 ],
   alphaCSR[ 83 ][ 325 ],
   alphaCSR[ 83 ][ 326 ],
   alphaCSR[ 83 ][ 327 ],
   alphaCSR[ 83 ][ 328 ],
   alphaCSR[ 83 ][ 329 ],
   alphaCSR[ 83 ][ 330 ],
   alphaCSR[ 83 ][ 331 ],
   alphaCSR[ 83 ][ 332 ],
   alphaCSR[ 83 ][ 333 ],
   alphaCSR[ 83 ][ 334 ],
   alphaCSR[ 83 ][ 335 ],
   alphaCSR[ 83 ][ 336 ],
   alphaCSR[ 83 ][ 337 ],
   alphaCSR[ 83 ][ 338 ],
   alphaCSR[ 83 ][ 339 ],
   alphaCSR[ 83 ][ 340 ],
   alphaCSR[ 83 ][ 341 ],
   alphaCSR[ 83 ][ 342 ],
   alphaCSR[ 83 ][ 343 ],
   alphaCSR[ 83 ][ 344 ],
   alphaCSR[ 83 ][ 345 ],
   alphaCSR[ 83 ][ 346 ],
   alphaCSR[ 83 ][ 347 ],
   alphaCSR[ 83 ][ 348 ],
   alphaCSR[ 83 ][ 349 ],
   alphaCSR[ 83 ][ 350 ],
   alphaCSR[ 83 ][ 351 ],
   alphaCSR[ 83 ][ 352 ],
   alphaCSR[ 83 ][ 353 ],
   alphaCSR[ 83 ][ 354 ],
   alphaCSR[ 83 ][ 355 ],
   alphaCSR[ 83 ][ 356 ],
   alphaCSR[ 83 ][ 357 ],
   alphaCSR[ 83 ][ 358 ],
   alphaCSR[ 83 ][ 359 ],
   alphaCSR[ 83 ][ 360 ],
   alphaCSR[ 83 ][ 361 ],
   alphaCSR[ 83 ][ 362 ],
   alphaCSR[ 83 ][ 363 ],
   alphaCSR[ 83 ][ 364 ],
   alphaCSR[ 83 ][ 365 ],
   alphaCSR[ 83 ][ 366 ],
   alphaCSR[ 83 ][ 367 ],
   alphaCSR[ 83 ][ 368 ],
   alphaCSR[ 83 ][ 369 ],
   alphaCSR[ 83 ][ 370 ],
   alphaCSR[ 83 ][ 371 ],
   alphaCSR[ 83 ][ 372 ],
   alphaCSR[ 83 ][ 373 ],
   alphaCSR[ 83 ][ 374 ],
   alphaCSR[ 83 ][ 375 ],
   alphaCSR[ 83 ][ 376 ],
   alphaCSR[ 83 ][ 377 ],
   alphaCSR[ 83 ][ 378 ],
   alphaCSR[ 83 ][ 379 ],
   alphaCSR[ 83 ][ 380 ],
   alphaCSR[ 83 ][ 381 ],
   alphaCSR[ 83 ][ 382 ],
   alphaCSR[ 83 ][ 383 ],
   alphaCSR[ 84 ][ 0 ],
   alphaCSR[ 84 ][ 1 ],
   alphaCSR[ 84 ][ 2 ],
   alphaCSR[ 84 ][ 3 ],
   alphaCSR[ 84 ][ 4 ],
   alphaCSR[ 84 ][ 5 ],
   alphaCSR[ 84 ][ 6 ],
   alphaCSR[ 84 ][ 7 ],
   alphaCSR[ 84 ][ 8 ],
   alphaCSR[ 84 ][ 9 ],
   alphaCSR[ 84 ][ 10 ],
   alphaCSR[ 84 ][ 11 ],
   alphaCSR[ 84 ][ 12 ],
   alphaCSR[ 84 ][ 13 ],
   alphaCSR[ 84 ][ 14 ],
   alphaCSR[ 84 ][ 15 ],
   alphaCSR[ 84 ][ 16 ],
   alphaCSR[ 84 ][ 17 ],
   alphaCSR[ 84 ][ 18 ],
   alphaCSR[ 84 ][ 19 ],
   alphaCSR[ 84 ][ 20 ],
   alphaCSR[ 84 ][ 21 ],
   alphaCSR[ 84 ][ 22 ],
   alphaCSR[ 84 ][ 23 ],
   alphaCSR[ 84 ][ 24 ],
   alphaCSR[ 84 ][ 25 ],
   alphaCSR[ 84 ][ 26 ],
   alphaCSR[ 84 ][ 27 ],
   alphaCSR[ 84 ][ 28 ],
   alphaCSR[ 84 ][ 29 ],
   alphaCSR[ 84 ][ 30 ],
   alphaCSR[ 84 ][ 31 ],
   alphaCSR[ 84 ][ 32 ],
   alphaCSR[ 84 ][ 33 ],
   alphaCSR[ 84 ][ 34 ],
   alphaCSR[ 84 ][ 35 ],
   alphaCSR[ 84 ][ 36 ],
   alphaCSR[ 84 ][ 37 ],
   alphaCSR[ 84 ][ 38 ],
   alphaCSR[ 84 ][ 39 ],
   alphaCSR[ 84 ][ 40 ],
   alphaCSR[ 84 ][ 41 ],
   alphaCSR[ 84 ][ 42 ],
   alphaCSR[ 84 ][ 43 ],
   alphaCSR[ 84 ][ 44 ],
   alphaCSR[ 84 ][ 45 ],
   alphaCSR[ 84 ][ 46 ],
   alphaCSR[ 84 ][ 47 ],
   alphaCSR[ 84 ][ 48 ],
   alphaCSR[ 84 ][ 49 ],
   alphaCSR[ 84 ][ 50 ],
   alphaCSR[ 84 ][ 51 ],
   alphaCSR[ 84 ][ 52 ],
   alphaCSR[ 84 ][ 53 ],
   alphaCSR[ 84 ][ 54 ],
   alphaCSR[ 84 ][ 55 ],
   alphaCSR[ 84 ][ 56 ],
   alphaCSR[ 84 ][ 57 ],
   alphaCSR[ 84 ][ 58 ],
   alphaCSR[ 84 ][ 59 ],
   alphaCSR[ 84 ][ 60 ],
   alphaCSR[ 84 ][ 61 ],
   alphaCSR[ 84 ][ 62 ],
   alphaCSR[ 84 ][ 63 ],
   alphaCSR[ 84 ][ 64 ],
   alphaCSR[ 84 ][ 65 ],
   alphaCSR[ 84 ][ 66 ],
   alphaCSR[ 84 ][ 67 ],
   alphaCSR[ 84 ][ 68 ],
   alphaCSR[ 84 ][ 69 ],
   alphaCSR[ 84 ][ 70 ],
   alphaCSR[ 84 ][ 71 ],
   alphaCSR[ 84 ][ 72 ],
   alphaCSR[ 84 ][ 73 ],
   alphaCSR[ 84 ][ 74 ],
   alphaCSR[ 84 ][ 75 ],
   alphaCSR[ 84 ][ 76 ],
   alphaCSR[ 84 ][ 77 ],
   alphaCSR[ 84 ][ 78 ],
   alphaCSR[ 84 ][ 79 ],
   alphaCSR[ 84 ][ 80 ],
   alphaCSR[ 84 ][ 81 ],
   alphaCSR[ 84 ][ 82 ],
   alphaCSR[ 84 ][ 83 ],
   alphaCSR[ 84 ][ 84 ],
   alphaCSR[ 84 ][ 85 ],
   alphaCSR[ 84 ][ 86 ],
   alphaCSR[ 84 ][ 87 ],
   alphaCSR[ 84 ][ 88 ],
   alphaCSR[ 84 ][ 89 ],
   alphaCSR[ 84 ][ 90 ],
   alphaCSR[ 84 ][ 91 ],
   alphaCSR[ 84 ][ 92 ],
   alphaCSR[ 84 ][ 93 ],
   alphaCSR[ 84 ][ 94 ],
   alphaCSR[ 84 ][ 95 ],
   alphaCSR[ 84 ][ 96 ],
   alphaCSR[ 84 ][ 97 ],
   alphaCSR[ 84 ][ 98 ],
   alphaCSR[ 84 ][ 99 ],
   alphaCSR[ 84 ][ 100 ],
   alphaCSR[ 84 ][ 101 ],
   alphaCSR[ 84 ][ 102 ],
   alphaCSR[ 84 ][ 103 ],
   alphaCSR[ 84 ][ 104 ],
   alphaCSR[ 84 ][ 105 ],
   alphaCSR[ 84 ][ 106 ],
   alphaCSR[ 84 ][ 107 ],
   alphaCSR[ 84 ][ 108 ],
   alphaCSR[ 84 ][ 109 ],
   alphaCSR[ 84 ][ 110 ],
   alphaCSR[ 84 ][ 111 ],
   alphaCSR[ 84 ][ 112 ],
   alphaCSR[ 84 ][ 113 ],
   alphaCSR[ 84 ][ 114 ],
   alphaCSR[ 84 ][ 115 ],
   alphaCSR[ 84 ][ 116 ],
   alphaCSR[ 84 ][ 117 ],
   alphaCSR[ 84 ][ 118 ],
   alphaCSR[ 84 ][ 119 ],
   alphaCSR[ 84 ][ 120 ],
   alphaCSR[ 84 ][ 121 ],
   alphaCSR[ 84 ][ 122 ],
   alphaCSR[ 84 ][ 123 ],
   alphaCSR[ 84 ][ 124 ],
   alphaCSR[ 84 ][ 125 ],
   alphaCSR[ 84 ][ 126 ],
   alphaCSR[ 84 ][ 127 ],
   alphaCSR[ 84 ][ 128 ],
   alphaCSR[ 84 ][ 129 ],
   alphaCSR[ 84 ][ 130 ],
   alphaCSR[ 84 ][ 131 ],
   alphaCSR[ 84 ][ 132 ],
   alphaCSR[ 84 ][ 133 ],
   alphaCSR[ 84 ][ 134 ],
   alphaCSR[ 84 ][ 135 ],
   alphaCSR[ 84 ][ 136 ],
   alphaCSR[ 84 ][ 137 ],
   alphaCSR[ 84 ][ 138 ],
   alphaCSR[ 84 ][ 139 ],
   alphaCSR[ 84 ][ 140 ],
   alphaCSR[ 84 ][ 141 ],
   alphaCSR[ 84 ][ 142 ],
   alphaCSR[ 84 ][ 143 ],
   alphaCSR[ 84 ][ 144 ],
   alphaCSR[ 84 ][ 145 ],
   alphaCSR[ 84 ][ 146 ],
   alphaCSR[ 84 ][ 147 ],
   alphaCSR[ 84 ][ 148 ],
   alphaCSR[ 84 ][ 149 ],
   alphaCSR[ 84 ][ 150 ],
   alphaCSR[ 84 ][ 151 ],
   alphaCSR[ 84 ][ 152 ],
   alphaCSR[ 84 ][ 153 ],
   alphaCSR[ 84 ][ 154 ],
   alphaCSR[ 84 ][ 155 ],
   alphaCSR[ 84 ][ 156 ],
   alphaCSR[ 84 ][ 157 ],
   alphaCSR[ 84 ][ 158 ],
   alphaCSR[ 84 ][ 159 ],
   alphaCSR[ 84 ][ 160 ],
   alphaCSR[ 84 ][ 161 ],
   alphaCSR[ 84 ][ 162 ],
   alphaCSR[ 84 ][ 163 ],
   alphaCSR[ 84 ][ 164 ],
   alphaCSR[ 84 ][ 165 ],
   alphaCSR[ 84 ][ 166 ],
   alphaCSR[ 84 ][ 167 ],
   alphaCSR[ 84 ][ 168 ],
   alphaCSR[ 84 ][ 169 ],
   alphaCSR[ 84 ][ 170 ],
   alphaCSR[ 84 ][ 171 ],
   alphaCSR[ 84 ][ 172 ],
   alphaCSR[ 84 ][ 173 ],
   alphaCSR[ 84 ][ 174 ],
   alphaCSR[ 84 ][ 175 ],
   alphaCSR[ 84 ][ 176 ],
   alphaCSR[ 84 ][ 177 ],
   alphaCSR[ 84 ][ 178 ],
   alphaCSR[ 84 ][ 179 ],
   alphaCSR[ 84 ][ 180 ],
   alphaCSR[ 84 ][ 181 ],
   alphaCSR[ 84 ][ 182 ],
   alphaCSR[ 84 ][ 183 ],
   alphaCSR[ 84 ][ 184 ],
   alphaCSR[ 84 ][ 185 ],
   alphaCSR[ 84 ][ 186 ],
   alphaCSR[ 84 ][ 187 ],
   alphaCSR[ 84 ][ 188 ],
   alphaCSR[ 84 ][ 189 ],
   alphaCSR[ 84 ][ 190 ],
   alphaCSR[ 84 ][ 191 ],
   alphaCSR[ 84 ][ 192 ],
   alphaCSR[ 84 ][ 193 ],
   alphaCSR[ 84 ][ 194 ],
   alphaCSR[ 84 ][ 195 ],
   alphaCSR[ 84 ][ 196 ],
   alphaCSR[ 84 ][ 197 ],
   alphaCSR[ 84 ][ 198 ],
   alphaCSR[ 84 ][ 199 ],
   alphaCSR[ 84 ][ 200 ],
   alphaCSR[ 84 ][ 201 ],
   alphaCSR[ 84 ][ 202 ],
   alphaCSR[ 84 ][ 203 ],
   alphaCSR[ 84 ][ 204 ],
   alphaCSR[ 84 ][ 205 ],
   alphaCSR[ 84 ][ 206 ],
   alphaCSR[ 84 ][ 207 ],
   alphaCSR[ 84 ][ 208 ],
   alphaCSR[ 84 ][ 209 ],
   alphaCSR[ 84 ][ 210 ],
   alphaCSR[ 84 ][ 211 ],
   alphaCSR[ 84 ][ 212 ],
   alphaCSR[ 84 ][ 213 ],
   alphaCSR[ 84 ][ 214 ],
   alphaCSR[ 84 ][ 215 ],
   alphaCSR[ 84 ][ 216 ],
   alphaCSR[ 84 ][ 217 ],
   alphaCSR[ 84 ][ 218 ],
   alphaCSR[ 84 ][ 219 ],
   alphaCSR[ 84 ][ 220 ],
   alphaCSR[ 84 ][ 221 ],
   alphaCSR[ 84 ][ 222 ],
   alphaCSR[ 84 ][ 223 ],
   alphaCSR[ 84 ][ 224 ],
   alphaCSR[ 84 ][ 225 ],
   alphaCSR[ 84 ][ 226 ],
   alphaCSR[ 84 ][ 227 ],
   alphaCSR[ 84 ][ 228 ],
   alphaCSR[ 84 ][ 229 ],
   alphaCSR[ 84 ][ 230 ],
   alphaCSR[ 84 ][ 231 ],
   alphaCSR[ 84 ][ 232 ],
   alphaCSR[ 84 ][ 233 ],
   alphaCSR[ 84 ][ 234 ],
   alphaCSR[ 84 ][ 235 ],
   alphaCSR[ 84 ][ 236 ],
   alphaCSR[ 84 ][ 237 ],
   alphaCSR[ 84 ][ 238 ],
   alphaCSR[ 84 ][ 239 ],
   alphaCSR[ 84 ][ 240 ],
   alphaCSR[ 84 ][ 241 ],
   alphaCSR[ 84 ][ 242 ],
   alphaCSR[ 84 ][ 243 ],
   alphaCSR[ 84 ][ 244 ],
   alphaCSR[ 84 ][ 245 ],
   alphaCSR[ 84 ][ 246 ],
   alphaCSR[ 84 ][ 247 ],
   alphaCSR[ 84 ][ 248 ],
   alphaCSR[ 84 ][ 249 ],
   alphaCSR[ 84 ][ 250 ],
   alphaCSR[ 84 ][ 251 ],
   alphaCSR[ 84 ][ 252 ],
   alphaCSR[ 84 ][ 253 ],
   alphaCSR[ 84 ][ 254 ],
   alphaCSR[ 84 ][ 255 ],
   alphaCSR[ 84 ][ 256 ],
   alphaCSR[ 84 ][ 257 ],
   alphaCSR[ 84 ][ 258 ],
   alphaCSR[ 84 ][ 259 ],
   alphaCSR[ 84 ][ 260 ],
   alphaCSR[ 84 ][ 261 ],
   alphaCSR[ 84 ][ 262 ],
   alphaCSR[ 84 ][ 263 ],
   alphaCSR[ 84 ][ 264 ],
   alphaCSR[ 84 ][ 265 ],
   alphaCSR[ 84 ][ 266 ],
   alphaCSR[ 84 ][ 267 ],
   alphaCSR[ 84 ][ 268 ],
   alphaCSR[ 84 ][ 269 ],
   alphaCSR[ 84 ][ 270 ],
   alphaCSR[ 84 ][ 271 ],
   alphaCSR[ 84 ][ 272 ],
   alphaCSR[ 84 ][ 273 ],
   alphaCSR[ 84 ][ 274 ],
   alphaCSR[ 84 ][ 275 ],
   alphaCSR[ 84 ][ 276 ],
   alphaCSR[ 84 ][ 277 ],
   alphaCSR[ 84 ][ 278 ],
   alphaCSR[ 84 ][ 279 ],
   alphaCSR[ 84 ][ 280 ],
   alphaCSR[ 84 ][ 281 ],
   alphaCSR[ 84 ][ 282 ],
   alphaCSR[ 84 ][ 283 ],
   alphaCSR[ 84 ][ 284 ],
   alphaCSR[ 84 ][ 285 ],
   alphaCSR[ 84 ][ 286 ],
   alphaCSR[ 84 ][ 287 ],
   alphaCSR[ 84 ][ 288 ],
   alphaCSR[ 84 ][ 289 ],
   alphaCSR[ 84 ][ 290 ],
   alphaCSR[ 84 ][ 291 ],
   alphaCSR[ 84 ][ 292 ],
   alphaCSR[ 84 ][ 293 ],
   alphaCSR[ 84 ][ 294 ],
   alphaCSR[ 84 ][ 295 ],
   alphaCSR[ 84 ][ 296 ],
   alphaCSR[ 84 ][ 297 ],
   alphaCSR[ 84 ][ 298 ],
   alphaCSR[ 84 ][ 299 ],
   alphaCSR[ 84 ][ 300 ],
   alphaCSR[ 84 ][ 301 ],
   alphaCSR[ 84 ][ 302 ],
   alphaCSR[ 84 ][ 303 ],
   alphaCSR[ 84 ][ 304 ],
   alphaCSR[ 84 ][ 305 ],
   alphaCSR[ 84 ][ 306 ],
   alphaCSR[ 84 ][ 307 ],
   alphaCSR[ 84 ][ 308 ],
   alphaCSR[ 84 ][ 309 ],
   alphaCSR[ 84 ][ 310 ],
   alphaCSR[ 84 ][ 311 ],
   alphaCSR[ 84 ][ 312 ],
   alphaCSR[ 84 ][ 313 ],
   alphaCSR[ 84 ][ 314 ],
   alphaCSR[ 84 ][ 315 ],
   alphaCSR[ 84 ][ 316 ],
   alphaCSR[ 84 ][ 317 ],
   alphaCSR[ 84 ][ 318 ],
   alphaCSR[ 84 ][ 319 ],
   alphaCSR[ 84 ][ 320 ],
   alphaCSR[ 84 ][ 321 ],
   alphaCSR[ 84 ][ 322 ],
   alphaCSR[ 84 ][ 323 ],
   alphaCSR[ 84 ][ 324 ],
   alphaCSR[ 84 ][ 325 ],
   alphaCSR[ 84 ][ 326 ],
   alphaCSR[ 84 ][ 327 ],
   alphaCSR[ 84 ][ 328 ],
   alphaCSR[ 84 ][ 329 ],
   alphaCSR[ 84 ][ 330 ],
   alphaCSR[ 84 ][ 331 ],
   alphaCSR[ 84 ][ 332 ],
   alphaCSR[ 84 ][ 333 ],
   alphaCSR[ 84 ][ 334 ],
   alphaCSR[ 84 ][ 335 ],
   alphaCSR[ 84 ][ 336 ],
   alphaCSR[ 84 ][ 337 ],
   alphaCSR[ 84 ][ 338 ],
   alphaCSR[ 84 ][ 339 ],
   alphaCSR[ 84 ][ 340 ],
   alphaCSR[ 84 ][ 341 ],
   alphaCSR[ 84 ][ 342 ],
   alphaCSR[ 84 ][ 343 ],
   alphaCSR[ 84 ][ 344 ],
   alphaCSR[ 84 ][ 345 ],
   alphaCSR[ 84 ][ 346 ],
   alphaCSR[ 84 ][ 347 ],
   alphaCSR[ 84 ][ 348 ],
   alphaCSR[ 84 ][ 349 ],
   alphaCSR[ 84 ][ 350 ],
   alphaCSR[ 84 ][ 351 ],
   alphaCSR[ 84 ][ 352 ],
   alphaCSR[ 84 ][ 353 ],
   alphaCSR[ 84 ][ 354 ],
   alphaCSR[ 84 ][ 355 ],
   alphaCSR[ 84 ][ 356 ],
   alphaCSR[ 84 ][ 357 ],
   alphaCSR[ 84 ][ 358 ],
   alphaCSR[ 84 ][ 359 ],
   alphaCSR[ 84 ][ 360 ],
   alphaCSR[ 84 ][ 361 ],
   alphaCSR[ 84 ][ 362 ],
   alphaCSR[ 84 ][ 363 ],
   alphaCSR[ 84 ][ 364 ],
   alphaCSR[ 84 ][ 365 ],
   alphaCSR[ 84 ][ 366 ],
   alphaCSR[ 84 ][ 367 ],
   alphaCSR[ 84 ][ 368 ],
   alphaCSR[ 84 ][ 369 ],
   alphaCSR[ 84 ][ 370 ],
   alphaCSR[ 84 ][ 371 ],
   alphaCSR[ 84 ][ 372 ],
   alphaCSR[ 84 ][ 373 ],
   alphaCSR[ 84 ][ 374 ],
   alphaCSR[ 84 ][ 375 ],
   alphaCSR[ 84 ][ 376 ],
   alphaCSR[ 84 ][ 377 ],
   alphaCSR[ 84 ][ 378 ],
   alphaCSR[ 84 ][ 379 ],
   alphaCSR[ 84 ][ 380 ],
   alphaCSR[ 84 ][ 381 ],
   alphaCSR[ 84 ][ 382 ],
   alphaCSR[ 84 ][ 383 ],
   alphaCSR[ 85 ][ 0 ],
   alphaCSR[ 85 ][ 1 ],
   alphaCSR[ 85 ][ 2 ],
   alphaCSR[ 85 ][ 3 ],
   alphaCSR[ 85 ][ 4 ],
   alphaCSR[ 85 ][ 5 ],
   alphaCSR[ 85 ][ 6 ],
   alphaCSR[ 85 ][ 7 ],
   alphaCSR[ 85 ][ 8 ],
   alphaCSR[ 85 ][ 9 ],
   alphaCSR[ 85 ][ 10 ],
   alphaCSR[ 85 ][ 11 ],
   alphaCSR[ 85 ][ 12 ],
   alphaCSR[ 85 ][ 13 ],
   alphaCSR[ 85 ][ 14 ],
   alphaCSR[ 85 ][ 15 ],
   alphaCSR[ 85 ][ 16 ],
   alphaCSR[ 85 ][ 17 ],
   alphaCSR[ 85 ][ 18 ],
   alphaCSR[ 85 ][ 19 ],
   alphaCSR[ 85 ][ 20 ],
   alphaCSR[ 85 ][ 21 ],
   alphaCSR[ 85 ][ 22 ],
   alphaCSR[ 85 ][ 23 ],
   alphaCSR[ 85 ][ 24 ],
   alphaCSR[ 85 ][ 25 ],
   alphaCSR[ 85 ][ 26 ],
   alphaCSR[ 85 ][ 27 ],
   alphaCSR[ 85 ][ 28 ],
   alphaCSR[ 85 ][ 29 ],
   alphaCSR[ 85 ][ 30 ],
   alphaCSR[ 85 ][ 31 ],
   alphaCSR[ 85 ][ 32 ],
   alphaCSR[ 85 ][ 33 ],
   alphaCSR[ 85 ][ 34 ],
   alphaCSR[ 85 ][ 35 ],
   alphaCSR[ 85 ][ 36 ],
   alphaCSR[ 85 ][ 37 ],
   alphaCSR[ 85 ][ 38 ],
   alphaCSR[ 85 ][ 39 ],
   alphaCSR[ 85 ][ 40 ],
   alphaCSR[ 85 ][ 41 ],
   alphaCSR[ 85 ][ 42 ],
   alphaCSR[ 85 ][ 43 ],
   alphaCSR[ 85 ][ 44 ],
   alphaCSR[ 85 ][ 45 ],
   alphaCSR[ 85 ][ 46 ],
   alphaCSR[ 85 ][ 47 ],
   alphaCSR[ 85 ][ 48 ],
   alphaCSR[ 85 ][ 49 ],
   alphaCSR[ 85 ][ 50 ],
   alphaCSR[ 85 ][ 51 ],
   alphaCSR[ 85 ][ 52 ],
   alphaCSR[ 85 ][ 53 ],
   alphaCSR[ 85 ][ 54 ],
   alphaCSR[ 85 ][ 55 ],
   alphaCSR[ 85 ][ 56 ],
   alphaCSR[ 85 ][ 57 ],
   alphaCSR[ 85 ][ 58 ],
   alphaCSR[ 85 ][ 59 ],
   alphaCSR[ 85 ][ 60 ],
   alphaCSR[ 85 ][ 61 ],
   alphaCSR[ 85 ][ 62 ],
   alphaCSR[ 85 ][ 63 ],
   alphaCSR[ 85 ][ 64 ],
   alphaCSR[ 85 ][ 65 ],
   alphaCSR[ 85 ][ 66 ],
   alphaCSR[ 85 ][ 67 ],
   alphaCSR[ 85 ][ 68 ],
   alphaCSR[ 85 ][ 69 ],
   alphaCSR[ 85 ][ 70 ],
   alphaCSR[ 85 ][ 71 ],
   alphaCSR[ 85 ][ 72 ],
   alphaCSR[ 85 ][ 73 ],
   alphaCSR[ 85 ][ 74 ],
   alphaCSR[ 85 ][ 75 ],
   alphaCSR[ 85 ][ 76 ],
   alphaCSR[ 85 ][ 77 ],
   alphaCSR[ 85 ][ 78 ],
   alphaCSR[ 85 ][ 79 ],
   alphaCSR[ 85 ][ 80 ],
   alphaCSR[ 85 ][ 81 ],
   alphaCSR[ 85 ][ 82 ],
   alphaCSR[ 85 ][ 83 ],
   alphaCSR[ 85 ][ 84 ],
   alphaCSR[ 85 ][ 85 ],
   alphaCSR[ 85 ][ 86 ],
   alphaCSR[ 85 ][ 87 ],
   alphaCSR[ 85 ][ 88 ],
   alphaCSR[ 85 ][ 89 ],
   alphaCSR[ 85 ][ 90 ],
   alphaCSR[ 85 ][ 91 ],
   alphaCSR[ 85 ][ 92 ],
   alphaCSR[ 85 ][ 93 ],
   alphaCSR[ 85 ][ 94 ],
   alphaCSR[ 85 ][ 95 ],
   alphaCSR[ 85 ][ 96 ],
   alphaCSR[ 85 ][ 97 ],
   alphaCSR[ 85 ][ 98 ],
   alphaCSR[ 85 ][ 99 ],
   alphaCSR[ 85 ][ 100 ],
   alphaCSR[ 85 ][ 101 ],
   alphaCSR[ 85 ][ 102 ],
   alphaCSR[ 85 ][ 103 ],
   alphaCSR[ 85 ][ 104 ],
   alphaCSR[ 85 ][ 105 ],
   alphaCSR[ 85 ][ 106 ],
   alphaCSR[ 85 ][ 107 ],
   alphaCSR[ 85 ][ 108 ],
   alphaCSR[ 85 ][ 109 ],
   alphaCSR[ 85 ][ 110 ],
   alphaCSR[ 85 ][ 111 ],
   alphaCSR[ 85 ][ 112 ],
   alphaCSR[ 85 ][ 113 ],
   alphaCSR[ 85 ][ 114 ],
   alphaCSR[ 85 ][ 115 ],
   alphaCSR[ 85 ][ 116 ],
   alphaCSR[ 85 ][ 117 ],
   alphaCSR[ 85 ][ 118 ],
   alphaCSR[ 85 ][ 119 ],
   alphaCSR[ 85 ][ 120 ],
   alphaCSR[ 85 ][ 121 ],
   alphaCSR[ 85 ][ 122 ],
   alphaCSR[ 85 ][ 123 ],
   alphaCSR[ 85 ][ 124 ],
   alphaCSR[ 85 ][ 125 ],
   alphaCSR[ 85 ][ 126 ],
   alphaCSR[ 85 ][ 127 ],
   alphaCSR[ 85 ][ 128 ],
   alphaCSR[ 85 ][ 129 ],
   alphaCSR[ 85 ][ 130 ],
   alphaCSR[ 85 ][ 131 ],
   alphaCSR[ 85 ][ 132 ],
   alphaCSR[ 85 ][ 133 ],
   alphaCSR[ 85 ][ 134 ],
   alphaCSR[ 85 ][ 135 ],
   alphaCSR[ 85 ][ 136 ],
   alphaCSR[ 85 ][ 137 ],
   alphaCSR[ 85 ][ 138 ],
   alphaCSR[ 85 ][ 139 ],
   alphaCSR[ 85 ][ 140 ],
   alphaCSR[ 85 ][ 141 ],
   alphaCSR[ 85 ][ 142 ],
   alphaCSR[ 85 ][ 143 ],
   alphaCSR[ 85 ][ 144 ],
   alphaCSR[ 85 ][ 145 ],
   alphaCSR[ 85 ][ 146 ],
   alphaCSR[ 85 ][ 147 ],
   alphaCSR[ 85 ][ 148 ],
   alphaCSR[ 85 ][ 149 ],
   alphaCSR[ 85 ][ 150 ],
   alphaCSR[ 85 ][ 151 ],
   alphaCSR[ 85 ][ 152 ],
   alphaCSR[ 85 ][ 153 ],
   alphaCSR[ 85 ][ 154 ],
   alphaCSR[ 85 ][ 155 ],
   alphaCSR[ 85 ][ 156 ],
   alphaCSR[ 85 ][ 157 ],
   alphaCSR[ 85 ][ 158 ],
   alphaCSR[ 85 ][ 159 ],
   alphaCSR[ 85 ][ 160 ],
   alphaCSR[ 85 ][ 161 ],
   alphaCSR[ 85 ][ 162 ],
   alphaCSR[ 85 ][ 163 ],
   alphaCSR[ 85 ][ 164 ],
   alphaCSR[ 85 ][ 165 ],
   alphaCSR[ 85 ][ 166 ],
   alphaCSR[ 85 ][ 167 ],
   alphaCSR[ 85 ][ 168 ],
   alphaCSR[ 85 ][ 169 ],
   alphaCSR[ 85 ][ 170 ],
   alphaCSR[ 85 ][ 171 ],
   alphaCSR[ 85 ][ 172 ],
   alphaCSR[ 85 ][ 173 ],
   alphaCSR[ 85 ][ 174 ],
   alphaCSR[ 85 ][ 175 ],
   alphaCSR[ 85 ][ 176 ],
   alphaCSR[ 85 ][ 177 ],
   alphaCSR[ 85 ][ 178 ],
   alphaCSR[ 85 ][ 179 ],
   alphaCSR[ 85 ][ 180 ],
   alphaCSR[ 85 ][ 181 ],
   alphaCSR[ 85 ][ 182 ],
   alphaCSR[ 85 ][ 183 ],
   alphaCSR[ 85 ][ 184 ],
   alphaCSR[ 85 ][ 185 ],
   alphaCSR[ 85 ][ 186 ],
   alphaCSR[ 85 ][ 187 ],
   alphaCSR[ 85 ][ 188 ],
   alphaCSR[ 85 ][ 189 ],
   alphaCSR[ 85 ][ 190 ],
   alphaCSR[ 85 ][ 191 ],
   alphaCSR[ 85 ][ 192 ],
   alphaCSR[ 85 ][ 193 ],
   alphaCSR[ 85 ][ 194 ],
   alphaCSR[ 85 ][ 195 ],
   alphaCSR[ 85 ][ 196 ],
   alphaCSR[ 85 ][ 197 ],
   alphaCSR[ 85 ][ 198 ],
   alphaCSR[ 85 ][ 199 ],
   alphaCSR[ 85 ][ 200 ],
   alphaCSR[ 85 ][ 201 ],
   alphaCSR[ 85 ][ 202 ],
   alphaCSR[ 85 ][ 203 ],
   alphaCSR[ 85 ][ 204 ],
   alphaCSR[ 85 ][ 205 ],
   alphaCSR[ 85 ][ 206 ],
   alphaCSR[ 85 ][ 207 ],
   alphaCSR[ 85 ][ 208 ],
   alphaCSR[ 85 ][ 209 ],
   alphaCSR[ 85 ][ 210 ],
   alphaCSR[ 85 ][ 211 ],
   alphaCSR[ 85 ][ 212 ],
   alphaCSR[ 85 ][ 213 ],
   alphaCSR[ 85 ][ 214 ],
   alphaCSR[ 85 ][ 215 ],
   alphaCSR[ 85 ][ 216 ],
   alphaCSR[ 85 ][ 217 ],
   alphaCSR[ 85 ][ 218 ],
   alphaCSR[ 85 ][ 219 ],
   alphaCSR[ 85 ][ 220 ],
   alphaCSR[ 85 ][ 221 ],
   alphaCSR[ 85 ][ 222 ],
   alphaCSR[ 85 ][ 223 ],
   alphaCSR[ 85 ][ 224 ],
   alphaCSR[ 85 ][ 225 ],
   alphaCSR[ 85 ][ 226 ],
   alphaCSR[ 85 ][ 227 ],
   alphaCSR[ 85 ][ 228 ],
   alphaCSR[ 85 ][ 229 ],
   alphaCSR[ 85 ][ 230 ],
   alphaCSR[ 85 ][ 231 ],
   alphaCSR[ 85 ][ 232 ],
   alphaCSR[ 85 ][ 233 ],
   alphaCSR[ 85 ][ 234 ],
   alphaCSR[ 85 ][ 235 ],
   alphaCSR[ 85 ][ 236 ],
   alphaCSR[ 85 ][ 237 ],
   alphaCSR[ 85 ][ 238 ],
   alphaCSR[ 85 ][ 239 ],
   alphaCSR[ 85 ][ 240 ],
   alphaCSR[ 85 ][ 241 ],
   alphaCSR[ 85 ][ 242 ],
   alphaCSR[ 85 ][ 243 ],
   alphaCSR[ 85 ][ 244 ],
   alphaCSR[ 85 ][ 245 ],
   alphaCSR[ 85 ][ 246 ],
   alphaCSR[ 85 ][ 247 ],
   alphaCSR[ 85 ][ 248 ],
   alphaCSR[ 85 ][ 249 ],
   alphaCSR[ 85 ][ 250 ],
   alphaCSR[ 85 ][ 251 ],
   alphaCSR[ 85 ][ 252 ],
   alphaCSR[ 85 ][ 253 ],
   alphaCSR[ 85 ][ 254 ],
   alphaCSR[ 85 ][ 255 ],
   alphaCSR[ 85 ][ 256 ],
   alphaCSR[ 85 ][ 257 ],
   alphaCSR[ 85 ][ 258 ],
   alphaCSR[ 85 ][ 259 ],
   alphaCSR[ 85 ][ 260 ],
   alphaCSR[ 85 ][ 261 ],
   alphaCSR[ 85 ][ 262 ],
   alphaCSR[ 85 ][ 263 ],
   alphaCSR[ 85 ][ 264 ],
   alphaCSR[ 85 ][ 265 ],
   alphaCSR[ 85 ][ 266 ],
   alphaCSR[ 85 ][ 267 ],
   alphaCSR[ 85 ][ 268 ],
   alphaCSR[ 85 ][ 269 ],
   alphaCSR[ 85 ][ 270 ],
   alphaCSR[ 85 ][ 271 ],
   alphaCSR[ 85 ][ 272 ],
   alphaCSR[ 85 ][ 273 ],
   alphaCSR[ 85 ][ 274 ],
   alphaCSR[ 85 ][ 275 ],
   alphaCSR[ 85 ][ 276 ],
   alphaCSR[ 85 ][ 277 ],
   alphaCSR[ 85 ][ 278 ],
   alphaCSR[ 85 ][ 279 ],
   alphaCSR[ 85 ][ 280 ],
   alphaCSR[ 85 ][ 281 ],
   alphaCSR[ 85 ][ 282 ],
   alphaCSR[ 85 ][ 283 ],
   alphaCSR[ 85 ][ 284 ],
   alphaCSR[ 85 ][ 285 ],
   alphaCSR[ 85 ][ 286 ],
   alphaCSR[ 85 ][ 287 ],
   alphaCSR[ 85 ][ 288 ],
   alphaCSR[ 85 ][ 289 ],
   alphaCSR[ 85 ][ 290 ],
   alphaCSR[ 85 ][ 291 ],
   alphaCSR[ 85 ][ 292 ],
   alphaCSR[ 85 ][ 293 ],
   alphaCSR[ 85 ][ 294 ],
   alphaCSR[ 85 ][ 295 ],
   alphaCSR[ 85 ][ 296 ],
   alphaCSR[ 85 ][ 297 ],
   alphaCSR[ 85 ][ 298 ],
   alphaCSR[ 85 ][ 299 ],
   alphaCSR[ 85 ][ 300 ],
   alphaCSR[ 85 ][ 301 ],
   alphaCSR[ 85 ][ 302 ],
   alphaCSR[ 85 ][ 303 ],
   alphaCSR[ 85 ][ 304 ],
   alphaCSR[ 85 ][ 305 ],
   alphaCSR[ 85 ][ 306 ],
   alphaCSR[ 85 ][ 307 ],
   alphaCSR[ 85 ][ 308 ],
   alphaCSR[ 85 ][ 309 ],
   alphaCSR[ 85 ][ 310 ],
   alphaCSR[ 85 ][ 311 ],
   alphaCSR[ 85 ][ 312 ],
   alphaCSR[ 85 ][ 313 ],
   alphaCSR[ 85 ][ 314 ],
   alphaCSR[ 85 ][ 315 ],
   alphaCSR[ 85 ][ 316 ],
   alphaCSR[ 85 ][ 317 ],
   alphaCSR[ 85 ][ 318 ],
   alphaCSR[ 85 ][ 319 ],
   alphaCSR[ 85 ][ 320 ],
   alphaCSR[ 85 ][ 321 ],
   alphaCSR[ 85 ][ 322 ],
   alphaCSR[ 85 ][ 323 ],
   alphaCSR[ 85 ][ 324 ],
   alphaCSR[ 85 ][ 325 ],
   alphaCSR[ 85 ][ 326 ],
   alphaCSR[ 85 ][ 327 ],
   alphaCSR[ 85 ][ 328 ],
   alphaCSR[ 85 ][ 329 ],
   alphaCSR[ 85 ][ 330 ],
   alphaCSR[ 85 ][ 331 ],
   alphaCSR[ 85 ][ 332 ],
   alphaCSR[ 85 ][ 333 ],
   alphaCSR[ 85 ][ 334 ],
   alphaCSR[ 85 ][ 335 ],
   alphaCSR[ 85 ][ 336 ],
   alphaCSR[ 85 ][ 337 ],
   alphaCSR[ 85 ][ 338 ],
   alphaCSR[ 85 ][ 339 ],
   alphaCSR[ 85 ][ 340 ],
   alphaCSR[ 85 ][ 341 ],
   alphaCSR[ 85 ][ 342 ],
   alphaCSR[ 85 ][ 343 ],
   alphaCSR[ 85 ][ 344 ],
   alphaCSR[ 85 ][ 345 ],
   alphaCSR[ 85 ][ 346 ],
   alphaCSR[ 85 ][ 347 ],
   alphaCSR[ 85 ][ 348 ],
   alphaCSR[ 85 ][ 349 ],
   alphaCSR[ 85 ][ 350 ],
   alphaCSR[ 85 ][ 351 ],
   alphaCSR[ 85 ][ 352 ],
   alphaCSR[ 85 ][ 353 ],
   alphaCSR[ 85 ][ 354 ],
   alphaCSR[ 85 ][ 355 ],
   alphaCSR[ 85 ][ 356 ],
   alphaCSR[ 85 ][ 357 ],
   alphaCSR[ 85 ][ 358 ],
   alphaCSR[ 85 ][ 359 ],
   alphaCSR[ 85 ][ 360 ],
   alphaCSR[ 85 ][ 361 ],
   alphaCSR[ 85 ][ 362 ],
   alphaCSR[ 85 ][ 363 ],
   alphaCSR[ 85 ][ 364 ],
   alphaCSR[ 85 ][ 365 ],
   alphaCSR[ 85 ][ 366 ],
   alphaCSR[ 85 ][ 367 ],
   alphaCSR[ 85 ][ 368 ],
   alphaCSR[ 85 ][ 369 ],
   alphaCSR[ 85 ][ 370 ],
   alphaCSR[ 85 ][ 371 ],
   alphaCSR[ 85 ][ 372 ],
   alphaCSR[ 85 ][ 373 ],
   alphaCSR[ 85 ][ 374 ],
   alphaCSR[ 85 ][ 375 ],
   alphaCSR[ 85 ][ 376 ],
   alphaCSR[ 85 ][ 377 ],
   alphaCSR[ 85 ][ 378 ],
   alphaCSR[ 85 ][ 379 ],
   alphaCSR[ 85 ][ 380 ],
   alphaCSR[ 85 ][ 381 ],
   alphaCSR[ 85 ][ 382 ],
   alphaCSR[ 85 ][ 383 ],
   alphaCSR[ 86 ][ 0 ],
   alphaCSR[ 86 ][ 1 ],
   alphaCSR[ 86 ][ 2 ],
   alphaCSR[ 86 ][ 3 ],
   alphaCSR[ 86 ][ 4 ],
   alphaCSR[ 86 ][ 5 ],
   alphaCSR[ 86 ][ 6 ],
   alphaCSR[ 86 ][ 7 ],
   alphaCSR[ 86 ][ 8 ],
   alphaCSR[ 86 ][ 9 ],
   alphaCSR[ 86 ][ 10 ],
   alphaCSR[ 86 ][ 11 ],
   alphaCSR[ 86 ][ 12 ],
   alphaCSR[ 86 ][ 13 ],
   alphaCSR[ 86 ][ 14 ],
   alphaCSR[ 86 ][ 15 ],
   alphaCSR[ 86 ][ 16 ],
   alphaCSR[ 86 ][ 17 ],
   alphaCSR[ 86 ][ 18 ],
   alphaCSR[ 86 ][ 19 ],
   alphaCSR[ 86 ][ 20 ],
   alphaCSR[ 86 ][ 21 ],
   alphaCSR[ 86 ][ 22 ],
   alphaCSR[ 86 ][ 23 ],
   alphaCSR[ 86 ][ 24 ],
   alphaCSR[ 86 ][ 25 ],
   alphaCSR[ 86 ][ 26 ],
   alphaCSR[ 86 ][ 27 ],
   alphaCSR[ 86 ][ 28 ],
   alphaCSR[ 86 ][ 29 ],
   alphaCSR[ 86 ][ 30 ],
   alphaCSR[ 86 ][ 31 ],
   alphaCSR[ 86 ][ 32 ],
   alphaCSR[ 86 ][ 33 ],
   alphaCSR[ 86 ][ 34 ],
   alphaCSR[ 86 ][ 35 ],
   alphaCSR[ 86 ][ 36 ],
   alphaCSR[ 86 ][ 37 ],
   alphaCSR[ 86 ][ 38 ],
   alphaCSR[ 86 ][ 39 ],
   alphaCSR[ 86 ][ 40 ],
   alphaCSR[ 86 ][ 41 ],
   alphaCSR[ 86 ][ 42 ],
   alphaCSR[ 86 ][ 43 ],
   alphaCSR[ 86 ][ 44 ],
   alphaCSR[ 86 ][ 45 ],
   alphaCSR[ 86 ][ 46 ],
   alphaCSR[ 86 ][ 47 ],
   alphaCSR[ 86 ][ 48 ],
   alphaCSR[ 86 ][ 49 ],
   alphaCSR[ 86 ][ 50 ],
   alphaCSR[ 86 ][ 51 ],
   alphaCSR[ 86 ][ 52 ],
   alphaCSR[ 86 ][ 53 ],
   alphaCSR[ 86 ][ 54 ],
   alphaCSR[ 86 ][ 55 ],
   alphaCSR[ 86 ][ 56 ],
   alphaCSR[ 86 ][ 57 ],
   alphaCSR[ 86 ][ 58 ],
   alphaCSR[ 86 ][ 59 ],
   alphaCSR[ 86 ][ 60 ],
   alphaCSR[ 86 ][ 61 ],
   alphaCSR[ 86 ][ 62 ],
   alphaCSR[ 86 ][ 63 ],
   alphaCSR[ 86 ][ 64 ],
   alphaCSR[ 86 ][ 65 ],
   alphaCSR[ 86 ][ 66 ],
   alphaCSR[ 86 ][ 67 ],
   alphaCSR[ 86 ][ 68 ],
   alphaCSR[ 86 ][ 69 ],
   alphaCSR[ 86 ][ 70 ],
   alphaCSR[ 86 ][ 71 ],
   alphaCSR[ 86 ][ 72 ],
   alphaCSR[ 86 ][ 73 ],
   alphaCSR[ 86 ][ 74 ],
   alphaCSR[ 86 ][ 75 ],
   alphaCSR[ 86 ][ 76 ],
   alphaCSR[ 86 ][ 77 ],
   alphaCSR[ 86 ][ 78 ],
   alphaCSR[ 86 ][ 79 ],
   alphaCSR[ 86 ][ 80 ],
   alphaCSR[ 86 ][ 81 ],
   alphaCSR[ 86 ][ 82 ],
   alphaCSR[ 86 ][ 83 ],
   alphaCSR[ 86 ][ 84 ],
   alphaCSR[ 86 ][ 85 ],
   alphaCSR[ 86 ][ 86 ],
   alphaCSR[ 86 ][ 87 ],
   alphaCSR[ 86 ][ 88 ],
   alphaCSR[ 86 ][ 89 ],
   alphaCSR[ 86 ][ 90 ],
   alphaCSR[ 86 ][ 91 ],
   alphaCSR[ 86 ][ 92 ],
   alphaCSR[ 86 ][ 93 ],
   alphaCSR[ 86 ][ 94 ],
   alphaCSR[ 86 ][ 95 ],
   alphaCSR[ 86 ][ 96 ],
   alphaCSR[ 86 ][ 97 ],
   alphaCSR[ 86 ][ 98 ],
   alphaCSR[ 86 ][ 99 ],
   alphaCSR[ 86 ][ 100 ],
   alphaCSR[ 86 ][ 101 ],
   alphaCSR[ 86 ][ 102 ],
   alphaCSR[ 86 ][ 103 ],
   alphaCSR[ 86 ][ 104 ],
   alphaCSR[ 86 ][ 105 ],
   alphaCSR[ 86 ][ 106 ],
   alphaCSR[ 86 ][ 107 ],
   alphaCSR[ 86 ][ 108 ],
   alphaCSR[ 86 ][ 109 ],
   alphaCSR[ 86 ][ 110 ],
   alphaCSR[ 86 ][ 111 ],
   alphaCSR[ 86 ][ 112 ],
   alphaCSR[ 86 ][ 113 ],
   alphaCSR[ 86 ][ 114 ],
   alphaCSR[ 86 ][ 115 ],
   alphaCSR[ 86 ][ 116 ],
   alphaCSR[ 86 ][ 117 ],
   alphaCSR[ 86 ][ 118 ],
   alphaCSR[ 86 ][ 119 ],
   alphaCSR[ 86 ][ 120 ],
   alphaCSR[ 86 ][ 121 ],
   alphaCSR[ 86 ][ 122 ],
   alphaCSR[ 86 ][ 123 ],
   alphaCSR[ 86 ][ 124 ],
   alphaCSR[ 86 ][ 125 ],
   alphaCSR[ 86 ][ 126 ],
   alphaCSR[ 86 ][ 127 ],
   alphaCSR[ 86 ][ 128 ],
   alphaCSR[ 86 ][ 129 ],
   alphaCSR[ 86 ][ 130 ],
   alphaCSR[ 86 ][ 131 ],
   alphaCSR[ 86 ][ 132 ],
   alphaCSR[ 86 ][ 133 ],
   alphaCSR[ 86 ][ 134 ],
   alphaCSR[ 86 ][ 135 ],
   alphaCSR[ 86 ][ 136 ],
   alphaCSR[ 86 ][ 137 ],
   alphaCSR[ 86 ][ 138 ],
   alphaCSR[ 86 ][ 139 ],
   alphaCSR[ 86 ][ 140 ],
   alphaCSR[ 86 ][ 141 ],
   alphaCSR[ 86 ][ 142 ],
   alphaCSR[ 86 ][ 143 ],
   alphaCSR[ 86 ][ 144 ],
   alphaCSR[ 86 ][ 145 ],
   alphaCSR[ 86 ][ 146 ],
   alphaCSR[ 86 ][ 147 ],
   alphaCSR[ 86 ][ 148 ],
   alphaCSR[ 86 ][ 149 ],
   alphaCSR[ 86 ][ 150 ],
   alphaCSR[ 86 ][ 151 ],
   alphaCSR[ 86 ][ 152 ],
   alphaCSR[ 86 ][ 153 ],
   alphaCSR[ 86 ][ 154 ],
   alphaCSR[ 86 ][ 155 ],
   alphaCSR[ 86 ][ 156 ],
   alphaCSR[ 86 ][ 157 ],
   alphaCSR[ 86 ][ 158 ],
   alphaCSR[ 86 ][ 159 ],
   alphaCSR[ 86 ][ 160 ],
   alphaCSR[ 86 ][ 161 ],
   alphaCSR[ 86 ][ 162 ],
   alphaCSR[ 86 ][ 163 ],
   alphaCSR[ 86 ][ 164 ],
   alphaCSR[ 86 ][ 165 ],
   alphaCSR[ 86 ][ 166 ],
   alphaCSR[ 86 ][ 167 ],
   alphaCSR[ 86 ][ 168 ],
   alphaCSR[ 86 ][ 169 ],
   alphaCSR[ 86 ][ 170 ],
   alphaCSR[ 86 ][ 171 ],
   alphaCSR[ 86 ][ 172 ],
   alphaCSR[ 86 ][ 173 ],
   alphaCSR[ 86 ][ 174 ],
   alphaCSR[ 86 ][ 175 ],
   alphaCSR[ 86 ][ 176 ],
   alphaCSR[ 86 ][ 177 ],
   alphaCSR[ 86 ][ 178 ],
   alphaCSR[ 86 ][ 179 ],
   alphaCSR[ 86 ][ 180 ],
   alphaCSR[ 86 ][ 181 ],
   alphaCSR[ 86 ][ 182 ],
   alphaCSR[ 86 ][ 183 ],
   alphaCSR[ 86 ][ 184 ],
   alphaCSR[ 86 ][ 185 ],
   alphaCSR[ 86 ][ 186 ],
   alphaCSR[ 86 ][ 187 ],
   alphaCSR[ 86 ][ 188 ],
   alphaCSR[ 86 ][ 189 ],
   alphaCSR[ 86 ][ 190 ],
   alphaCSR[ 86 ][ 191 ],
   alphaCSR[ 86 ][ 192 ],
   alphaCSR[ 86 ][ 193 ],
   alphaCSR[ 86 ][ 194 ],
   alphaCSR[ 86 ][ 195 ],
   alphaCSR[ 86 ][ 196 ],
   alphaCSR[ 86 ][ 197 ],
   alphaCSR[ 86 ][ 198 ],
   alphaCSR[ 86 ][ 199 ],
   alphaCSR[ 86 ][ 200 ],
   alphaCSR[ 86 ][ 201 ],
   alphaCSR[ 86 ][ 202 ],
   alphaCSR[ 86 ][ 203 ],
   alphaCSR[ 86 ][ 204 ],
   alphaCSR[ 86 ][ 205 ],
   alphaCSR[ 86 ][ 206 ],
   alphaCSR[ 86 ][ 207 ],
   alphaCSR[ 86 ][ 208 ],
   alphaCSR[ 86 ][ 209 ],
   alphaCSR[ 86 ][ 210 ],
   alphaCSR[ 86 ][ 211 ],
   alphaCSR[ 86 ][ 212 ],
   alphaCSR[ 86 ][ 213 ],
   alphaCSR[ 86 ][ 214 ],
   alphaCSR[ 86 ][ 215 ],
   alphaCSR[ 86 ][ 216 ],
   alphaCSR[ 86 ][ 217 ],
   alphaCSR[ 86 ][ 218 ],
   alphaCSR[ 86 ][ 219 ],
   alphaCSR[ 86 ][ 220 ],
   alphaCSR[ 86 ][ 221 ],
   alphaCSR[ 86 ][ 222 ],
   alphaCSR[ 86 ][ 223 ],
   alphaCSR[ 86 ][ 224 ],
   alphaCSR[ 86 ][ 225 ],
   alphaCSR[ 86 ][ 226 ],
   alphaCSR[ 86 ][ 227 ],
   alphaCSR[ 86 ][ 228 ],
   alphaCSR[ 86 ][ 229 ],
   alphaCSR[ 86 ][ 230 ],
   alphaCSR[ 86 ][ 231 ],
   alphaCSR[ 86 ][ 232 ],
   alphaCSR[ 86 ][ 233 ],
   alphaCSR[ 86 ][ 234 ],
   alphaCSR[ 86 ][ 235 ],
   alphaCSR[ 86 ][ 236 ],
   alphaCSR[ 86 ][ 237 ],
   alphaCSR[ 86 ][ 238 ],
   alphaCSR[ 86 ][ 239 ],
   alphaCSR[ 86 ][ 240 ],
   alphaCSR[ 86 ][ 241 ],
   alphaCSR[ 86 ][ 242 ],
   alphaCSR[ 86 ][ 243 ],
   alphaCSR[ 86 ][ 244 ],
   alphaCSR[ 86 ][ 245 ],
   alphaCSR[ 86 ][ 246 ],
   alphaCSR[ 86 ][ 247 ],
   alphaCSR[ 86 ][ 248 ],
   alphaCSR[ 86 ][ 249 ],
   alphaCSR[ 86 ][ 250 ],
   alphaCSR[ 86 ][ 251 ],
   alphaCSR[ 86 ][ 252 ],
   alphaCSR[ 86 ][ 253 ],
   alphaCSR[ 86 ][ 254 ],
   alphaCSR[ 86 ][ 255 ],
   alphaCSR[ 86 ][ 256 ],
   alphaCSR[ 86 ][ 257 ],
   alphaCSR[ 86 ][ 258 ],
   alphaCSR[ 86 ][ 259 ],
   alphaCSR[ 86 ][ 260 ],
   alphaCSR[ 86 ][ 261 ],
   alphaCSR[ 86 ][ 262 ],
   alphaCSR[ 86 ][ 263 ],
   alphaCSR[ 86 ][ 264 ],
   alphaCSR[ 86 ][ 265 ],
   alphaCSR[ 86 ][ 266 ],
   alphaCSR[ 86 ][ 267 ],
   alphaCSR[ 86 ][ 268 ],
   alphaCSR[ 86 ][ 269 ],
   alphaCSR[ 86 ][ 270 ],
   alphaCSR[ 86 ][ 271 ],
   alphaCSR[ 86 ][ 272 ],
   alphaCSR[ 86 ][ 273 ],
   alphaCSR[ 86 ][ 274 ],
   alphaCSR[ 86 ][ 275 ],
   alphaCSR[ 86 ][ 276 ],
   alphaCSR[ 86 ][ 277 ],
   alphaCSR[ 86 ][ 278 ],
   alphaCSR[ 86 ][ 279 ],
   alphaCSR[ 86 ][ 280 ],
   alphaCSR[ 86 ][ 281 ],
   alphaCSR[ 86 ][ 282 ],
   alphaCSR[ 86 ][ 283 ],
   alphaCSR[ 86 ][ 284 ],
   alphaCSR[ 86 ][ 285 ],
   alphaCSR[ 86 ][ 286 ],
   alphaCSR[ 86 ][ 287 ],
   alphaCSR[ 86 ][ 288 ],
   alphaCSR[ 86 ][ 289 ],
   alphaCSR[ 86 ][ 290 ],
   alphaCSR[ 86 ][ 291 ],
   alphaCSR[ 86 ][ 292 ],
   alphaCSR[ 86 ][ 293 ],
   alphaCSR[ 86 ][ 294 ],
   alphaCSR[ 86 ][ 295 ],
   alphaCSR[ 86 ][ 296 ],
   alphaCSR[ 86 ][ 297 ],
   alphaCSR[ 86 ][ 298 ],
   alphaCSR[ 86 ][ 299 ],
   alphaCSR[ 86 ][ 300 ],
   alphaCSR[ 86 ][ 301 ],
   alphaCSR[ 86 ][ 302 ],
   alphaCSR[ 86 ][ 303 ],
   alphaCSR[ 86 ][ 304 ],
   alphaCSR[ 86 ][ 305 ],
   alphaCSR[ 86 ][ 306 ],
   alphaCSR[ 86 ][ 307 ],
   alphaCSR[ 86 ][ 308 ],
   alphaCSR[ 86 ][ 309 ],
   alphaCSR[ 86 ][ 310 ],
   alphaCSR[ 86 ][ 311 ],
   alphaCSR[ 86 ][ 312 ],
   alphaCSR[ 86 ][ 313 ],
   alphaCSR[ 86 ][ 314 ],
   alphaCSR[ 86 ][ 315 ],
   alphaCSR[ 86 ][ 316 ],
   alphaCSR[ 86 ][ 317 ],
   alphaCSR[ 86 ][ 318 ],
   alphaCSR[ 86 ][ 319 ],
   alphaCSR[ 86 ][ 320 ],
   alphaCSR[ 86 ][ 321 ],
   alphaCSR[ 86 ][ 322 ],
   alphaCSR[ 86 ][ 323 ],
   alphaCSR[ 86 ][ 324 ],
   alphaCSR[ 86 ][ 325 ],
   alphaCSR[ 86 ][ 326 ],
   alphaCSR[ 86 ][ 327 ],
   alphaCSR[ 86 ][ 328 ],
   alphaCSR[ 86 ][ 329 ],
   alphaCSR[ 86 ][ 330 ],
   alphaCSR[ 86 ][ 331 ],
   alphaCSR[ 86 ][ 332 ],
   alphaCSR[ 86 ][ 333 ],
   alphaCSR[ 86 ][ 334 ],
   alphaCSR[ 86 ][ 335 ],
   alphaCSR[ 86 ][ 336 ],
   alphaCSR[ 86 ][ 337 ],
   alphaCSR[ 86 ][ 338 ],
   alphaCSR[ 86 ][ 339 ],
   alphaCSR[ 86 ][ 340 ],
   alphaCSR[ 86 ][ 341 ],
   alphaCSR[ 86 ][ 342 ],
   alphaCSR[ 86 ][ 343 ],
   alphaCSR[ 86 ][ 344 ],
   alphaCSR[ 86 ][ 345 ],
   alphaCSR[ 86 ][ 346 ],
   alphaCSR[ 86 ][ 347 ],
   alphaCSR[ 86 ][ 348 ],
   alphaCSR[ 86 ][ 349 ],
   alphaCSR[ 86 ][ 350 ],
   alphaCSR[ 86 ][ 351 ],
   alphaCSR[ 86 ][ 352 ],
   alphaCSR[ 86 ][ 353 ],
   alphaCSR[ 86 ][ 354 ],
   alphaCSR[ 86 ][ 355 ],
   alphaCSR[ 86 ][ 356 ],
   alphaCSR[ 86 ][ 357 ],
   alphaCSR[ 86 ][ 358 ],
   alphaCSR[ 86 ][ 359 ],
   alphaCSR[ 86 ][ 360 ],
   alphaCSR[ 86 ][ 361 ],
   alphaCSR[ 86 ][ 362 ],
   alphaCSR[ 86 ][ 363 ],
   alphaCSR[ 86 ][ 364 ],
   alphaCSR[ 86 ][ 365 ],
   alphaCSR[ 86 ][ 366 ],
   alphaCSR[ 86 ][ 367 ],
   alphaCSR[ 86 ][ 368 ],
   alphaCSR[ 86 ][ 369 ],
   alphaCSR[ 86 ][ 370 ],
   alphaCSR[ 86 ][ 371 ],
   alphaCSR[ 86 ][ 372 ],
   alphaCSR[ 86 ][ 373 ],
   alphaCSR[ 86 ][ 374 ],
   alphaCSR[ 86 ][ 375 ],
   alphaCSR[ 86 ][ 376 ],
   alphaCSR[ 86 ][ 377 ],
   alphaCSR[ 86 ][ 378 ],
   alphaCSR[ 86 ][ 379 ],
   alphaCSR[ 86 ][ 380 ],
   alphaCSR[ 86 ][ 381 ],
   alphaCSR[ 86 ][ 382 ],
   alphaCSR[ 86 ][ 383 ],
   alphaCSR[ 87 ][ 0 ],
   alphaCSR[ 87 ][ 1 ],
   alphaCSR[ 87 ][ 2 ],
   alphaCSR[ 87 ][ 3 ],
   alphaCSR[ 87 ][ 4 ],
   alphaCSR[ 87 ][ 5 ],
   alphaCSR[ 87 ][ 6 ],
   alphaCSR[ 87 ][ 7 ],
   alphaCSR[ 87 ][ 8 ],
   alphaCSR[ 87 ][ 9 ],
   alphaCSR[ 87 ][ 10 ],
   alphaCSR[ 87 ][ 11 ],
   alphaCSR[ 87 ][ 12 ],
   alphaCSR[ 87 ][ 13 ],
   alphaCSR[ 87 ][ 14 ],
   alphaCSR[ 87 ][ 15 ],
   alphaCSR[ 87 ][ 16 ],
   alphaCSR[ 87 ][ 17 ],
   alphaCSR[ 87 ][ 18 ],
   alphaCSR[ 87 ][ 19 ],
   alphaCSR[ 87 ][ 20 ],
   alphaCSR[ 87 ][ 21 ],
   alphaCSR[ 87 ][ 22 ],
   alphaCSR[ 87 ][ 23 ],
   alphaCSR[ 87 ][ 24 ],
   alphaCSR[ 87 ][ 25 ],
   alphaCSR[ 87 ][ 26 ],
   alphaCSR[ 87 ][ 27 ],
   alphaCSR[ 87 ][ 28 ],
   alphaCSR[ 87 ][ 29 ],
   alphaCSR[ 87 ][ 30 ],
   alphaCSR[ 87 ][ 31 ],
   alphaCSR[ 87 ][ 32 ],
   alphaCSR[ 87 ][ 33 ],
   alphaCSR[ 87 ][ 34 ],
   alphaCSR[ 87 ][ 35 ],
   alphaCSR[ 87 ][ 36 ],
   alphaCSR[ 87 ][ 37 ],
   alphaCSR[ 87 ][ 38 ],
   alphaCSR[ 87 ][ 39 ],
   alphaCSR[ 87 ][ 40 ],
   alphaCSR[ 87 ][ 41 ],
   alphaCSR[ 87 ][ 42 ],
   alphaCSR[ 87 ][ 43 ],
   alphaCSR[ 87 ][ 44 ],
   alphaCSR[ 87 ][ 45 ],
   alphaCSR[ 87 ][ 46 ],
   alphaCSR[ 87 ][ 47 ],
   alphaCSR[ 87 ][ 48 ],
   alphaCSR[ 87 ][ 49 ],
   alphaCSR[ 87 ][ 50 ],
   alphaCSR[ 87 ][ 51 ],
   alphaCSR[ 87 ][ 52 ],
   alphaCSR[ 87 ][ 53 ],
   alphaCSR[ 87 ][ 54 ],
   alphaCSR[ 87 ][ 55 ],
   alphaCSR[ 87 ][ 56 ],
   alphaCSR[ 87 ][ 57 ],
   alphaCSR[ 87 ][ 58 ],
   alphaCSR[ 87 ][ 59 ],
   alphaCSR[ 87 ][ 60 ],
   alphaCSR[ 87 ][ 61 ],
   alphaCSR[ 87 ][ 62 ],
   alphaCSR[ 87 ][ 63 ],
   alphaCSR[ 87 ][ 64 ],
   alphaCSR[ 87 ][ 65 ],
   alphaCSR[ 87 ][ 66 ],
   alphaCSR[ 87 ][ 67 ],
   alphaCSR[ 87 ][ 68 ],
   alphaCSR[ 87 ][ 69 ],
   alphaCSR[ 87 ][ 70 ],
   alphaCSR[ 87 ][ 71 ],
   alphaCSR[ 87 ][ 72 ],
   alphaCSR[ 87 ][ 73 ],
   alphaCSR[ 87 ][ 74 ],
   alphaCSR[ 87 ][ 75 ],
   alphaCSR[ 87 ][ 76 ],
   alphaCSR[ 87 ][ 77 ],
   alphaCSR[ 87 ][ 78 ],
   alphaCSR[ 87 ][ 79 ],
   alphaCSR[ 87 ][ 80 ],
   alphaCSR[ 87 ][ 81 ],
   alphaCSR[ 87 ][ 82 ],
   alphaCSR[ 87 ][ 83 ],
   alphaCSR[ 87 ][ 84 ],
   alphaCSR[ 87 ][ 85 ],
   alphaCSR[ 87 ][ 86 ],
   alphaCSR[ 87 ][ 87 ],
   alphaCSR[ 87 ][ 88 ],
   alphaCSR[ 87 ][ 89 ],
   alphaCSR[ 87 ][ 90 ],
   alphaCSR[ 87 ][ 91 ],
   alphaCSR[ 87 ][ 92 ],
   alphaCSR[ 87 ][ 93 ],
   alphaCSR[ 87 ][ 94 ],
   alphaCSR[ 87 ][ 95 ],
   alphaCSR[ 87 ][ 96 ],
   alphaCSR[ 87 ][ 97 ],
   alphaCSR[ 87 ][ 98 ],
   alphaCSR[ 87 ][ 99 ],
   alphaCSR[ 87 ][ 100 ],
   alphaCSR[ 87 ][ 101 ],
   alphaCSR[ 87 ][ 102 ],
   alphaCSR[ 87 ][ 103 ],
   alphaCSR[ 87 ][ 104 ],
   alphaCSR[ 87 ][ 105 ],
   alphaCSR[ 87 ][ 106 ],
   alphaCSR[ 87 ][ 107 ],
   alphaCSR[ 87 ][ 108 ],
   alphaCSR[ 87 ][ 109 ],
   alphaCSR[ 87 ][ 110 ],
   alphaCSR[ 87 ][ 111 ],
   alphaCSR[ 87 ][ 112 ],
   alphaCSR[ 87 ][ 113 ],
   alphaCSR[ 87 ][ 114 ],
   alphaCSR[ 87 ][ 115 ],
   alphaCSR[ 87 ][ 116 ],
   alphaCSR[ 87 ][ 117 ],
   alphaCSR[ 87 ][ 118 ],
   alphaCSR[ 87 ][ 119 ],
   alphaCSR[ 87 ][ 120 ],
   alphaCSR[ 87 ][ 121 ],
   alphaCSR[ 87 ][ 122 ],
   alphaCSR[ 87 ][ 123 ],
   alphaCSR[ 87 ][ 124 ],
   alphaCSR[ 87 ][ 125 ],
   alphaCSR[ 87 ][ 126 ],
   alphaCSR[ 87 ][ 127 ],
   alphaCSR[ 87 ][ 128 ],
   alphaCSR[ 87 ][ 129 ],
   alphaCSR[ 87 ][ 130 ],
   alphaCSR[ 87 ][ 131 ],
   alphaCSR[ 87 ][ 132 ],
   alphaCSR[ 87 ][ 133 ],
   alphaCSR[ 87 ][ 134 ],
   alphaCSR[ 87 ][ 135 ],
   alphaCSR[ 87 ][ 136 ],
   alphaCSR[ 87 ][ 137 ],
   alphaCSR[ 87 ][ 138 ],
   alphaCSR[ 87 ][ 139 ],
   alphaCSR[ 87 ][ 140 ],
   alphaCSR[ 87 ][ 141 ],
   alphaCSR[ 87 ][ 142 ],
   alphaCSR[ 87 ][ 143 ],
   alphaCSR[ 87 ][ 144 ],
   alphaCSR[ 87 ][ 145 ],
   alphaCSR[ 87 ][ 146 ],
   alphaCSR[ 87 ][ 147 ],
   alphaCSR[ 87 ][ 148 ],
   alphaCSR[ 87 ][ 149 ],
   alphaCSR[ 87 ][ 150 ],
   alphaCSR[ 87 ][ 151 ],
   alphaCSR[ 87 ][ 152 ],
   alphaCSR[ 87 ][ 153 ],
   alphaCSR[ 87 ][ 154 ],
   alphaCSR[ 87 ][ 155 ],
   alphaCSR[ 87 ][ 156 ],
   alphaCSR[ 87 ][ 157 ],
   alphaCSR[ 87 ][ 158 ],
   alphaCSR[ 87 ][ 159 ],
   alphaCSR[ 87 ][ 160 ],
   alphaCSR[ 87 ][ 161 ],
   alphaCSR[ 87 ][ 162 ],
   alphaCSR[ 87 ][ 163 ],
   alphaCSR[ 87 ][ 164 ],
   alphaCSR[ 87 ][ 165 ],
   alphaCSR[ 87 ][ 166 ],
   alphaCSR[ 87 ][ 167 ],
   alphaCSR[ 87 ][ 168 ],
   alphaCSR[ 87 ][ 169 ],
   alphaCSR[ 87 ][ 170 ],
   alphaCSR[ 87 ][ 171 ],
   alphaCSR[ 87 ][ 172 ],
   alphaCSR[ 87 ][ 173 ],
   alphaCSR[ 87 ][ 174 ],
   alphaCSR[ 87 ][ 175 ],
   alphaCSR[ 87 ][ 176 ],
   alphaCSR[ 87 ][ 177 ],
   alphaCSR[ 87 ][ 178 ],
   alphaCSR[ 87 ][ 179 ],
   alphaCSR[ 87 ][ 180 ],
   alphaCSR[ 87 ][ 181 ],
   alphaCSR[ 87 ][ 182 ],
   alphaCSR[ 87 ][ 183 ],
   alphaCSR[ 87 ][ 184 ],
   alphaCSR[ 87 ][ 185 ],
   alphaCSR[ 87 ][ 186 ],
   alphaCSR[ 87 ][ 187 ],
   alphaCSR[ 87 ][ 188 ],
   alphaCSR[ 87 ][ 189 ],
   alphaCSR[ 87 ][ 190 ],
   alphaCSR[ 87 ][ 191 ],
   alphaCSR[ 87 ][ 192 ],
   alphaCSR[ 87 ][ 193 ],
   alphaCSR[ 87 ][ 194 ],
   alphaCSR[ 87 ][ 195 ],
   alphaCSR[ 87 ][ 196 ],
   alphaCSR[ 87 ][ 197 ],
   alphaCSR[ 87 ][ 198 ],
   alphaCSR[ 87 ][ 199 ],
   alphaCSR[ 87 ][ 200 ],
   alphaCSR[ 87 ][ 201 ],
   alphaCSR[ 87 ][ 202 ],
   alphaCSR[ 87 ][ 203 ],
   alphaCSR[ 87 ][ 204 ],
   alphaCSR[ 87 ][ 205 ],
   alphaCSR[ 87 ][ 206 ],
   alphaCSR[ 87 ][ 207 ],
   alphaCSR[ 87 ][ 208 ],
   alphaCSR[ 87 ][ 209 ],
   alphaCSR[ 87 ][ 210 ],
   alphaCSR[ 87 ][ 211 ],
   alphaCSR[ 87 ][ 212 ],
   alphaCSR[ 87 ][ 213 ],
   alphaCSR[ 87 ][ 214 ],
   alphaCSR[ 87 ][ 215 ],
   alphaCSR[ 87 ][ 216 ],
   alphaCSR[ 87 ][ 217 ],
   alphaCSR[ 87 ][ 218 ],
   alphaCSR[ 87 ][ 219 ],
   alphaCSR[ 87 ][ 220 ],
   alphaCSR[ 87 ][ 221 ],
   alphaCSR[ 87 ][ 222 ],
   alphaCSR[ 87 ][ 223 ],
   alphaCSR[ 87 ][ 224 ],
   alphaCSR[ 87 ][ 225 ],
   alphaCSR[ 87 ][ 226 ],
   alphaCSR[ 87 ][ 227 ],
   alphaCSR[ 87 ][ 228 ],
   alphaCSR[ 87 ][ 229 ],
   alphaCSR[ 87 ][ 230 ],
   alphaCSR[ 87 ][ 231 ],
   alphaCSR[ 87 ][ 232 ],
   alphaCSR[ 87 ][ 233 ],
   alphaCSR[ 87 ][ 234 ],
   alphaCSR[ 87 ][ 235 ],
   alphaCSR[ 87 ][ 236 ],
   alphaCSR[ 87 ][ 237 ],
   alphaCSR[ 87 ][ 238 ],
   alphaCSR[ 87 ][ 239 ],
   alphaCSR[ 87 ][ 240 ],
   alphaCSR[ 87 ][ 241 ],
   alphaCSR[ 87 ][ 242 ],
   alphaCSR[ 87 ][ 243 ],
   alphaCSR[ 87 ][ 244 ],
   alphaCSR[ 87 ][ 245 ],
   alphaCSR[ 87 ][ 246 ],
   alphaCSR[ 87 ][ 247 ],
   alphaCSR[ 87 ][ 248 ],
   alphaCSR[ 87 ][ 249 ],
   alphaCSR[ 87 ][ 250 ],
   alphaCSR[ 87 ][ 251 ],
   alphaCSR[ 87 ][ 252 ],
   alphaCSR[ 87 ][ 253 ],
   alphaCSR[ 87 ][ 254 ],
   alphaCSR[ 87 ][ 255 ],
   alphaCSR[ 87 ][ 256 ],
   alphaCSR[ 87 ][ 257 ],
   alphaCSR[ 87 ][ 258 ],
   alphaCSR[ 87 ][ 259 ],
   alphaCSR[ 87 ][ 260 ],
   alphaCSR[ 87 ][ 261 ],
   alphaCSR[ 87 ][ 262 ],
   alphaCSR[ 87 ][ 263 ],
   alphaCSR[ 87 ][ 264 ],
   alphaCSR[ 87 ][ 265 ],
   alphaCSR[ 87 ][ 266 ],
   alphaCSR[ 87 ][ 267 ],
   alphaCSR[ 87 ][ 268 ],
   alphaCSR[ 87 ][ 269 ],
   alphaCSR[ 87 ][ 270 ],
   alphaCSR[ 87 ][ 271 ],
   alphaCSR[ 87 ][ 272 ],
   alphaCSR[ 87 ][ 273 ],
   alphaCSR[ 87 ][ 274 ],
   alphaCSR[ 87 ][ 275 ],
   alphaCSR[ 87 ][ 276 ],
   alphaCSR[ 87 ][ 277 ],
   alphaCSR[ 87 ][ 278 ],
   alphaCSR[ 87 ][ 279 ],
   alphaCSR[ 87 ][ 280 ],
   alphaCSR[ 87 ][ 281 ],
   alphaCSR[ 87 ][ 282 ],
   alphaCSR[ 87 ][ 283 ],
   alphaCSR[ 87 ][ 284 ],
   alphaCSR[ 87 ][ 285 ],
   alphaCSR[ 87 ][ 286 ],
   alphaCSR[ 87 ][ 287 ],
   alphaCSR[ 87 ][ 288 ],
   alphaCSR[ 87 ][ 289 ],
   alphaCSR[ 87 ][ 290 ],
   alphaCSR[ 87 ][ 291 ],
   alphaCSR[ 87 ][ 292 ],
   alphaCSR[ 87 ][ 293 ],
   alphaCSR[ 87 ][ 294 ],
   alphaCSR[ 87 ][ 295 ],
   alphaCSR[ 87 ][ 296 ],
   alphaCSR[ 87 ][ 297 ],
   alphaCSR[ 87 ][ 298 ],
   alphaCSR[ 87 ][ 299 ],
   alphaCSR[ 87 ][ 300 ],
   alphaCSR[ 87 ][ 301 ],
   alphaCSR[ 87 ][ 302 ],
   alphaCSR[ 87 ][ 303 ],
   alphaCSR[ 87 ][ 304 ],
   alphaCSR[ 87 ][ 305 ],
   alphaCSR[ 87 ][ 306 ],
   alphaCSR[ 87 ][ 307 ],
   alphaCSR[ 87 ][ 308 ],
   alphaCSR[ 87 ][ 309 ],
   alphaCSR[ 87 ][ 310 ],
   alphaCSR[ 87 ][ 311 ],
   alphaCSR[ 87 ][ 312 ],
   alphaCSR[ 87 ][ 313 ],
   alphaCSR[ 87 ][ 314 ],
   alphaCSR[ 87 ][ 315 ],
   alphaCSR[ 87 ][ 316 ],
   alphaCSR[ 87 ][ 317 ],
   alphaCSR[ 87 ][ 318 ],
   alphaCSR[ 87 ][ 319 ],
   alphaCSR[ 87 ][ 320 ],
   alphaCSR[ 87 ][ 321 ],
   alphaCSR[ 87 ][ 322 ],
   alphaCSR[ 87 ][ 323 ],
   alphaCSR[ 87 ][ 324 ],
   alphaCSR[ 87 ][ 325 ],
   alphaCSR[ 87 ][ 326 ],
   alphaCSR[ 87 ][ 327 ],
   alphaCSR[ 87 ][ 328 ],
   alphaCSR[ 87 ][ 329 ],
   alphaCSR[ 87 ][ 330 ],
   alphaCSR[ 87 ][ 331 ],
   alphaCSR[ 87 ][ 332 ],
   alphaCSR[ 87 ][ 333 ],
   alphaCSR[ 87 ][ 334 ],
   alphaCSR[ 87 ][ 335 ],
   alphaCSR[ 87 ][ 336 ],
   alphaCSR[ 87 ][ 337 ],
   alphaCSR[ 87 ][ 338 ],
   alphaCSR[ 87 ][ 339 ],
   alphaCSR[ 87 ][ 340 ],
   alphaCSR[ 87 ][ 341 ],
   alphaCSR[ 87 ][ 342 ],
   alphaCSR[ 87 ][ 343 ],
   alphaCSR[ 87 ][ 344 ],
   alphaCSR[ 87 ][ 345 ],
   alphaCSR[ 87 ][ 346 ],
   alphaCSR[ 87 ][ 347 ],
   alphaCSR[ 87 ][ 348 ],
   alphaCSR[ 87 ][ 349 ],
   alphaCSR[ 87 ][ 350 ],
   alphaCSR[ 87 ][ 351 ],
   alphaCSR[ 87 ][ 352 ],
   alphaCSR[ 87 ][ 353 ],
   alphaCSR[ 87 ][ 354 ],
   alphaCSR[ 87 ][ 355 ],
   alphaCSR[ 87 ][ 356 ],
   alphaCSR[ 87 ][ 357 ],
   alphaCSR[ 87 ][ 358 ],
   alphaCSR[ 87 ][ 359 ],
   alphaCSR[ 87 ][ 360 ],
   alphaCSR[ 87 ][ 361 ],
   alphaCSR[ 87 ][ 362 ],
   alphaCSR[ 87 ][ 363 ],
   alphaCSR[ 87 ][ 364 ],
   alphaCSR[ 87 ][ 365 ],
   alphaCSR[ 87 ][ 366 ],
   alphaCSR[ 87 ][ 367 ],
   alphaCSR[ 87 ][ 368 ],
   alphaCSR[ 87 ][ 369 ],
   alphaCSR[ 87 ][ 370 ],
   alphaCSR[ 87 ][ 371 ],
   alphaCSR[ 87 ][ 372 ],
   alphaCSR[ 87 ][ 373 ],
   alphaCSR[ 87 ][ 374 ],
   alphaCSR[ 87 ][ 375 ],
   alphaCSR[ 87 ][ 376 ],
   alphaCSR[ 87 ][ 377 ],
   alphaCSR[ 87 ][ 378 ],
   alphaCSR[ 87 ][ 379 ],
   alphaCSR[ 87 ][ 380 ],
   alphaCSR[ 87 ][ 381 ],
   alphaCSR[ 87 ][ 382 ],
   alphaCSR[ 87 ][ 383 ],
   alphaCSR[ 88 ][ 0 ],
   alphaCSR[ 88 ][ 1 ],
   alphaCSR[ 88 ][ 2 ],
   alphaCSR[ 88 ][ 3 ],
   alphaCSR[ 88 ][ 4 ],
   alphaCSR[ 88 ][ 5 ],
   alphaCSR[ 88 ][ 6 ],
   alphaCSR[ 88 ][ 7 ],
   alphaCSR[ 88 ][ 8 ],
   alphaCSR[ 88 ][ 9 ],
   alphaCSR[ 88 ][ 10 ],
   alphaCSR[ 88 ][ 11 ],
   alphaCSR[ 88 ][ 12 ],
   alphaCSR[ 88 ][ 13 ],
   alphaCSR[ 88 ][ 14 ],
   alphaCSR[ 88 ][ 15 ],
   alphaCSR[ 88 ][ 16 ],
   alphaCSR[ 88 ][ 17 ],
   alphaCSR[ 88 ][ 18 ],
   alphaCSR[ 88 ][ 19 ],
   alphaCSR[ 88 ][ 20 ],
   alphaCSR[ 88 ][ 21 ],
   alphaCSR[ 88 ][ 22 ],
   alphaCSR[ 88 ][ 23 ],
   alphaCSR[ 88 ][ 24 ],
   alphaCSR[ 88 ][ 25 ],
   alphaCSR[ 88 ][ 26 ],
   alphaCSR[ 88 ][ 27 ],
   alphaCSR[ 88 ][ 28 ],
   alphaCSR[ 88 ][ 29 ],
   alphaCSR[ 88 ][ 30 ],
   alphaCSR[ 88 ][ 31 ],
   alphaCSR[ 88 ][ 32 ],
   alphaCSR[ 88 ][ 33 ],
   alphaCSR[ 88 ][ 34 ],
   alphaCSR[ 88 ][ 35 ],
   alphaCSR[ 88 ][ 36 ],
   alphaCSR[ 88 ][ 37 ],
   alphaCSR[ 88 ][ 38 ],
   alphaCSR[ 88 ][ 39 ],
   alphaCSR[ 88 ][ 40 ],
   alphaCSR[ 88 ][ 41 ],
   alphaCSR[ 88 ][ 42 ],
   alphaCSR[ 88 ][ 43 ],
   alphaCSR[ 88 ][ 44 ],
   alphaCSR[ 88 ][ 45 ],
   alphaCSR[ 88 ][ 46 ],
   alphaCSR[ 88 ][ 47 ],
   alphaCSR[ 88 ][ 48 ],
   alphaCSR[ 88 ][ 49 ],
   alphaCSR[ 88 ][ 50 ],
   alphaCSR[ 88 ][ 51 ],
   alphaCSR[ 88 ][ 52 ],
   alphaCSR[ 88 ][ 53 ],
   alphaCSR[ 88 ][ 54 ],
   alphaCSR[ 88 ][ 55 ],
   alphaCSR[ 88 ][ 56 ],
   alphaCSR[ 88 ][ 57 ],
   alphaCSR[ 88 ][ 58 ],
   alphaCSR[ 88 ][ 59 ],
   alphaCSR[ 88 ][ 60 ],
   alphaCSR[ 88 ][ 61 ],
   alphaCSR[ 88 ][ 62 ],
   alphaCSR[ 88 ][ 63 ],
   alphaCSR[ 88 ][ 64 ],
   alphaCSR[ 88 ][ 65 ],
   alphaCSR[ 88 ][ 66 ],
   alphaCSR[ 88 ][ 67 ],
   alphaCSR[ 88 ][ 68 ],
   alphaCSR[ 88 ][ 69 ],
   alphaCSR[ 88 ][ 70 ],
   alphaCSR[ 88 ][ 71 ],
   alphaCSR[ 88 ][ 72 ],
   alphaCSR[ 88 ][ 73 ],
   alphaCSR[ 88 ][ 74 ],
   alphaCSR[ 88 ][ 75 ],
   alphaCSR[ 88 ][ 76 ],
   alphaCSR[ 88 ][ 77 ],
   alphaCSR[ 88 ][ 78 ],
   alphaCSR[ 88 ][ 79 ],
   alphaCSR[ 88 ][ 80 ],
   alphaCSR[ 88 ][ 81 ],
   alphaCSR[ 88 ][ 82 ],
   alphaCSR[ 88 ][ 83 ],
   alphaCSR[ 88 ][ 84 ],
   alphaCSR[ 88 ][ 85 ],
   alphaCSR[ 88 ][ 86 ],
   alphaCSR[ 88 ][ 87 ],
   alphaCSR[ 88 ][ 88 ],
   alphaCSR[ 88 ][ 89 ],
   alphaCSR[ 88 ][ 90 ],
   alphaCSR[ 88 ][ 91 ],
   alphaCSR[ 88 ][ 92 ],
   alphaCSR[ 88 ][ 93 ],
   alphaCSR[ 88 ][ 94 ],
   alphaCSR[ 88 ][ 95 ],
   alphaCSR[ 88 ][ 96 ],
   alphaCSR[ 88 ][ 97 ],
   alphaCSR[ 88 ][ 98 ],
   alphaCSR[ 88 ][ 99 ],
   alphaCSR[ 88 ][ 100 ],
   alphaCSR[ 88 ][ 101 ],
   alphaCSR[ 88 ][ 102 ],
   alphaCSR[ 88 ][ 103 ],
   alphaCSR[ 88 ][ 104 ],
   alphaCSR[ 88 ][ 105 ],
   alphaCSR[ 88 ][ 106 ],
   alphaCSR[ 88 ][ 107 ],
   alphaCSR[ 88 ][ 108 ],
   alphaCSR[ 88 ][ 109 ],
   alphaCSR[ 88 ][ 110 ],
   alphaCSR[ 88 ][ 111 ],
   alphaCSR[ 88 ][ 112 ],
   alphaCSR[ 88 ][ 113 ],
   alphaCSR[ 88 ][ 114 ],
   alphaCSR[ 88 ][ 115 ],
   alphaCSR[ 88 ][ 116 ],
   alphaCSR[ 88 ][ 117 ],
   alphaCSR[ 88 ][ 118 ],
   alphaCSR[ 88 ][ 119 ],
   alphaCSR[ 88 ][ 120 ],
   alphaCSR[ 88 ][ 121 ],
   alphaCSR[ 88 ][ 122 ],
   alphaCSR[ 88 ][ 123 ],
   alphaCSR[ 88 ][ 124 ],
   alphaCSR[ 88 ][ 125 ],
   alphaCSR[ 88 ][ 126 ],
   alphaCSR[ 88 ][ 127 ],
   alphaCSR[ 88 ][ 128 ],
   alphaCSR[ 88 ][ 129 ],
   alphaCSR[ 88 ][ 130 ],
   alphaCSR[ 88 ][ 131 ],
   alphaCSR[ 88 ][ 132 ],
   alphaCSR[ 88 ][ 133 ],
   alphaCSR[ 88 ][ 134 ],
   alphaCSR[ 88 ][ 135 ],
   alphaCSR[ 88 ][ 136 ],
   alphaCSR[ 88 ][ 137 ],
   alphaCSR[ 88 ][ 138 ],
   alphaCSR[ 88 ][ 139 ],
   alphaCSR[ 88 ][ 140 ],
   alphaCSR[ 88 ][ 141 ],
   alphaCSR[ 88 ][ 142 ],
   alphaCSR[ 88 ][ 143 ],
   alphaCSR[ 88 ][ 144 ],
   alphaCSR[ 88 ][ 145 ],
   alphaCSR[ 88 ][ 146 ],
   alphaCSR[ 88 ][ 147 ],
   alphaCSR[ 88 ][ 148 ],
   alphaCSR[ 88 ][ 149 ],
   alphaCSR[ 88 ][ 150 ],
   alphaCSR[ 88 ][ 151 ],
   alphaCSR[ 88 ][ 152 ],
   alphaCSR[ 88 ][ 153 ],
   alphaCSR[ 88 ][ 154 ],
   alphaCSR[ 88 ][ 155 ],
   alphaCSR[ 88 ][ 156 ],
   alphaCSR[ 88 ][ 157 ],
   alphaCSR[ 88 ][ 158 ],
   alphaCSR[ 88 ][ 159 ],
   alphaCSR[ 88 ][ 160 ],
   alphaCSR[ 88 ][ 161 ],
   alphaCSR[ 88 ][ 162 ],
   alphaCSR[ 88 ][ 163 ],
   alphaCSR[ 88 ][ 164 ],
   alphaCSR[ 88 ][ 165 ],
   alphaCSR[ 88 ][ 166 ],
   alphaCSR[ 88 ][ 167 ],
   alphaCSR[ 88 ][ 168 ],
   alphaCSR[ 88 ][ 169 ],
   alphaCSR[ 88 ][ 170 ],
   alphaCSR[ 88 ][ 171 ],
   alphaCSR[ 88 ][ 172 ],
   alphaCSR[ 88 ][ 173 ],
   alphaCSR[ 88 ][ 174 ],
   alphaCSR[ 88 ][ 175 ],
   alphaCSR[ 88 ][ 176 ],
   alphaCSR[ 88 ][ 177 ],
   alphaCSR[ 88 ][ 178 ],
   alphaCSR[ 88 ][ 179 ],
   alphaCSR[ 88 ][ 180 ],
   alphaCSR[ 88 ][ 181 ],
   alphaCSR[ 88 ][ 182 ],
   alphaCSR[ 88 ][ 183 ],
   alphaCSR[ 88 ][ 184 ],
   alphaCSR[ 88 ][ 185 ],
   alphaCSR[ 88 ][ 186 ],
   alphaCSR[ 88 ][ 187 ],
   alphaCSR[ 88 ][ 188 ],
   alphaCSR[ 88 ][ 189 ],
   alphaCSR[ 88 ][ 190 ],
   alphaCSR[ 88 ][ 191 ],
   alphaCSR[ 88 ][ 192 ],
   alphaCSR[ 88 ][ 193 ],
   alphaCSR[ 88 ][ 194 ],
   alphaCSR[ 88 ][ 195 ],
   alphaCSR[ 88 ][ 196 ],
   alphaCSR[ 88 ][ 197 ],
   alphaCSR[ 88 ][ 198 ],
   alphaCSR[ 88 ][ 199 ],
   alphaCSR[ 88 ][ 200 ],
   alphaCSR[ 88 ][ 201 ],
   alphaCSR[ 88 ][ 202 ],
   alphaCSR[ 88 ][ 203 ],
   alphaCSR[ 88 ][ 204 ],
   alphaCSR[ 88 ][ 205 ],
   alphaCSR[ 88 ][ 206 ],
   alphaCSR[ 88 ][ 207 ],
   alphaCSR[ 88 ][ 208 ],
   alphaCSR[ 88 ][ 209 ],
   alphaCSR[ 88 ][ 210 ],
   alphaCSR[ 88 ][ 211 ],
   alphaCSR[ 88 ][ 212 ],
   alphaCSR[ 88 ][ 213 ],
   alphaCSR[ 88 ][ 214 ],
   alphaCSR[ 88 ][ 215 ],
   alphaCSR[ 88 ][ 216 ],
   alphaCSR[ 88 ][ 217 ],
   alphaCSR[ 88 ][ 218 ],
   alphaCSR[ 88 ][ 219 ],
   alphaCSR[ 88 ][ 220 ],
   alphaCSR[ 88 ][ 221 ],
   alphaCSR[ 88 ][ 222 ],
   alphaCSR[ 88 ][ 223 ],
   alphaCSR[ 88 ][ 224 ],
   alphaCSR[ 88 ][ 225 ],
   alphaCSR[ 88 ][ 226 ],
   alphaCSR[ 88 ][ 227 ],
   alphaCSR[ 88 ][ 228 ],
   alphaCSR[ 88 ][ 229 ],
   alphaCSR[ 88 ][ 230 ],
   alphaCSR[ 88 ][ 231 ],
   alphaCSR[ 88 ][ 232 ],
   alphaCSR[ 88 ][ 233 ],
   alphaCSR[ 88 ][ 234 ],
   alphaCSR[ 88 ][ 235 ],
   alphaCSR[ 88 ][ 236 ],
   alphaCSR[ 88 ][ 237 ],
   alphaCSR[ 88 ][ 238 ],
   alphaCSR[ 88 ][ 239 ],
   alphaCSR[ 88 ][ 240 ],
   alphaCSR[ 88 ][ 241 ],
   alphaCSR[ 88 ][ 242 ],
   alphaCSR[ 88 ][ 243 ],
   alphaCSR[ 88 ][ 244 ],
   alphaCSR[ 88 ][ 245 ],
   alphaCSR[ 88 ][ 246 ],
   alphaCSR[ 88 ][ 247 ],
   alphaCSR[ 88 ][ 248 ],
   alphaCSR[ 88 ][ 249 ],
   alphaCSR[ 88 ][ 250 ],
   alphaCSR[ 88 ][ 251 ],
   alphaCSR[ 88 ][ 252 ],
   alphaCSR[ 88 ][ 253 ],
   alphaCSR[ 88 ][ 254 ],
   alphaCSR[ 88 ][ 255 ],
   alphaCSR[ 88 ][ 256 ],
   alphaCSR[ 88 ][ 257 ],
   alphaCSR[ 88 ][ 258 ],
   alphaCSR[ 88 ][ 259 ],
   alphaCSR[ 88 ][ 260 ],
   alphaCSR[ 88 ][ 261 ],
   alphaCSR[ 88 ][ 262 ],
   alphaCSR[ 88 ][ 263 ],
   alphaCSR[ 88 ][ 264 ],
   alphaCSR[ 88 ][ 265 ],
   alphaCSR[ 88 ][ 266 ],
   alphaCSR[ 88 ][ 267 ],
   alphaCSR[ 88 ][ 268 ],
   alphaCSR[ 88 ][ 269 ],
   alphaCSR[ 88 ][ 270 ],
   alphaCSR[ 88 ][ 271 ],
   alphaCSR[ 88 ][ 272 ],
   alphaCSR[ 88 ][ 273 ],
   alphaCSR[ 88 ][ 274 ],
   alphaCSR[ 88 ][ 275 ],
   alphaCSR[ 88 ][ 276 ],
   alphaCSR[ 88 ][ 277 ],
   alphaCSR[ 88 ][ 278 ],
   alphaCSR[ 88 ][ 279 ],
   alphaCSR[ 88 ][ 280 ],
   alphaCSR[ 88 ][ 281 ],
   alphaCSR[ 88 ][ 282 ],
   alphaCSR[ 88 ][ 283 ],
   alphaCSR[ 88 ][ 284 ],
   alphaCSR[ 88 ][ 285 ],
   alphaCSR[ 88 ][ 286 ],
   alphaCSR[ 88 ][ 287 ],
   alphaCSR[ 88 ][ 288 ],
   alphaCSR[ 88 ][ 289 ],
   alphaCSR[ 88 ][ 290 ],
   alphaCSR[ 88 ][ 291 ],
   alphaCSR[ 88 ][ 292 ],
   alphaCSR[ 88 ][ 293 ],
   alphaCSR[ 88 ][ 294 ],
   alphaCSR[ 88 ][ 295 ],
   alphaCSR[ 88 ][ 296 ],
   alphaCSR[ 88 ][ 297 ],
   alphaCSR[ 88 ][ 298 ],
   alphaCSR[ 88 ][ 299 ],
   alphaCSR[ 88 ][ 300 ],
   alphaCSR[ 88 ][ 301 ],
   alphaCSR[ 88 ][ 302 ],
   alphaCSR[ 88 ][ 303 ],
   alphaCSR[ 88 ][ 304 ],
   alphaCSR[ 88 ][ 305 ],
   alphaCSR[ 88 ][ 306 ],
   alphaCSR[ 88 ][ 307 ],
   alphaCSR[ 88 ][ 308 ],
   alphaCSR[ 88 ][ 309 ],
   alphaCSR[ 88 ][ 310 ],
   alphaCSR[ 88 ][ 311 ],
   alphaCSR[ 88 ][ 312 ],
   alphaCSR[ 88 ][ 313 ],
   alphaCSR[ 88 ][ 314 ],
   alphaCSR[ 88 ][ 315 ],
   alphaCSR[ 88 ][ 316 ],
   alphaCSR[ 88 ][ 317 ],
   alphaCSR[ 88 ][ 318 ],
   alphaCSR[ 88 ][ 319 ],
   alphaCSR[ 88 ][ 320 ],
   alphaCSR[ 88 ][ 321 ],
   alphaCSR[ 88 ][ 322 ],
   alphaCSR[ 88 ][ 323 ],
   alphaCSR[ 88 ][ 324 ],
   alphaCSR[ 88 ][ 325 ],
   alphaCSR[ 88 ][ 326 ],
   alphaCSR[ 88 ][ 327 ],
   alphaCSR[ 88 ][ 328 ],
   alphaCSR[ 88 ][ 329 ],
   alphaCSR[ 88 ][ 330 ],
   alphaCSR[ 88 ][ 331 ],
   alphaCSR[ 88 ][ 332 ],
   alphaCSR[ 88 ][ 333 ],
   alphaCSR[ 88 ][ 334 ],
   alphaCSR[ 88 ][ 335 ],
   alphaCSR[ 88 ][ 336 ],
   alphaCSR[ 88 ][ 337 ],
   alphaCSR[ 88 ][ 338 ],
   alphaCSR[ 88 ][ 339 ],
   alphaCSR[ 88 ][ 340 ],
   alphaCSR[ 88 ][ 341 ],
   alphaCSR[ 88 ][ 342 ],
   alphaCSR[ 88 ][ 343 ],
   alphaCSR[ 88 ][ 344 ],
   alphaCSR[ 88 ][ 345 ],
   alphaCSR[ 88 ][ 346 ],
   alphaCSR[ 88 ][ 347 ],
   alphaCSR[ 88 ][ 348 ],
   alphaCSR[ 88 ][ 349 ],
   alphaCSR[ 88 ][ 350 ],
   alphaCSR[ 88 ][ 351 ],
   alphaCSR[ 88 ][ 352 ],
   alphaCSR[ 88 ][ 353 ],
   alphaCSR[ 88 ][ 354 ],
   alphaCSR[ 88 ][ 355 ],
   alphaCSR[ 88 ][ 356 ],
   alphaCSR[ 88 ][ 357 ],
   alphaCSR[ 88 ][ 358 ],
   alphaCSR[ 88 ][ 359 ],
   alphaCSR[ 88 ][ 360 ],
   alphaCSR[ 88 ][ 361 ],
   alphaCSR[ 88 ][ 362 ],
   alphaCSR[ 88 ][ 363 ],
   alphaCSR[ 88 ][ 364 ],
   alphaCSR[ 88 ][ 365 ],
   alphaCSR[ 88 ][ 366 ],
   alphaCSR[ 88 ][ 367 ],
   alphaCSR[ 88 ][ 368 ],
   alphaCSR[ 88 ][ 369 ],
   alphaCSR[ 88 ][ 370 ],
   alphaCSR[ 88 ][ 371 ],
   alphaCSR[ 88 ][ 372 ],
   alphaCSR[ 88 ][ 373 ],
   alphaCSR[ 88 ][ 374 ],
   alphaCSR[ 88 ][ 375 ],
   alphaCSR[ 88 ][ 376 ],
   alphaCSR[ 88 ][ 377 ],
   alphaCSR[ 88 ][ 378 ],
   alphaCSR[ 88 ][ 379 ],
   alphaCSR[ 88 ][ 380 ],
   alphaCSR[ 88 ][ 381 ],
   alphaCSR[ 88 ][ 382 ],
   alphaCSR[ 88 ][ 383 ],
   alphaCSR[ 89 ][ 0 ],
   alphaCSR[ 89 ][ 1 ],
   alphaCSR[ 89 ][ 2 ],
   alphaCSR[ 89 ][ 3 ],
   alphaCSR[ 89 ][ 4 ],
   alphaCSR[ 89 ][ 5 ],
   alphaCSR[ 89 ][ 6 ],
   alphaCSR[ 89 ][ 7 ],
   alphaCSR[ 89 ][ 8 ],
   alphaCSR[ 89 ][ 9 ],
   alphaCSR[ 89 ][ 10 ],
   alphaCSR[ 89 ][ 11 ],
   alphaCSR[ 89 ][ 12 ],
   alphaCSR[ 89 ][ 13 ],
   alphaCSR[ 89 ][ 14 ],
   alphaCSR[ 89 ][ 15 ],
   alphaCSR[ 89 ][ 16 ],
   alphaCSR[ 89 ][ 17 ],
   alphaCSR[ 89 ][ 18 ],
   alphaCSR[ 89 ][ 19 ],
   alphaCSR[ 89 ][ 20 ],
   alphaCSR[ 89 ][ 21 ],
   alphaCSR[ 89 ][ 22 ],
   alphaCSR[ 89 ][ 23 ],
   alphaCSR[ 89 ][ 24 ],
   alphaCSR[ 89 ][ 25 ],
   alphaCSR[ 89 ][ 26 ],
   alphaCSR[ 89 ][ 27 ],
   alphaCSR[ 89 ][ 28 ],
   alphaCSR[ 89 ][ 29 ],
   alphaCSR[ 89 ][ 30 ],
   alphaCSR[ 89 ][ 31 ],
   alphaCSR[ 89 ][ 32 ],
   alphaCSR[ 89 ][ 33 ],
   alphaCSR[ 89 ][ 34 ],
   alphaCSR[ 89 ][ 35 ],
   alphaCSR[ 89 ][ 36 ],
   alphaCSR[ 89 ][ 37 ],
   alphaCSR[ 89 ][ 38 ],
   alphaCSR[ 89 ][ 39 ],
   alphaCSR[ 89 ][ 40 ],
   alphaCSR[ 89 ][ 41 ],
   alphaCSR[ 89 ][ 42 ],
   alphaCSR[ 89 ][ 43 ],
   alphaCSR[ 89 ][ 44 ],
   alphaCSR[ 89 ][ 45 ],
   alphaCSR[ 89 ][ 46 ],
   alphaCSR[ 89 ][ 47 ],
   alphaCSR[ 89 ][ 48 ],
   alphaCSR[ 89 ][ 49 ],
   alphaCSR[ 89 ][ 50 ],
   alphaCSR[ 89 ][ 51 ],
   alphaCSR[ 89 ][ 52 ],
   alphaCSR[ 89 ][ 53 ],
   alphaCSR[ 89 ][ 54 ],
   alphaCSR[ 89 ][ 55 ],
   alphaCSR[ 89 ][ 56 ],
   alphaCSR[ 89 ][ 57 ],
   alphaCSR[ 89 ][ 58 ],
   alphaCSR[ 89 ][ 59 ],
   alphaCSR[ 89 ][ 60 ],
   alphaCSR[ 89 ][ 61 ],
   alphaCSR[ 89 ][ 62 ],
   alphaCSR[ 89 ][ 63 ],
   alphaCSR[ 89 ][ 64 ],
   alphaCSR[ 89 ][ 65 ],
   alphaCSR[ 89 ][ 66 ],
   alphaCSR[ 89 ][ 67 ],
   alphaCSR[ 89 ][ 68 ],
   alphaCSR[ 89 ][ 69 ],
   alphaCSR[ 89 ][ 70 ],
   alphaCSR[ 89 ][ 71 ],
   alphaCSR[ 89 ][ 72 ],
   alphaCSR[ 89 ][ 73 ],
   alphaCSR[ 89 ][ 74 ],
   alphaCSR[ 89 ][ 75 ],
   alphaCSR[ 89 ][ 76 ],
   alphaCSR[ 89 ][ 77 ],
   alphaCSR[ 89 ][ 78 ],
   alphaCSR[ 89 ][ 79 ],
   alphaCSR[ 89 ][ 80 ],
   alphaCSR[ 89 ][ 81 ],
   alphaCSR[ 89 ][ 82 ],
   alphaCSR[ 89 ][ 83 ],
   alphaCSR[ 89 ][ 84 ],
   alphaCSR[ 89 ][ 85 ],
   alphaCSR[ 89 ][ 86 ],
   alphaCSR[ 89 ][ 87 ],
   alphaCSR[ 89 ][ 88 ],
   alphaCSR[ 89 ][ 89 ],
   alphaCSR[ 89 ][ 90 ],
   alphaCSR[ 89 ][ 91 ],
   alphaCSR[ 89 ][ 92 ],
   alphaCSR[ 89 ][ 93 ],
   alphaCSR[ 89 ][ 94 ],
   alphaCSR[ 89 ][ 95 ],
   alphaCSR[ 89 ][ 96 ],
   alphaCSR[ 89 ][ 97 ],
   alphaCSR[ 89 ][ 98 ],
   alphaCSR[ 89 ][ 99 ],
   alphaCSR[ 89 ][ 100 ],
   alphaCSR[ 89 ][ 101 ],
   alphaCSR[ 89 ][ 102 ],
   alphaCSR[ 89 ][ 103 ],
   alphaCSR[ 89 ][ 104 ],
   alphaCSR[ 89 ][ 105 ],
   alphaCSR[ 89 ][ 106 ],
   alphaCSR[ 89 ][ 107 ],
   alphaCSR[ 89 ][ 108 ],
   alphaCSR[ 89 ][ 109 ],
   alphaCSR[ 89 ][ 110 ],
   alphaCSR[ 89 ][ 111 ],
   alphaCSR[ 89 ][ 112 ],
   alphaCSR[ 89 ][ 113 ],
   alphaCSR[ 89 ][ 114 ],
   alphaCSR[ 89 ][ 115 ],
   alphaCSR[ 89 ][ 116 ],
   alphaCSR[ 89 ][ 117 ],
   alphaCSR[ 89 ][ 118 ],
   alphaCSR[ 89 ][ 119 ],
   alphaCSR[ 89 ][ 120 ],
   alphaCSR[ 89 ][ 121 ],
   alphaCSR[ 89 ][ 122 ],
   alphaCSR[ 89 ][ 123 ],
   alphaCSR[ 89 ][ 124 ],
   alphaCSR[ 89 ][ 125 ],
   alphaCSR[ 89 ][ 126 ],
   alphaCSR[ 89 ][ 127 ],
   alphaCSR[ 89 ][ 128 ],
   alphaCSR[ 89 ][ 129 ],
   alphaCSR[ 89 ][ 130 ],
   alphaCSR[ 89 ][ 131 ],
   alphaCSR[ 89 ][ 132 ],
   alphaCSR[ 89 ][ 133 ],
   alphaCSR[ 89 ][ 134 ],
   alphaCSR[ 89 ][ 135 ],
   alphaCSR[ 89 ][ 136 ],
   alphaCSR[ 89 ][ 137 ],
   alphaCSR[ 89 ][ 138 ],
   alphaCSR[ 89 ][ 139 ],
   alphaCSR[ 89 ][ 140 ],
   alphaCSR[ 89 ][ 141 ],
   alphaCSR[ 89 ][ 142 ],
   alphaCSR[ 89 ][ 143 ],
   alphaCSR[ 89 ][ 144 ],
   alphaCSR[ 89 ][ 145 ],
   alphaCSR[ 89 ][ 146 ],
   alphaCSR[ 89 ][ 147 ],
   alphaCSR[ 89 ][ 148 ],
   alphaCSR[ 89 ][ 149 ],
   alphaCSR[ 89 ][ 150 ],
   alphaCSR[ 89 ][ 151 ],
   alphaCSR[ 89 ][ 152 ],
   alphaCSR[ 89 ][ 153 ],
   alphaCSR[ 89 ][ 154 ],
   alphaCSR[ 89 ][ 155 ],
   alphaCSR[ 89 ][ 156 ],
   alphaCSR[ 89 ][ 157 ],
   alphaCSR[ 89 ][ 158 ],
   alphaCSR[ 89 ][ 159 ],
   alphaCSR[ 89 ][ 160 ],
   alphaCSR[ 89 ][ 161 ],
   alphaCSR[ 89 ][ 162 ],
   alphaCSR[ 89 ][ 163 ],
   alphaCSR[ 89 ][ 164 ],
   alphaCSR[ 89 ][ 165 ],
   alphaCSR[ 89 ][ 166 ],
   alphaCSR[ 89 ][ 167 ],
   alphaCSR[ 89 ][ 168 ],
   alphaCSR[ 89 ][ 169 ],
   alphaCSR[ 89 ][ 170 ],
   alphaCSR[ 89 ][ 171 ],
   alphaCSR[ 89 ][ 172 ],
   alphaCSR[ 89 ][ 173 ],
   alphaCSR[ 89 ][ 174 ],
   alphaCSR[ 89 ][ 175 ],
   alphaCSR[ 89 ][ 176 ],
   alphaCSR[ 89 ][ 177 ],
   alphaCSR[ 89 ][ 178 ],
   alphaCSR[ 89 ][ 179 ],
   alphaCSR[ 89 ][ 180 ],
   alphaCSR[ 89 ][ 181 ],
   alphaCSR[ 89 ][ 182 ],
   alphaCSR[ 89 ][ 183 ],
   alphaCSR[ 89 ][ 184 ],
   alphaCSR[ 89 ][ 185 ],
   alphaCSR[ 89 ][ 186 ],
   alphaCSR[ 89 ][ 187 ],
   alphaCSR[ 89 ][ 188 ],
   alphaCSR[ 89 ][ 189 ],
   alphaCSR[ 89 ][ 190 ],
   alphaCSR[ 89 ][ 191 ],
   alphaCSR[ 89 ][ 192 ],
   alphaCSR[ 89 ][ 193 ],
   alphaCSR[ 89 ][ 194 ],
   alphaCSR[ 89 ][ 195 ],
   alphaCSR[ 89 ][ 196 ],
   alphaCSR[ 89 ][ 197 ],
   alphaCSR[ 89 ][ 198 ],
   alphaCSR[ 89 ][ 199 ],
   alphaCSR[ 89 ][ 200 ],
   alphaCSR[ 89 ][ 201 ],
   alphaCSR[ 89 ][ 202 ],
   alphaCSR[ 89 ][ 203 ],
   alphaCSR[ 89 ][ 204 ],
   alphaCSR[ 89 ][ 205 ],
   alphaCSR[ 89 ][ 206 ],
   alphaCSR[ 89 ][ 207 ],
   alphaCSR[ 89 ][ 208 ],
   alphaCSR[ 89 ][ 209 ],
   alphaCSR[ 89 ][ 210 ],
   alphaCSR[ 89 ][ 211 ],
   alphaCSR[ 89 ][ 212 ],
   alphaCSR[ 89 ][ 213 ],
   alphaCSR[ 89 ][ 214 ],
   alphaCSR[ 89 ][ 215 ],
   alphaCSR[ 89 ][ 216 ],
   alphaCSR[ 89 ][ 217 ],
   alphaCSR[ 89 ][ 218 ],
   alphaCSR[ 89 ][ 219 ],
   alphaCSR[ 89 ][ 220 ],
   alphaCSR[ 89 ][ 221 ],
   alphaCSR[ 89 ][ 222 ],
   alphaCSR[ 89 ][ 223 ],
   alphaCSR[ 89 ][ 224 ],
   alphaCSR[ 89 ][ 225 ],
   alphaCSR[ 89 ][ 226 ],
   alphaCSR[ 89 ][ 227 ],
   alphaCSR[ 89 ][ 228 ],
   alphaCSR[ 89 ][ 229 ],
   alphaCSR[ 89 ][ 230 ],
   alphaCSR[ 89 ][ 231 ],
   alphaCSR[ 89 ][ 232 ],
   alphaCSR[ 89 ][ 233 ],
   alphaCSR[ 89 ][ 234 ],
   alphaCSR[ 89 ][ 235 ],
   alphaCSR[ 89 ][ 236 ],
   alphaCSR[ 89 ][ 237 ],
   alphaCSR[ 89 ][ 238 ],
   alphaCSR[ 89 ][ 239 ],
   alphaCSR[ 89 ][ 240 ],
   alphaCSR[ 89 ][ 241 ],
   alphaCSR[ 89 ][ 242 ],
   alphaCSR[ 89 ][ 243 ],
   alphaCSR[ 89 ][ 244 ],
   alphaCSR[ 89 ][ 245 ],
   alphaCSR[ 89 ][ 246 ],
   alphaCSR[ 89 ][ 247 ],
   alphaCSR[ 89 ][ 248 ],
   alphaCSR[ 89 ][ 249 ],
   alphaCSR[ 89 ][ 250 ],
   alphaCSR[ 89 ][ 251 ],
   alphaCSR[ 89 ][ 252 ],
   alphaCSR[ 89 ][ 253 ],
   alphaCSR[ 89 ][ 254 ],
   alphaCSR[ 89 ][ 255 ],
   alphaCSR[ 89 ][ 256 ],
   alphaCSR[ 89 ][ 257 ],
   alphaCSR[ 89 ][ 258 ],
   alphaCSR[ 89 ][ 259 ],
   alphaCSR[ 89 ][ 260 ],
   alphaCSR[ 89 ][ 261 ],
   alphaCSR[ 89 ][ 262 ],
   alphaCSR[ 89 ][ 263 ],
   alphaCSR[ 89 ][ 264 ],
   alphaCSR[ 89 ][ 265 ],
   alphaCSR[ 89 ][ 266 ],
   alphaCSR[ 89 ][ 267 ],
   alphaCSR[ 89 ][ 268 ],
   alphaCSR[ 89 ][ 269 ],
   alphaCSR[ 89 ][ 270 ],
   alphaCSR[ 89 ][ 271 ],
   alphaCSR[ 89 ][ 272 ],
   alphaCSR[ 89 ][ 273 ],
   alphaCSR[ 89 ][ 274 ],
   alphaCSR[ 89 ][ 275 ],
   alphaCSR[ 89 ][ 276 ],
   alphaCSR[ 89 ][ 277 ],
   alphaCSR[ 89 ][ 278 ],
   alphaCSR[ 89 ][ 279 ],
   alphaCSR[ 89 ][ 280 ],
   alphaCSR[ 89 ][ 281 ],
   alphaCSR[ 89 ][ 282 ],
   alphaCSR[ 89 ][ 283 ],
   alphaCSR[ 89 ][ 284 ],
   alphaCSR[ 89 ][ 285 ],
   alphaCSR[ 89 ][ 286 ],
   alphaCSR[ 89 ][ 287 ],
   alphaCSR[ 89 ][ 288 ],
   alphaCSR[ 89 ][ 289 ],
   alphaCSR[ 89 ][ 290 ],
   alphaCSR[ 89 ][ 291 ],
   alphaCSR[ 89 ][ 292 ],
   alphaCSR[ 89 ][ 293 ],
   alphaCSR[ 89 ][ 294 ],
   alphaCSR[ 89 ][ 295 ],
   alphaCSR[ 89 ][ 296 ],
   alphaCSR[ 89 ][ 297 ],
   alphaCSR[ 89 ][ 298 ],
   alphaCSR[ 89 ][ 299 ],
   alphaCSR[ 89 ][ 300 ],
   alphaCSR[ 89 ][ 301 ],
   alphaCSR[ 89 ][ 302 ],
   alphaCSR[ 89 ][ 303 ],
   alphaCSR[ 89 ][ 304 ],
   alphaCSR[ 89 ][ 305 ],
   alphaCSR[ 89 ][ 306 ],
   alphaCSR[ 89 ][ 307 ],
   alphaCSR[ 89 ][ 308 ],
   alphaCSR[ 89 ][ 309 ],
   alphaCSR[ 89 ][ 310 ],
   alphaCSR[ 89 ][ 311 ],
   alphaCSR[ 89 ][ 312 ],
   alphaCSR[ 89 ][ 313 ],
   alphaCSR[ 89 ][ 314 ],
   alphaCSR[ 89 ][ 315 ],
   alphaCSR[ 89 ][ 316 ],
   alphaCSR[ 89 ][ 317 ],
   alphaCSR[ 89 ][ 318 ],
   alphaCSR[ 89 ][ 319 ],
   alphaCSR[ 89 ][ 320 ],
   alphaCSR[ 89 ][ 321 ],
   alphaCSR[ 89 ][ 322 ],
   alphaCSR[ 89 ][ 323 ],
   alphaCSR[ 89 ][ 324 ],
   alphaCSR[ 89 ][ 325 ],
   alphaCSR[ 89 ][ 326 ],
   alphaCSR[ 89 ][ 327 ],
   alphaCSR[ 89 ][ 328 ],
   alphaCSR[ 89 ][ 329 ],
   alphaCSR[ 89 ][ 330 ],
   alphaCSR[ 89 ][ 331 ],
   alphaCSR[ 89 ][ 332 ],
   alphaCSR[ 89 ][ 333 ],
   alphaCSR[ 89 ][ 334 ],
   alphaCSR[ 89 ][ 335 ],
   alphaCSR[ 89 ][ 336 ],
   alphaCSR[ 89 ][ 337 ],
   alphaCSR[ 89 ][ 338 ],
   alphaCSR[ 89 ][ 339 ],
   alphaCSR[ 89 ][ 340 ],
   alphaCSR[ 89 ][ 341 ],
   alphaCSR[ 89 ][ 342 ],
   alphaCSR[ 89 ][ 343 ],
   alphaCSR[ 89 ][ 344 ],
   alphaCSR[ 89 ][ 345 ],
   alphaCSR[ 89 ][ 346 ],
   alphaCSR[ 89 ][ 347 ],
   alphaCSR[ 89 ][ 348 ],
   alphaCSR[ 89 ][ 349 ],
   alphaCSR[ 89 ][ 350 ],
   alphaCSR[ 89 ][ 351 ],
   alphaCSR[ 89 ][ 352 ],
   alphaCSR[ 89 ][ 353 ],
   alphaCSR[ 89 ][ 354 ],
   alphaCSR[ 89 ][ 355 ],
   alphaCSR[ 89 ][ 356 ],
   alphaCSR[ 89 ][ 357 ],
   alphaCSR[ 89 ][ 358 ],
   alphaCSR[ 89 ][ 359 ],
   alphaCSR[ 89 ][ 360 ],
   alphaCSR[ 89 ][ 361 ],
   alphaCSR[ 89 ][ 362 ],
   alphaCSR[ 89 ][ 363 ],
   alphaCSR[ 89 ][ 364 ],
   alphaCSR[ 89 ][ 365 ],
   alphaCSR[ 89 ][ 366 ],
   alphaCSR[ 89 ][ 367 ],
   alphaCSR[ 89 ][ 368 ],
   alphaCSR[ 89 ][ 369 ],
   alphaCSR[ 89 ][ 370 ],
   alphaCSR[ 89 ][ 371 ],
   alphaCSR[ 89 ][ 372 ],
   alphaCSR[ 89 ][ 373 ],
   alphaCSR[ 89 ][ 374 ],
   alphaCSR[ 89 ][ 375 ],
   alphaCSR[ 89 ][ 376 ],
   alphaCSR[ 89 ][ 377 ],
   alphaCSR[ 89 ][ 378 ],
   alphaCSR[ 89 ][ 379 ],
   alphaCSR[ 89 ][ 380 ],
   alphaCSR[ 89 ][ 381 ],
   alphaCSR[ 89 ][ 382 ],
   alphaCSR[ 89 ][ 383 ],
   alphaCSR[ 90 ][ 0 ],
   alphaCSR[ 90 ][ 1 ],
   alphaCSR[ 90 ][ 2 ],
   alphaCSR[ 90 ][ 3 ],
   alphaCSR[ 90 ][ 4 ],
   alphaCSR[ 90 ][ 5 ],
   alphaCSR[ 90 ][ 6 ],
   alphaCSR[ 90 ][ 7 ],
   alphaCSR[ 90 ][ 8 ],
   alphaCSR[ 90 ][ 9 ],
   alphaCSR[ 90 ][ 10 ],
   alphaCSR[ 90 ][ 11 ],
   alphaCSR[ 90 ][ 12 ],
   alphaCSR[ 90 ][ 13 ],
   alphaCSR[ 90 ][ 14 ],
   alphaCSR[ 90 ][ 15 ],
   alphaCSR[ 90 ][ 16 ],
   alphaCSR[ 90 ][ 17 ],
   alphaCSR[ 90 ][ 18 ],
   alphaCSR[ 90 ][ 19 ],
   alphaCSR[ 90 ][ 20 ],
   alphaCSR[ 90 ][ 21 ],
   alphaCSR[ 90 ][ 22 ],
   alphaCSR[ 90 ][ 23 ],
   alphaCSR[ 90 ][ 24 ],
   alphaCSR[ 90 ][ 25 ],
   alphaCSR[ 90 ][ 26 ],
   alphaCSR[ 90 ][ 27 ],
   alphaCSR[ 90 ][ 28 ],
   alphaCSR[ 90 ][ 29 ],
   alphaCSR[ 90 ][ 30 ],
   alphaCSR[ 90 ][ 31 ],
   alphaCSR[ 90 ][ 32 ],
   alphaCSR[ 90 ][ 33 ],
   alphaCSR[ 90 ][ 34 ],
   alphaCSR[ 90 ][ 35 ],
   alphaCSR[ 90 ][ 36 ],
   alphaCSR[ 90 ][ 37 ],
   alphaCSR[ 90 ][ 38 ],
   alphaCSR[ 90 ][ 39 ],
   alphaCSR[ 90 ][ 40 ],
   alphaCSR[ 90 ][ 41 ],
   alphaCSR[ 90 ][ 42 ],
   alphaCSR[ 90 ][ 43 ],
   alphaCSR[ 90 ][ 44 ],
   alphaCSR[ 90 ][ 45 ],
   alphaCSR[ 90 ][ 46 ],
   alphaCSR[ 90 ][ 47 ],
   alphaCSR[ 90 ][ 48 ],
   alphaCSR[ 90 ][ 49 ],
   alphaCSR[ 90 ][ 50 ],
   alphaCSR[ 90 ][ 51 ],
   alphaCSR[ 90 ][ 52 ],
   alphaCSR[ 90 ][ 53 ],
   alphaCSR[ 90 ][ 54 ],
   alphaCSR[ 90 ][ 55 ],
   alphaCSR[ 90 ][ 56 ],
   alphaCSR[ 90 ][ 57 ],
   alphaCSR[ 90 ][ 58 ],
   alphaCSR[ 90 ][ 59 ],
   alphaCSR[ 90 ][ 60 ],
   alphaCSR[ 90 ][ 61 ],
   alphaCSR[ 90 ][ 62 ],
   alphaCSR[ 90 ][ 63 ],
   alphaCSR[ 90 ][ 64 ],
   alphaCSR[ 90 ][ 65 ],
   alphaCSR[ 90 ][ 66 ],
   alphaCSR[ 90 ][ 67 ],
   alphaCSR[ 90 ][ 68 ],
   alphaCSR[ 90 ][ 69 ],
   alphaCSR[ 90 ][ 70 ],
   alphaCSR[ 90 ][ 71 ],
   alphaCSR[ 90 ][ 72 ],
   alphaCSR[ 90 ][ 73 ],
   alphaCSR[ 90 ][ 74 ],
   alphaCSR[ 90 ][ 75 ],
   alphaCSR[ 90 ][ 76 ],
   alphaCSR[ 90 ][ 77 ],
   alphaCSR[ 90 ][ 78 ],
   alphaCSR[ 90 ][ 79 ],
   alphaCSR[ 90 ][ 80 ],
   alphaCSR[ 90 ][ 81 ],
   alphaCSR[ 90 ][ 82 ],
   alphaCSR[ 90 ][ 83 ],
   alphaCSR[ 90 ][ 84 ],
   alphaCSR[ 90 ][ 85 ],
   alphaCSR[ 90 ][ 86 ],
   alphaCSR[ 90 ][ 87 ],
   alphaCSR[ 90 ][ 88 ],
   alphaCSR[ 90 ][ 89 ],
   alphaCSR[ 90 ][ 90 ],
   alphaCSR[ 90 ][ 91 ],
   alphaCSR[ 90 ][ 92 ],
   alphaCSR[ 90 ][ 93 ],
   alphaCSR[ 90 ][ 94 ],
   alphaCSR[ 90 ][ 95 ],
   alphaCSR[ 90 ][ 96 ],
   alphaCSR[ 90 ][ 97 ],
   alphaCSR[ 90 ][ 98 ],
   alphaCSR[ 90 ][ 99 ],
   alphaCSR[ 90 ][ 100 ],
   alphaCSR[ 90 ][ 101 ],
   alphaCSR[ 90 ][ 102 ],
   alphaCSR[ 90 ][ 103 ],
   alphaCSR[ 90 ][ 104 ],
   alphaCSR[ 90 ][ 105 ],
   alphaCSR[ 90 ][ 106 ],
   alphaCSR[ 90 ][ 107 ],
   alphaCSR[ 90 ][ 108 ],
   alphaCSR[ 90 ][ 109 ],
   alphaCSR[ 90 ][ 110 ],
   alphaCSR[ 90 ][ 111 ],
   alphaCSR[ 90 ][ 112 ],
   alphaCSR[ 90 ][ 113 ],
   alphaCSR[ 90 ][ 114 ],
   alphaCSR[ 90 ][ 115 ],
   alphaCSR[ 90 ][ 116 ],
   alphaCSR[ 90 ][ 117 ],
   alphaCSR[ 90 ][ 118 ],
   alphaCSR[ 90 ][ 119 ],
   alphaCSR[ 90 ][ 120 ],
   alphaCSR[ 90 ][ 121 ],
   alphaCSR[ 90 ][ 122 ],
   alphaCSR[ 90 ][ 123 ],
   alphaCSR[ 90 ][ 124 ],
   alphaCSR[ 90 ][ 125 ],
   alphaCSR[ 90 ][ 126 ],
   alphaCSR[ 90 ][ 127 ],
   alphaCSR[ 90 ][ 128 ],
   alphaCSR[ 90 ][ 129 ],
   alphaCSR[ 90 ][ 130 ],
   alphaCSR[ 90 ][ 131 ],
   alphaCSR[ 90 ][ 132 ],
   alphaCSR[ 90 ][ 133 ],
   alphaCSR[ 90 ][ 134 ],
   alphaCSR[ 90 ][ 135 ],
   alphaCSR[ 90 ][ 136 ],
   alphaCSR[ 90 ][ 137 ],
   alphaCSR[ 90 ][ 138 ],
   alphaCSR[ 90 ][ 139 ],
   alphaCSR[ 90 ][ 140 ],
   alphaCSR[ 90 ][ 141 ],
   alphaCSR[ 90 ][ 142 ],
   alphaCSR[ 90 ][ 143 ],
   alphaCSR[ 90 ][ 144 ],
   alphaCSR[ 90 ][ 145 ],
   alphaCSR[ 90 ][ 146 ],
   alphaCSR[ 90 ][ 147 ],
   alphaCSR[ 90 ][ 148 ],
   alphaCSR[ 90 ][ 149 ],
   alphaCSR[ 90 ][ 150 ],
   alphaCSR[ 90 ][ 151 ],
   alphaCSR[ 90 ][ 152 ],
   alphaCSR[ 90 ][ 153 ],
   alphaCSR[ 90 ][ 154 ],
   alphaCSR[ 90 ][ 155 ],
   alphaCSR[ 90 ][ 156 ],
   alphaCSR[ 90 ][ 157 ],
   alphaCSR[ 90 ][ 158 ],
   alphaCSR[ 90 ][ 159 ],
   alphaCSR[ 90 ][ 160 ],
   alphaCSR[ 90 ][ 161 ],
   alphaCSR[ 90 ][ 162 ],
   alphaCSR[ 90 ][ 163 ],
   alphaCSR[ 90 ][ 164 ],
   alphaCSR[ 90 ][ 165 ],
   alphaCSR[ 90 ][ 166 ],
   alphaCSR[ 90 ][ 167 ],
   alphaCSR[ 90 ][ 168 ],
   alphaCSR[ 90 ][ 169 ],
   alphaCSR[ 90 ][ 170 ],
   alphaCSR[ 90 ][ 171 ],
   alphaCSR[ 90 ][ 172 ],
   alphaCSR[ 90 ][ 173 ],
   alphaCSR[ 90 ][ 174 ],
   alphaCSR[ 90 ][ 175 ],
   alphaCSR[ 90 ][ 176 ],
   alphaCSR[ 90 ][ 177 ],
   alphaCSR[ 90 ][ 178 ],
   alphaCSR[ 90 ][ 179 ],
   alphaCSR[ 90 ][ 180 ],
   alphaCSR[ 90 ][ 181 ],
   alphaCSR[ 90 ][ 182 ],
   alphaCSR[ 90 ][ 183 ],
   alphaCSR[ 90 ][ 184 ],
   alphaCSR[ 90 ][ 185 ],
   alphaCSR[ 90 ][ 186 ],
   alphaCSR[ 90 ][ 187 ],
   alphaCSR[ 90 ][ 188 ],
   alphaCSR[ 90 ][ 189 ],
   alphaCSR[ 90 ][ 190 ],
   alphaCSR[ 90 ][ 191 ],
   alphaCSR[ 90 ][ 192 ],
   alphaCSR[ 90 ][ 193 ],
   alphaCSR[ 90 ][ 194 ],
   alphaCSR[ 90 ][ 195 ],
   alphaCSR[ 90 ][ 196 ],
   alphaCSR[ 90 ][ 197 ],
   alphaCSR[ 90 ][ 198 ],
   alphaCSR[ 90 ][ 199 ],
   alphaCSR[ 90 ][ 200 ],
   alphaCSR[ 90 ][ 201 ],
   alphaCSR[ 90 ][ 202 ],
   alphaCSR[ 90 ][ 203 ],
   alphaCSR[ 90 ][ 204 ],
   alphaCSR[ 90 ][ 205 ],
   alphaCSR[ 90 ][ 206 ],
   alphaCSR[ 90 ][ 207 ],
   alphaCSR[ 90 ][ 208 ],
   alphaCSR[ 90 ][ 209 ],
   alphaCSR[ 90 ][ 210 ],
   alphaCSR[ 90 ][ 211 ],
   alphaCSR[ 90 ][ 212 ],
   alphaCSR[ 90 ][ 213 ],
   alphaCSR[ 90 ][ 214 ],
   alphaCSR[ 90 ][ 215 ],
   alphaCSR[ 90 ][ 216 ],
   alphaCSR[ 90 ][ 217 ],
   alphaCSR[ 90 ][ 218 ],
   alphaCSR[ 90 ][ 219 ],
   alphaCSR[ 90 ][ 220 ],
   alphaCSR[ 90 ][ 221 ],
   alphaCSR[ 90 ][ 222 ],
   alphaCSR[ 90 ][ 223 ],
   alphaCSR[ 90 ][ 224 ],
   alphaCSR[ 90 ][ 225 ],
   alphaCSR[ 90 ][ 226 ],
   alphaCSR[ 90 ][ 227 ],
   alphaCSR[ 90 ][ 228 ],
   alphaCSR[ 90 ][ 229 ],
   alphaCSR[ 90 ][ 230 ],
   alphaCSR[ 90 ][ 231 ],
   alphaCSR[ 90 ][ 232 ],
   alphaCSR[ 90 ][ 233 ],
   alphaCSR[ 90 ][ 234 ],
   alphaCSR[ 90 ][ 235 ],
   alphaCSR[ 90 ][ 236 ],
   alphaCSR[ 90 ][ 237 ],
   alphaCSR[ 90 ][ 238 ],
   alphaCSR[ 90 ][ 239 ],
   alphaCSR[ 90 ][ 240 ],
   alphaCSR[ 90 ][ 241 ],
   alphaCSR[ 90 ][ 242 ],
   alphaCSR[ 90 ][ 243 ],
   alphaCSR[ 90 ][ 244 ],
   alphaCSR[ 90 ][ 245 ],
   alphaCSR[ 90 ][ 246 ],
   alphaCSR[ 90 ][ 247 ],
   alphaCSR[ 90 ][ 248 ],
   alphaCSR[ 90 ][ 249 ],
   alphaCSR[ 90 ][ 250 ],
   alphaCSR[ 90 ][ 251 ],
   alphaCSR[ 90 ][ 252 ],
   alphaCSR[ 90 ][ 253 ],
   alphaCSR[ 90 ][ 254 ],
   alphaCSR[ 90 ][ 255 ],
   alphaCSR[ 90 ][ 256 ],
   alphaCSR[ 90 ][ 257 ],
   alphaCSR[ 90 ][ 258 ],
   alphaCSR[ 90 ][ 259 ],
   alphaCSR[ 90 ][ 260 ],
   alphaCSR[ 90 ][ 261 ],
   alphaCSR[ 90 ][ 262 ],
   alphaCSR[ 90 ][ 263 ],
   alphaCSR[ 90 ][ 264 ],
   alphaCSR[ 90 ][ 265 ],
   alphaCSR[ 90 ][ 266 ],
   alphaCSR[ 90 ][ 267 ],
   alphaCSR[ 90 ][ 268 ],
   alphaCSR[ 90 ][ 269 ],
   alphaCSR[ 90 ][ 270 ],
   alphaCSR[ 90 ][ 271 ],
   alphaCSR[ 90 ][ 272 ],
   alphaCSR[ 90 ][ 273 ],
   alphaCSR[ 90 ][ 274 ],
   alphaCSR[ 90 ][ 275 ],
   alphaCSR[ 90 ][ 276 ],
   alphaCSR[ 90 ][ 277 ],
   alphaCSR[ 90 ][ 278 ],
   alphaCSR[ 90 ][ 279 ],
   alphaCSR[ 90 ][ 280 ],
   alphaCSR[ 90 ][ 281 ],
   alphaCSR[ 90 ][ 282 ],
   alphaCSR[ 90 ][ 283 ],
   alphaCSR[ 90 ][ 284 ],
   alphaCSR[ 90 ][ 285 ],
   alphaCSR[ 90 ][ 286 ],
   alphaCSR[ 90 ][ 287 ],
   alphaCSR[ 90 ][ 288 ],
   alphaCSR[ 90 ][ 289 ],
   alphaCSR[ 90 ][ 290 ],
   alphaCSR[ 90 ][ 291 ],
   alphaCSR[ 90 ][ 292 ],
   alphaCSR[ 90 ][ 293 ],
   alphaCSR[ 90 ][ 294 ],
   alphaCSR[ 90 ][ 295 ],
   alphaCSR[ 90 ][ 296 ],
   alphaCSR[ 90 ][ 297 ],
   alphaCSR[ 90 ][ 298 ],
   alphaCSR[ 90 ][ 299 ],
   alphaCSR[ 90 ][ 300 ],
   alphaCSR[ 90 ][ 301 ],
   alphaCSR[ 90 ][ 302 ],
   alphaCSR[ 90 ][ 303 ],
   alphaCSR[ 90 ][ 304 ],
   alphaCSR[ 90 ][ 305 ],
   alphaCSR[ 90 ][ 306 ],
   alphaCSR[ 90 ][ 307 ],
   alphaCSR[ 90 ][ 308 ],
   alphaCSR[ 90 ][ 309 ],
   alphaCSR[ 90 ][ 310 ],
   alphaCSR[ 90 ][ 311 ],
   alphaCSR[ 90 ][ 312 ],
   alphaCSR[ 90 ][ 313 ],
   alphaCSR[ 90 ][ 314 ],
   alphaCSR[ 90 ][ 315 ],
   alphaCSR[ 90 ][ 316 ],
   alphaCSR[ 90 ][ 317 ],
   alphaCSR[ 90 ][ 318 ],
   alphaCSR[ 90 ][ 319 ],
   alphaCSR[ 90 ][ 320 ],
   alphaCSR[ 90 ][ 321 ],
   alphaCSR[ 90 ][ 322 ],
   alphaCSR[ 90 ][ 323 ],
   alphaCSR[ 90 ][ 324 ],
   alphaCSR[ 90 ][ 325 ],
   alphaCSR[ 90 ][ 326 ],
   alphaCSR[ 90 ][ 327 ],
   alphaCSR[ 90 ][ 328 ],
   alphaCSR[ 90 ][ 329 ],
   alphaCSR[ 90 ][ 330 ],
   alphaCSR[ 90 ][ 331 ],
   alphaCSR[ 90 ][ 332 ],
   alphaCSR[ 90 ][ 333 ],
   alphaCSR[ 90 ][ 334 ],
   alphaCSR[ 90 ][ 335 ],
   alphaCSR[ 90 ][ 336 ],
   alphaCSR[ 90 ][ 337 ],
   alphaCSR[ 90 ][ 338 ],
   alphaCSR[ 90 ][ 339 ],
   alphaCSR[ 90 ][ 340 ],
   alphaCSR[ 90 ][ 341 ],
   alphaCSR[ 90 ][ 342 ],
   alphaCSR[ 90 ][ 343 ],
   alphaCSR[ 90 ][ 344 ],
   alphaCSR[ 90 ][ 345 ],
   alphaCSR[ 90 ][ 346 ],
   alphaCSR[ 90 ][ 347 ],
   alphaCSR[ 90 ][ 348 ],
   alphaCSR[ 90 ][ 349 ],
   alphaCSR[ 90 ][ 350 ],
   alphaCSR[ 90 ][ 351 ],
   alphaCSR[ 90 ][ 352 ],
   alphaCSR[ 90 ][ 353 ],
   alphaCSR[ 90 ][ 354 ],
   alphaCSR[ 90 ][ 355 ],
   alphaCSR[ 90 ][ 356 ],
   alphaCSR[ 90 ][ 357 ],
   alphaCSR[ 90 ][ 358 ],
   alphaCSR[ 90 ][ 359 ],
   alphaCSR[ 90 ][ 360 ],
   alphaCSR[ 90 ][ 361 ],
   alphaCSR[ 90 ][ 362 ],
   alphaCSR[ 90 ][ 363 ],
   alphaCSR[ 90 ][ 364 ],
   alphaCSR[ 90 ][ 365 ],
   alphaCSR[ 90 ][ 366 ],
   alphaCSR[ 90 ][ 367 ],
   alphaCSR[ 90 ][ 368 ],
   alphaCSR[ 90 ][ 369 ],
   alphaCSR[ 90 ][ 370 ],
   alphaCSR[ 90 ][ 371 ],
   alphaCSR[ 90 ][ 372 ],
   alphaCSR[ 90 ][ 373 ],
   alphaCSR[ 90 ][ 374 ],
   alphaCSR[ 90 ][ 375 ],
   alphaCSR[ 90 ][ 376 ],
   alphaCSR[ 90 ][ 377 ],
   alphaCSR[ 90 ][ 378 ],
   alphaCSR[ 90 ][ 379 ],
   alphaCSR[ 90 ][ 380 ],
   alphaCSR[ 90 ][ 381 ],
   alphaCSR[ 90 ][ 382 ],
   alphaCSR[ 90 ][ 383 ],
   alphaCSR[ 91 ][ 0 ],
   alphaCSR[ 91 ][ 1 ],
   alphaCSR[ 91 ][ 2 ],
   alphaCSR[ 91 ][ 3 ],
   alphaCSR[ 91 ][ 4 ],
   alphaCSR[ 91 ][ 5 ],
   alphaCSR[ 91 ][ 6 ],
   alphaCSR[ 91 ][ 7 ],
   alphaCSR[ 91 ][ 8 ],
   alphaCSR[ 91 ][ 9 ],
   alphaCSR[ 91 ][ 10 ],
   alphaCSR[ 91 ][ 11 ],
   alphaCSR[ 91 ][ 12 ],
   alphaCSR[ 91 ][ 13 ],
   alphaCSR[ 91 ][ 14 ],
   alphaCSR[ 91 ][ 15 ],
   alphaCSR[ 91 ][ 16 ],
   alphaCSR[ 91 ][ 17 ],
   alphaCSR[ 91 ][ 18 ],
   alphaCSR[ 91 ][ 19 ],
   alphaCSR[ 91 ][ 20 ],
   alphaCSR[ 91 ][ 21 ],
   alphaCSR[ 91 ][ 22 ],
   alphaCSR[ 91 ][ 23 ],
   alphaCSR[ 91 ][ 24 ],
   alphaCSR[ 91 ][ 25 ],
   alphaCSR[ 91 ][ 26 ],
   alphaCSR[ 91 ][ 27 ],
   alphaCSR[ 91 ][ 28 ],
   alphaCSR[ 91 ][ 29 ],
   alphaCSR[ 91 ][ 30 ],
   alphaCSR[ 91 ][ 31 ],
   alphaCSR[ 91 ][ 32 ],
   alphaCSR[ 91 ][ 33 ],
   alphaCSR[ 91 ][ 34 ],
   alphaCSR[ 91 ][ 35 ],
   alphaCSR[ 91 ][ 36 ],
   alphaCSR[ 91 ][ 37 ],
   alphaCSR[ 91 ][ 38 ],
   alphaCSR[ 91 ][ 39 ],
   alphaCSR[ 91 ][ 40 ],
   alphaCSR[ 91 ][ 41 ],
   alphaCSR[ 91 ][ 42 ],
   alphaCSR[ 91 ][ 43 ],
   alphaCSR[ 91 ][ 44 ],
   alphaCSR[ 91 ][ 45 ],
   alphaCSR[ 91 ][ 46 ],
   alphaCSR[ 91 ][ 47 ],
   alphaCSR[ 91 ][ 48 ],
   alphaCSR[ 91 ][ 49 ],
   alphaCSR[ 91 ][ 50 ],
   alphaCSR[ 91 ][ 51 ],
   alphaCSR[ 91 ][ 52 ],
   alphaCSR[ 91 ][ 53 ],
   alphaCSR[ 91 ][ 54 ],
   alphaCSR[ 91 ][ 55 ],
   alphaCSR[ 91 ][ 56 ],
   alphaCSR[ 91 ][ 57 ],
   alphaCSR[ 91 ][ 58 ],
   alphaCSR[ 91 ][ 59 ],
   alphaCSR[ 91 ][ 60 ],
   alphaCSR[ 91 ][ 61 ],
   alphaCSR[ 91 ][ 62 ],
   alphaCSR[ 91 ][ 63 ],
   alphaCSR[ 91 ][ 64 ],
   alphaCSR[ 91 ][ 65 ],
   alphaCSR[ 91 ][ 66 ],
   alphaCSR[ 91 ][ 67 ],
   alphaCSR[ 91 ][ 68 ],
   alphaCSR[ 91 ][ 69 ],
   alphaCSR[ 91 ][ 70 ],
   alphaCSR[ 91 ][ 71 ],
   alphaCSR[ 91 ][ 72 ],
   alphaCSR[ 91 ][ 73 ],
   alphaCSR[ 91 ][ 74 ],
   alphaCSR[ 91 ][ 75 ],
   alphaCSR[ 91 ][ 76 ],
   alphaCSR[ 91 ][ 77 ],
   alphaCSR[ 91 ][ 78 ],
   alphaCSR[ 91 ][ 79 ],
   alphaCSR[ 91 ][ 80 ],
   alphaCSR[ 91 ][ 81 ],
   alphaCSR[ 91 ][ 82 ],
   alphaCSR[ 91 ][ 83 ],
   alphaCSR[ 91 ][ 84 ],
   alphaCSR[ 91 ][ 85 ],
   alphaCSR[ 91 ][ 86 ],
   alphaCSR[ 91 ][ 87 ],
   alphaCSR[ 91 ][ 88 ],
   alphaCSR[ 91 ][ 89 ],
   alphaCSR[ 91 ][ 90 ],
   alphaCSR[ 91 ][ 91 ],
   alphaCSR[ 91 ][ 92 ],
   alphaCSR[ 91 ][ 93 ],
   alphaCSR[ 91 ][ 94 ],
   alphaCSR[ 91 ][ 95 ],
   alphaCSR[ 91 ][ 96 ],
   alphaCSR[ 91 ][ 97 ],
   alphaCSR[ 91 ][ 98 ],
   alphaCSR[ 91 ][ 99 ],
   alphaCSR[ 91 ][ 100 ],
   alphaCSR[ 91 ][ 101 ],
   alphaCSR[ 91 ][ 102 ],
   alphaCSR[ 91 ][ 103 ],
   alphaCSR[ 91 ][ 104 ],
   alphaCSR[ 91 ][ 105 ],
   alphaCSR[ 91 ][ 106 ],
   alphaCSR[ 91 ][ 107 ],
   alphaCSR[ 91 ][ 108 ],
   alphaCSR[ 91 ][ 109 ],
   alphaCSR[ 91 ][ 110 ],
   alphaCSR[ 91 ][ 111 ],
   alphaCSR[ 91 ][ 112 ],
   alphaCSR[ 91 ][ 113 ],
   alphaCSR[ 91 ][ 114 ],
   alphaCSR[ 91 ][ 115 ],
   alphaCSR[ 91 ][ 116 ],
   alphaCSR[ 91 ][ 117 ],
   alphaCSR[ 91 ][ 118 ],
   alphaCSR[ 91 ][ 119 ],
   alphaCSR[ 91 ][ 120 ],
   alphaCSR[ 91 ][ 121 ],
   alphaCSR[ 91 ][ 122 ],
   alphaCSR[ 91 ][ 123 ],
   alphaCSR[ 91 ][ 124 ],
   alphaCSR[ 91 ][ 125 ],
   alphaCSR[ 91 ][ 126 ],
   alphaCSR[ 91 ][ 127 ],
   alphaCSR[ 91 ][ 128 ],
   alphaCSR[ 91 ][ 129 ],
   alphaCSR[ 91 ][ 130 ],
   alphaCSR[ 91 ][ 131 ],
   alphaCSR[ 91 ][ 132 ],
   alphaCSR[ 91 ][ 133 ],
   alphaCSR[ 91 ][ 134 ],
   alphaCSR[ 91 ][ 135 ],
   alphaCSR[ 91 ][ 136 ],
   alphaCSR[ 91 ][ 137 ],
   alphaCSR[ 91 ][ 138 ],
   alphaCSR[ 91 ][ 139 ],
   alphaCSR[ 91 ][ 140 ],
   alphaCSR[ 91 ][ 141 ],
   alphaCSR[ 91 ][ 142 ],
   alphaCSR[ 91 ][ 143 ],
   alphaCSR[ 91 ][ 144 ],
   alphaCSR[ 91 ][ 145 ],
   alphaCSR[ 91 ][ 146 ],
   alphaCSR[ 91 ][ 147 ],
   alphaCSR[ 91 ][ 148 ],
   alphaCSR[ 91 ][ 149 ],
   alphaCSR[ 91 ][ 150 ],
   alphaCSR[ 91 ][ 151 ],
   alphaCSR[ 91 ][ 152 ],
   alphaCSR[ 91 ][ 153 ],
   alphaCSR[ 91 ][ 154 ],
   alphaCSR[ 91 ][ 155 ],
   alphaCSR[ 91 ][ 156 ],
   alphaCSR[ 91 ][ 157 ],
   alphaCSR[ 91 ][ 158 ],
   alphaCSR[ 91 ][ 159 ],
   alphaCSR[ 91 ][ 160 ],
   alphaCSR[ 91 ][ 161 ],
   alphaCSR[ 91 ][ 162 ],
   alphaCSR[ 91 ][ 163 ],
   alphaCSR[ 91 ][ 164 ],
   alphaCSR[ 91 ][ 165 ],
   alphaCSR[ 91 ][ 166 ],
   alphaCSR[ 91 ][ 167 ],
   alphaCSR[ 91 ][ 168 ],
   alphaCSR[ 91 ][ 169 ],
   alphaCSR[ 91 ][ 170 ],
   alphaCSR[ 91 ][ 171 ],
   alphaCSR[ 91 ][ 172 ],
   alphaCSR[ 91 ][ 173 ],
   alphaCSR[ 91 ][ 174 ],
   alphaCSR[ 91 ][ 175 ],
   alphaCSR[ 91 ][ 176 ],
   alphaCSR[ 91 ][ 177 ],
   alphaCSR[ 91 ][ 178 ],
   alphaCSR[ 91 ][ 179 ],
   alphaCSR[ 91 ][ 180 ],
   alphaCSR[ 91 ][ 181 ],
   alphaCSR[ 91 ][ 182 ],
   alphaCSR[ 91 ][ 183 ],
   alphaCSR[ 91 ][ 184 ],
   alphaCSR[ 91 ][ 185 ],
   alphaCSR[ 91 ][ 186 ],
   alphaCSR[ 91 ][ 187 ],
   alphaCSR[ 91 ][ 188 ],
   alphaCSR[ 91 ][ 189 ],
   alphaCSR[ 91 ][ 190 ],
   alphaCSR[ 91 ][ 191 ],
   alphaCSR[ 91 ][ 192 ],
   alphaCSR[ 91 ][ 193 ],
   alphaCSR[ 91 ][ 194 ],
   alphaCSR[ 91 ][ 195 ],
   alphaCSR[ 91 ][ 196 ],
   alphaCSR[ 91 ][ 197 ],
   alphaCSR[ 91 ][ 198 ],
   alphaCSR[ 91 ][ 199 ],
   alphaCSR[ 91 ][ 200 ],
   alphaCSR[ 91 ][ 201 ],
   alphaCSR[ 91 ][ 202 ],
   alphaCSR[ 91 ][ 203 ],
   alphaCSR[ 91 ][ 204 ],
   alphaCSR[ 91 ][ 205 ],
   alphaCSR[ 91 ][ 206 ],
   alphaCSR[ 91 ][ 207 ],
   alphaCSR[ 91 ][ 208 ],
   alphaCSR[ 91 ][ 209 ],
   alphaCSR[ 91 ][ 210 ],
   alphaCSR[ 91 ][ 211 ],
   alphaCSR[ 91 ][ 212 ],
   alphaCSR[ 91 ][ 213 ],
   alphaCSR[ 91 ][ 214 ],
   alphaCSR[ 91 ][ 215 ],
   alphaCSR[ 91 ][ 216 ],
   alphaCSR[ 91 ][ 217 ],
   alphaCSR[ 91 ][ 218 ],
   alphaCSR[ 91 ][ 219 ],
   alphaCSR[ 91 ][ 220 ],
   alphaCSR[ 91 ][ 221 ],
   alphaCSR[ 91 ][ 222 ],
   alphaCSR[ 91 ][ 223 ],
   alphaCSR[ 91 ][ 224 ],
   alphaCSR[ 91 ][ 225 ],
   alphaCSR[ 91 ][ 226 ],
   alphaCSR[ 91 ][ 227 ],
   alphaCSR[ 91 ][ 228 ],
   alphaCSR[ 91 ][ 229 ],
   alphaCSR[ 91 ][ 230 ],
   alphaCSR[ 91 ][ 231 ],
   alphaCSR[ 91 ][ 232 ],
   alphaCSR[ 91 ][ 233 ],
   alphaCSR[ 91 ][ 234 ],
   alphaCSR[ 91 ][ 235 ],
   alphaCSR[ 91 ][ 236 ],
   alphaCSR[ 91 ][ 237 ],
   alphaCSR[ 91 ][ 238 ],
   alphaCSR[ 91 ][ 239 ],
   alphaCSR[ 91 ][ 240 ],
   alphaCSR[ 91 ][ 241 ],
   alphaCSR[ 91 ][ 242 ],
   alphaCSR[ 91 ][ 243 ],
   alphaCSR[ 91 ][ 244 ],
   alphaCSR[ 91 ][ 245 ],
   alphaCSR[ 91 ][ 246 ],
   alphaCSR[ 91 ][ 247 ],
   alphaCSR[ 91 ][ 248 ],
   alphaCSR[ 91 ][ 249 ],
   alphaCSR[ 91 ][ 250 ],
   alphaCSR[ 91 ][ 251 ],
   alphaCSR[ 91 ][ 252 ],
   alphaCSR[ 91 ][ 253 ],
   alphaCSR[ 91 ][ 254 ],
   alphaCSR[ 91 ][ 255 ],
   alphaCSR[ 91 ][ 256 ],
   alphaCSR[ 91 ][ 257 ],
   alphaCSR[ 91 ][ 258 ],
   alphaCSR[ 91 ][ 259 ],
   alphaCSR[ 91 ][ 260 ],
   alphaCSR[ 91 ][ 261 ],
   alphaCSR[ 91 ][ 262 ],
   alphaCSR[ 91 ][ 263 ],
   alphaCSR[ 91 ][ 264 ],
   alphaCSR[ 91 ][ 265 ],
   alphaCSR[ 91 ][ 266 ],
   alphaCSR[ 91 ][ 267 ],
   alphaCSR[ 91 ][ 268 ],
   alphaCSR[ 91 ][ 269 ],
   alphaCSR[ 91 ][ 270 ],
   alphaCSR[ 91 ][ 271 ],
   alphaCSR[ 91 ][ 272 ],
   alphaCSR[ 91 ][ 273 ],
   alphaCSR[ 91 ][ 274 ],
   alphaCSR[ 91 ][ 275 ],
   alphaCSR[ 91 ][ 276 ],
   alphaCSR[ 91 ][ 277 ],
   alphaCSR[ 91 ][ 278 ],
   alphaCSR[ 91 ][ 279 ],
   alphaCSR[ 91 ][ 280 ],
   alphaCSR[ 91 ][ 281 ],
   alphaCSR[ 91 ][ 282 ],
   alphaCSR[ 91 ][ 283 ],
   alphaCSR[ 91 ][ 284 ],
   alphaCSR[ 91 ][ 285 ],
   alphaCSR[ 91 ][ 286 ],
   alphaCSR[ 91 ][ 287 ],
   alphaCSR[ 91 ][ 288 ],
   alphaCSR[ 91 ][ 289 ],
   alphaCSR[ 91 ][ 290 ],
   alphaCSR[ 91 ][ 291 ],
   alphaCSR[ 91 ][ 292 ],
   alphaCSR[ 91 ][ 293 ],
   alphaCSR[ 91 ][ 294 ],
   alphaCSR[ 91 ][ 295 ],
   alphaCSR[ 91 ][ 296 ],
   alphaCSR[ 91 ][ 297 ],
   alphaCSR[ 91 ][ 298 ],
   alphaCSR[ 91 ][ 299 ],
   alphaCSR[ 91 ][ 300 ],
   alphaCSR[ 91 ][ 301 ],
   alphaCSR[ 91 ][ 302 ],
   alphaCSR[ 91 ][ 303 ],
   alphaCSR[ 91 ][ 304 ],
   alphaCSR[ 91 ][ 305 ],
   alphaCSR[ 91 ][ 306 ],
   alphaCSR[ 91 ][ 307 ],
   alphaCSR[ 91 ][ 308 ],
   alphaCSR[ 91 ][ 309 ],
   alphaCSR[ 91 ][ 310 ],
   alphaCSR[ 91 ][ 311 ],
   alphaCSR[ 91 ][ 312 ],
   alphaCSR[ 91 ][ 313 ],
   alphaCSR[ 91 ][ 314 ],
   alphaCSR[ 91 ][ 315 ],
   alphaCSR[ 91 ][ 316 ],
   alphaCSR[ 91 ][ 317 ],
   alphaCSR[ 91 ][ 318 ],
   alphaCSR[ 91 ][ 319 ],
   alphaCSR[ 91 ][ 320 ],
   alphaCSR[ 91 ][ 321 ],
   alphaCSR[ 91 ][ 322 ],
   alphaCSR[ 91 ][ 323 ],
   alphaCSR[ 91 ][ 324 ],
   alphaCSR[ 91 ][ 325 ],
   alphaCSR[ 91 ][ 326 ],
   alphaCSR[ 91 ][ 327 ],
   alphaCSR[ 91 ][ 328 ],
   alphaCSR[ 91 ][ 329 ],
   alphaCSR[ 91 ][ 330 ],
   alphaCSR[ 91 ][ 331 ],
   alphaCSR[ 91 ][ 332 ],
   alphaCSR[ 91 ][ 333 ],
   alphaCSR[ 91 ][ 334 ],
   alphaCSR[ 91 ][ 335 ],
   alphaCSR[ 91 ][ 336 ],
   alphaCSR[ 91 ][ 337 ],
   alphaCSR[ 91 ][ 338 ],
   alphaCSR[ 91 ][ 339 ],
   alphaCSR[ 91 ][ 340 ],
   alphaCSR[ 91 ][ 341 ],
   alphaCSR[ 91 ][ 342 ],
   alphaCSR[ 91 ][ 343 ],
   alphaCSR[ 91 ][ 344 ],
   alphaCSR[ 91 ][ 345 ],
   alphaCSR[ 91 ][ 346 ],
   alphaCSR[ 91 ][ 347 ],
   alphaCSR[ 91 ][ 348 ],
   alphaCSR[ 91 ][ 349 ],
   alphaCSR[ 91 ][ 350 ],
   alphaCSR[ 91 ][ 351 ],
   alphaCSR[ 91 ][ 352 ],
   alphaCSR[ 91 ][ 353 ],
   alphaCSR[ 91 ][ 354 ],
   alphaCSR[ 91 ][ 355 ],
   alphaCSR[ 91 ][ 356 ],
   alphaCSR[ 91 ][ 357 ],
   alphaCSR[ 91 ][ 358 ],
   alphaCSR[ 91 ][ 359 ],
   alphaCSR[ 91 ][ 360 ],
   alphaCSR[ 91 ][ 361 ],
   alphaCSR[ 91 ][ 362 ],
   alphaCSR[ 91 ][ 363 ],
   alphaCSR[ 91 ][ 364 ],
   alphaCSR[ 91 ][ 365 ],
   alphaCSR[ 91 ][ 366 ],
   alphaCSR[ 91 ][ 367 ],
   alphaCSR[ 91 ][ 368 ],
   alphaCSR[ 91 ][ 369 ],
   alphaCSR[ 91 ][ 370 ],
   alphaCSR[ 91 ][ 371 ],
   alphaCSR[ 91 ][ 372 ],
   alphaCSR[ 91 ][ 373 ],
   alphaCSR[ 91 ][ 374 ],
   alphaCSR[ 91 ][ 375 ],
   alphaCSR[ 91 ][ 376 ],
   alphaCSR[ 91 ][ 377 ],
   alphaCSR[ 91 ][ 378 ],
   alphaCSR[ 91 ][ 379 ],
   alphaCSR[ 91 ][ 380 ],
   alphaCSR[ 91 ][ 381 ],
   alphaCSR[ 91 ][ 382 ],
   alphaCSR[ 91 ][ 383 ],
   alphaCSR[ 92 ][ 0 ],
   alphaCSR[ 92 ][ 1 ],
   alphaCSR[ 92 ][ 2 ],
   alphaCSR[ 92 ][ 3 ],
   alphaCSR[ 92 ][ 4 ],
   alphaCSR[ 92 ][ 5 ],
   alphaCSR[ 92 ][ 6 ],
   alphaCSR[ 92 ][ 7 ],
   alphaCSR[ 92 ][ 8 ],
   alphaCSR[ 92 ][ 9 ],
   alphaCSR[ 92 ][ 10 ],
   alphaCSR[ 92 ][ 11 ],
   alphaCSR[ 92 ][ 12 ],
   alphaCSR[ 92 ][ 13 ],
   alphaCSR[ 92 ][ 14 ],
   alphaCSR[ 92 ][ 15 ],
   alphaCSR[ 92 ][ 16 ],
   alphaCSR[ 92 ][ 17 ],
   alphaCSR[ 92 ][ 18 ],
   alphaCSR[ 92 ][ 19 ],
   alphaCSR[ 92 ][ 20 ],
   alphaCSR[ 92 ][ 21 ],
   alphaCSR[ 92 ][ 22 ],
   alphaCSR[ 92 ][ 23 ],
   alphaCSR[ 92 ][ 24 ],
   alphaCSR[ 92 ][ 25 ],
   alphaCSR[ 92 ][ 26 ],
   alphaCSR[ 92 ][ 27 ],
   alphaCSR[ 92 ][ 28 ],
   alphaCSR[ 92 ][ 29 ],
   alphaCSR[ 92 ][ 30 ],
   alphaCSR[ 92 ][ 31 ],
   alphaCSR[ 92 ][ 32 ],
   alphaCSR[ 92 ][ 33 ],
   alphaCSR[ 92 ][ 34 ],
   alphaCSR[ 92 ][ 35 ],
   alphaCSR[ 92 ][ 36 ],
   alphaCSR[ 92 ][ 37 ],
   alphaCSR[ 92 ][ 38 ],
   alphaCSR[ 92 ][ 39 ],
   alphaCSR[ 92 ][ 40 ],
   alphaCSR[ 92 ][ 41 ],
   alphaCSR[ 92 ][ 42 ],
   alphaCSR[ 92 ][ 43 ],
   alphaCSR[ 92 ][ 44 ],
   alphaCSR[ 92 ][ 45 ],
   alphaCSR[ 92 ][ 46 ],
   alphaCSR[ 92 ][ 47 ],
   alphaCSR[ 92 ][ 48 ],
   alphaCSR[ 92 ][ 49 ],
   alphaCSR[ 92 ][ 50 ],
   alphaCSR[ 92 ][ 51 ],
   alphaCSR[ 92 ][ 52 ],
   alphaCSR[ 92 ][ 53 ],
   alphaCSR[ 92 ][ 54 ],
   alphaCSR[ 92 ][ 55 ],
   alphaCSR[ 92 ][ 56 ],
   alphaCSR[ 92 ][ 57 ],
   alphaCSR[ 92 ][ 58 ],
   alphaCSR[ 92 ][ 59 ],
   alphaCSR[ 92 ][ 60 ],
   alphaCSR[ 92 ][ 61 ],
   alphaCSR[ 92 ][ 62 ],
   alphaCSR[ 92 ][ 63 ],
   alphaCSR[ 92 ][ 64 ],
   alphaCSR[ 92 ][ 65 ],
   alphaCSR[ 92 ][ 66 ],
   alphaCSR[ 92 ][ 67 ],
   alphaCSR[ 92 ][ 68 ],
   alphaCSR[ 92 ][ 69 ],
   alphaCSR[ 92 ][ 70 ],
   alphaCSR[ 92 ][ 71 ],
   alphaCSR[ 92 ][ 72 ],
   alphaCSR[ 92 ][ 73 ],
   alphaCSR[ 92 ][ 74 ],
   alphaCSR[ 92 ][ 75 ],
   alphaCSR[ 92 ][ 76 ],
   alphaCSR[ 92 ][ 77 ],
   alphaCSR[ 92 ][ 78 ],
   alphaCSR[ 92 ][ 79 ],
   alphaCSR[ 92 ][ 80 ],
   alphaCSR[ 92 ][ 81 ],
   alphaCSR[ 92 ][ 82 ],
   alphaCSR[ 92 ][ 83 ],
   alphaCSR[ 92 ][ 84 ],
   alphaCSR[ 92 ][ 85 ],
   alphaCSR[ 92 ][ 86 ],
   alphaCSR[ 92 ][ 87 ],
   alphaCSR[ 92 ][ 88 ],
   alphaCSR[ 92 ][ 89 ],
   alphaCSR[ 92 ][ 90 ],
   alphaCSR[ 92 ][ 91 ],
   alphaCSR[ 92 ][ 92 ],
   alphaCSR[ 92 ][ 93 ],
   alphaCSR[ 92 ][ 94 ],
   alphaCSR[ 92 ][ 95 ],
   alphaCSR[ 92 ][ 96 ],
   alphaCSR[ 92 ][ 97 ],
   alphaCSR[ 92 ][ 98 ],
   alphaCSR[ 92 ][ 99 ],
   alphaCSR[ 92 ][ 100 ],
   alphaCSR[ 92 ][ 101 ],
   alphaCSR[ 92 ][ 102 ],
   alphaCSR[ 92 ][ 103 ],
   alphaCSR[ 92 ][ 104 ],
   alphaCSR[ 92 ][ 105 ],
   alphaCSR[ 92 ][ 106 ],
   alphaCSR[ 92 ][ 107 ],
   alphaCSR[ 92 ][ 108 ],
   alphaCSR[ 92 ][ 109 ],
   alphaCSR[ 92 ][ 110 ],
   alphaCSR[ 92 ][ 111 ],
   alphaCSR[ 92 ][ 112 ],
   alphaCSR[ 92 ][ 113 ],
   alphaCSR[ 92 ][ 114 ],
   alphaCSR[ 92 ][ 115 ],
   alphaCSR[ 92 ][ 116 ],
   alphaCSR[ 92 ][ 117 ],
   alphaCSR[ 92 ][ 118 ],
   alphaCSR[ 92 ][ 119 ],
   alphaCSR[ 92 ][ 120 ],
   alphaCSR[ 92 ][ 121 ],
   alphaCSR[ 92 ][ 122 ],
   alphaCSR[ 92 ][ 123 ],
   alphaCSR[ 92 ][ 124 ],
   alphaCSR[ 92 ][ 125 ],
   alphaCSR[ 92 ][ 126 ],
   alphaCSR[ 92 ][ 127 ],
   alphaCSR[ 92 ][ 128 ],
   alphaCSR[ 92 ][ 129 ],
   alphaCSR[ 92 ][ 130 ],
   alphaCSR[ 92 ][ 131 ],
   alphaCSR[ 92 ][ 132 ],
   alphaCSR[ 92 ][ 133 ],
   alphaCSR[ 92 ][ 134 ],
   alphaCSR[ 92 ][ 135 ],
   alphaCSR[ 92 ][ 136 ],
   alphaCSR[ 92 ][ 137 ],
   alphaCSR[ 92 ][ 138 ],
   alphaCSR[ 92 ][ 139 ],
   alphaCSR[ 92 ][ 140 ],
   alphaCSR[ 92 ][ 141 ],
   alphaCSR[ 92 ][ 142 ],
   alphaCSR[ 92 ][ 143 ],
   alphaCSR[ 92 ][ 144 ],
   alphaCSR[ 92 ][ 145 ],
   alphaCSR[ 92 ][ 146 ],
   alphaCSR[ 92 ][ 147 ],
   alphaCSR[ 92 ][ 148 ],
   alphaCSR[ 92 ][ 149 ],
   alphaCSR[ 92 ][ 150 ],
   alphaCSR[ 92 ][ 151 ],
   alphaCSR[ 92 ][ 152 ],
   alphaCSR[ 92 ][ 153 ],
   alphaCSR[ 92 ][ 154 ],
   alphaCSR[ 92 ][ 155 ],
   alphaCSR[ 92 ][ 156 ],
   alphaCSR[ 92 ][ 157 ],
   alphaCSR[ 92 ][ 158 ],
   alphaCSR[ 92 ][ 159 ],
   alphaCSR[ 92 ][ 160 ],
   alphaCSR[ 92 ][ 161 ],
   alphaCSR[ 92 ][ 162 ],
   alphaCSR[ 92 ][ 163 ],
   alphaCSR[ 92 ][ 164 ],
   alphaCSR[ 92 ][ 165 ],
   alphaCSR[ 92 ][ 166 ],
   alphaCSR[ 92 ][ 167 ],
   alphaCSR[ 92 ][ 168 ],
   alphaCSR[ 92 ][ 169 ],
   alphaCSR[ 92 ][ 170 ],
   alphaCSR[ 92 ][ 171 ],
   alphaCSR[ 92 ][ 172 ],
   alphaCSR[ 92 ][ 173 ],
   alphaCSR[ 92 ][ 174 ],
   alphaCSR[ 92 ][ 175 ],
   alphaCSR[ 92 ][ 176 ],
   alphaCSR[ 92 ][ 177 ],
   alphaCSR[ 92 ][ 178 ],
   alphaCSR[ 92 ][ 179 ],
   alphaCSR[ 92 ][ 180 ],
   alphaCSR[ 92 ][ 181 ],
   alphaCSR[ 92 ][ 182 ],
   alphaCSR[ 92 ][ 183 ],
   alphaCSR[ 92 ][ 184 ],
   alphaCSR[ 92 ][ 185 ],
   alphaCSR[ 92 ][ 186 ],
   alphaCSR[ 92 ][ 187 ],
   alphaCSR[ 92 ][ 188 ],
   alphaCSR[ 92 ][ 189 ],
   alphaCSR[ 92 ][ 190 ],
   alphaCSR[ 92 ][ 191 ],
   alphaCSR[ 92 ][ 192 ],
   alphaCSR[ 92 ][ 193 ],
   alphaCSR[ 92 ][ 194 ],
   alphaCSR[ 92 ][ 195 ],
   alphaCSR[ 92 ][ 196 ],
   alphaCSR[ 92 ][ 197 ],
   alphaCSR[ 92 ][ 198 ],
   alphaCSR[ 92 ][ 199 ],
   alphaCSR[ 92 ][ 200 ],
   alphaCSR[ 92 ][ 201 ],
   alphaCSR[ 92 ][ 202 ],
   alphaCSR[ 92 ][ 203 ],
   alphaCSR[ 92 ][ 204 ],
   alphaCSR[ 92 ][ 205 ],
   alphaCSR[ 92 ][ 206 ],
   alphaCSR[ 92 ][ 207 ],
   alphaCSR[ 92 ][ 208 ],
   alphaCSR[ 92 ][ 209 ],
   alphaCSR[ 92 ][ 210 ],
   alphaCSR[ 92 ][ 211 ],
   alphaCSR[ 92 ][ 212 ],
   alphaCSR[ 92 ][ 213 ],
   alphaCSR[ 92 ][ 214 ],
   alphaCSR[ 92 ][ 215 ],
   alphaCSR[ 92 ][ 216 ],
   alphaCSR[ 92 ][ 217 ],
   alphaCSR[ 92 ][ 218 ],
   alphaCSR[ 92 ][ 219 ],
   alphaCSR[ 92 ][ 220 ],
   alphaCSR[ 92 ][ 221 ],
   alphaCSR[ 92 ][ 222 ],
   alphaCSR[ 92 ][ 223 ],
   alphaCSR[ 92 ][ 224 ],
   alphaCSR[ 92 ][ 225 ],
   alphaCSR[ 92 ][ 226 ],
   alphaCSR[ 92 ][ 227 ],
   alphaCSR[ 92 ][ 228 ],
   alphaCSR[ 92 ][ 229 ],
   alphaCSR[ 92 ][ 230 ],
   alphaCSR[ 92 ][ 231 ],
   alphaCSR[ 92 ][ 232 ],
   alphaCSR[ 92 ][ 233 ],
   alphaCSR[ 92 ][ 234 ],
   alphaCSR[ 92 ][ 235 ],
   alphaCSR[ 92 ][ 236 ],
   alphaCSR[ 92 ][ 237 ],
   alphaCSR[ 92 ][ 238 ],
   alphaCSR[ 92 ][ 239 ],
   alphaCSR[ 92 ][ 240 ],
   alphaCSR[ 92 ][ 241 ],
   alphaCSR[ 92 ][ 242 ],
   alphaCSR[ 92 ][ 243 ],
   alphaCSR[ 92 ][ 244 ],
   alphaCSR[ 92 ][ 245 ],
   alphaCSR[ 92 ][ 246 ],
   alphaCSR[ 92 ][ 247 ],
   alphaCSR[ 92 ][ 248 ],
   alphaCSR[ 92 ][ 249 ],
   alphaCSR[ 92 ][ 250 ],
   alphaCSR[ 92 ][ 251 ],
   alphaCSR[ 92 ][ 252 ],
   alphaCSR[ 92 ][ 253 ],
   alphaCSR[ 92 ][ 254 ],
   alphaCSR[ 92 ][ 255 ],
   alphaCSR[ 92 ][ 256 ],
   alphaCSR[ 92 ][ 257 ],
   alphaCSR[ 92 ][ 258 ],
   alphaCSR[ 92 ][ 259 ],
   alphaCSR[ 92 ][ 260 ],
   alphaCSR[ 92 ][ 261 ],
   alphaCSR[ 92 ][ 262 ],
   alphaCSR[ 92 ][ 263 ],
   alphaCSR[ 92 ][ 264 ],
   alphaCSR[ 92 ][ 265 ],
   alphaCSR[ 92 ][ 266 ],
   alphaCSR[ 92 ][ 267 ],
   alphaCSR[ 92 ][ 268 ],
   alphaCSR[ 92 ][ 269 ],
   alphaCSR[ 92 ][ 270 ],
   alphaCSR[ 92 ][ 271 ],
   alphaCSR[ 92 ][ 272 ],
   alphaCSR[ 92 ][ 273 ],
   alphaCSR[ 92 ][ 274 ],
   alphaCSR[ 92 ][ 275 ],
   alphaCSR[ 92 ][ 276 ],
   alphaCSR[ 92 ][ 277 ],
   alphaCSR[ 92 ][ 278 ],
   alphaCSR[ 92 ][ 279 ],
   alphaCSR[ 92 ][ 280 ],
   alphaCSR[ 92 ][ 281 ],
   alphaCSR[ 92 ][ 282 ],
   alphaCSR[ 92 ][ 283 ],
   alphaCSR[ 92 ][ 284 ],
   alphaCSR[ 92 ][ 285 ],
   alphaCSR[ 92 ][ 286 ],
   alphaCSR[ 92 ][ 287 ],
   alphaCSR[ 92 ][ 288 ],
   alphaCSR[ 92 ][ 289 ],
   alphaCSR[ 92 ][ 290 ],
   alphaCSR[ 92 ][ 291 ],
   alphaCSR[ 92 ][ 292 ],
   alphaCSR[ 92 ][ 293 ],
   alphaCSR[ 92 ][ 294 ],
   alphaCSR[ 92 ][ 295 ],
   alphaCSR[ 92 ][ 296 ],
   alphaCSR[ 92 ][ 297 ],
   alphaCSR[ 92 ][ 298 ],
   alphaCSR[ 92 ][ 299 ],
   alphaCSR[ 92 ][ 300 ],
   alphaCSR[ 92 ][ 301 ],
   alphaCSR[ 92 ][ 302 ],
   alphaCSR[ 92 ][ 303 ],
   alphaCSR[ 92 ][ 304 ],
   alphaCSR[ 92 ][ 305 ],
   alphaCSR[ 92 ][ 306 ],
   alphaCSR[ 92 ][ 307 ],
   alphaCSR[ 92 ][ 308 ],
   alphaCSR[ 92 ][ 309 ],
   alphaCSR[ 92 ][ 310 ],
   alphaCSR[ 92 ][ 311 ],
   alphaCSR[ 92 ][ 312 ],
   alphaCSR[ 92 ][ 313 ],
   alphaCSR[ 92 ][ 314 ],
   alphaCSR[ 92 ][ 315 ],
   alphaCSR[ 92 ][ 316 ],
   alphaCSR[ 92 ][ 317 ],
   alphaCSR[ 92 ][ 318 ],
   alphaCSR[ 92 ][ 319 ],
   alphaCSR[ 92 ][ 320 ],
   alphaCSR[ 92 ][ 321 ],
   alphaCSR[ 92 ][ 322 ],
   alphaCSR[ 92 ][ 323 ],
   alphaCSR[ 92 ][ 324 ],
   alphaCSR[ 92 ][ 325 ],
   alphaCSR[ 92 ][ 326 ],
   alphaCSR[ 92 ][ 327 ],
   alphaCSR[ 92 ][ 328 ],
   alphaCSR[ 92 ][ 329 ],
   alphaCSR[ 92 ][ 330 ],
   alphaCSR[ 92 ][ 331 ],
   alphaCSR[ 92 ][ 332 ],
   alphaCSR[ 92 ][ 333 ],
   alphaCSR[ 92 ][ 334 ],
   alphaCSR[ 92 ][ 335 ],
   alphaCSR[ 92 ][ 336 ],
   alphaCSR[ 92 ][ 337 ],
   alphaCSR[ 92 ][ 338 ],
   alphaCSR[ 92 ][ 339 ],
   alphaCSR[ 92 ][ 340 ],
   alphaCSR[ 92 ][ 341 ],
   alphaCSR[ 92 ][ 342 ],
   alphaCSR[ 92 ][ 343 ],
   alphaCSR[ 92 ][ 344 ],
   alphaCSR[ 92 ][ 345 ],
   alphaCSR[ 92 ][ 346 ],
   alphaCSR[ 92 ][ 347 ],
   alphaCSR[ 92 ][ 348 ],
   alphaCSR[ 92 ][ 349 ],
   alphaCSR[ 92 ][ 350 ],
   alphaCSR[ 92 ][ 351 ],
   alphaCSR[ 92 ][ 352 ],
   alphaCSR[ 92 ][ 353 ],
   alphaCSR[ 92 ][ 354 ],
   alphaCSR[ 92 ][ 355 ],
   alphaCSR[ 92 ][ 356 ],
   alphaCSR[ 92 ][ 357 ],
   alphaCSR[ 92 ][ 358 ],
   alphaCSR[ 92 ][ 359 ],
   alphaCSR[ 92 ][ 360 ],
   alphaCSR[ 92 ][ 361 ],
   alphaCSR[ 92 ][ 362 ],
   alphaCSR[ 92 ][ 363 ],
   alphaCSR[ 92 ][ 364 ],
   alphaCSR[ 92 ][ 365 ],
   alphaCSR[ 92 ][ 366 ],
   alphaCSR[ 92 ][ 367 ],
   alphaCSR[ 92 ][ 368 ],
   alphaCSR[ 92 ][ 369 ],
   alphaCSR[ 92 ][ 370 ],
   alphaCSR[ 92 ][ 371 ],
   alphaCSR[ 92 ][ 372 ],
   alphaCSR[ 92 ][ 373 ],
   alphaCSR[ 92 ][ 374 ],
   alphaCSR[ 92 ][ 375 ],
   alphaCSR[ 92 ][ 376 ],
   alphaCSR[ 92 ][ 377 ],
   alphaCSR[ 92 ][ 378 ],
   alphaCSR[ 92 ][ 379 ],
   alphaCSR[ 92 ][ 380 ],
   alphaCSR[ 92 ][ 381 ],
   alphaCSR[ 92 ][ 382 ],
   alphaCSR[ 92 ][ 383 ],
   alphaCSR[ 93 ][ 0 ],
   alphaCSR[ 93 ][ 1 ],
   alphaCSR[ 93 ][ 2 ],
   alphaCSR[ 93 ][ 3 ],
   alphaCSR[ 93 ][ 4 ],
   alphaCSR[ 93 ][ 5 ],
   alphaCSR[ 93 ][ 6 ],
   alphaCSR[ 93 ][ 7 ],
   alphaCSR[ 93 ][ 8 ],
   alphaCSR[ 93 ][ 9 ],
   alphaCSR[ 93 ][ 10 ],
   alphaCSR[ 93 ][ 11 ],
   alphaCSR[ 93 ][ 12 ],
   alphaCSR[ 93 ][ 13 ],
   alphaCSR[ 93 ][ 14 ],
   alphaCSR[ 93 ][ 15 ],
   alphaCSR[ 93 ][ 16 ],
   alphaCSR[ 93 ][ 17 ],
   alphaCSR[ 93 ][ 18 ],
   alphaCSR[ 93 ][ 19 ],
   alphaCSR[ 93 ][ 20 ],
   alphaCSR[ 93 ][ 21 ],
   alphaCSR[ 93 ][ 22 ],
   alphaCSR[ 93 ][ 23 ],
   alphaCSR[ 93 ][ 24 ],
   alphaCSR[ 93 ][ 25 ],
   alphaCSR[ 93 ][ 26 ],
   alphaCSR[ 93 ][ 27 ],
   alphaCSR[ 93 ][ 28 ],
   alphaCSR[ 93 ][ 29 ],
   alphaCSR[ 93 ][ 30 ],
   alphaCSR[ 93 ][ 31 ],
   alphaCSR[ 93 ][ 32 ],
   alphaCSR[ 93 ][ 33 ],
   alphaCSR[ 93 ][ 34 ],
   alphaCSR[ 93 ][ 35 ],
   alphaCSR[ 93 ][ 36 ],
   alphaCSR[ 93 ][ 37 ],
   alphaCSR[ 93 ][ 38 ],
   alphaCSR[ 93 ][ 39 ],
   alphaCSR[ 93 ][ 40 ],
   alphaCSR[ 93 ][ 41 ],
   alphaCSR[ 93 ][ 42 ],
   alphaCSR[ 93 ][ 43 ],
   alphaCSR[ 93 ][ 44 ],
   alphaCSR[ 93 ][ 45 ],
   alphaCSR[ 93 ][ 46 ],
   alphaCSR[ 93 ][ 47 ],
   alphaCSR[ 93 ][ 48 ],
   alphaCSR[ 93 ][ 49 ],
   alphaCSR[ 93 ][ 50 ],
   alphaCSR[ 93 ][ 51 ],
   alphaCSR[ 93 ][ 52 ],
   alphaCSR[ 93 ][ 53 ],
   alphaCSR[ 93 ][ 54 ],
   alphaCSR[ 93 ][ 55 ],
   alphaCSR[ 93 ][ 56 ],
   alphaCSR[ 93 ][ 57 ],
   alphaCSR[ 93 ][ 58 ],
   alphaCSR[ 93 ][ 59 ],
   alphaCSR[ 93 ][ 60 ],
   alphaCSR[ 93 ][ 61 ],
   alphaCSR[ 93 ][ 62 ],
   alphaCSR[ 93 ][ 63 ],
   alphaCSR[ 93 ][ 64 ],
   alphaCSR[ 93 ][ 65 ],
   alphaCSR[ 93 ][ 66 ],
   alphaCSR[ 93 ][ 67 ],
   alphaCSR[ 93 ][ 68 ],
   alphaCSR[ 93 ][ 69 ],
   alphaCSR[ 93 ][ 70 ],
   alphaCSR[ 93 ][ 71 ],
   alphaCSR[ 93 ][ 72 ],
   alphaCSR[ 93 ][ 73 ],
   alphaCSR[ 93 ][ 74 ],
   alphaCSR[ 93 ][ 75 ],
   alphaCSR[ 93 ][ 76 ],
   alphaCSR[ 93 ][ 77 ],
   alphaCSR[ 93 ][ 78 ],
   alphaCSR[ 93 ][ 79 ],
   alphaCSR[ 93 ][ 80 ],
   alphaCSR[ 93 ][ 81 ],
   alphaCSR[ 93 ][ 82 ],
   alphaCSR[ 93 ][ 83 ],
   alphaCSR[ 93 ][ 84 ],
   alphaCSR[ 93 ][ 85 ],
   alphaCSR[ 93 ][ 86 ],
   alphaCSR[ 93 ][ 87 ],
   alphaCSR[ 93 ][ 88 ],
   alphaCSR[ 93 ][ 89 ],
   alphaCSR[ 93 ][ 90 ],
   alphaCSR[ 93 ][ 91 ],
   alphaCSR[ 93 ][ 92 ],
   alphaCSR[ 93 ][ 93 ],
   alphaCSR[ 93 ][ 94 ],
   alphaCSR[ 93 ][ 95 ],
   alphaCSR[ 93 ][ 96 ],
   alphaCSR[ 93 ][ 97 ],
   alphaCSR[ 93 ][ 98 ],
   alphaCSR[ 93 ][ 99 ],
   alphaCSR[ 93 ][ 100 ],
   alphaCSR[ 93 ][ 101 ],
   alphaCSR[ 93 ][ 102 ],
   alphaCSR[ 93 ][ 103 ],
   alphaCSR[ 93 ][ 104 ],
   alphaCSR[ 93 ][ 105 ],
   alphaCSR[ 93 ][ 106 ],
   alphaCSR[ 93 ][ 107 ],
   alphaCSR[ 93 ][ 108 ],
   alphaCSR[ 93 ][ 109 ],
   alphaCSR[ 93 ][ 110 ],
   alphaCSR[ 93 ][ 111 ],
   alphaCSR[ 93 ][ 112 ],
   alphaCSR[ 93 ][ 113 ],
   alphaCSR[ 93 ][ 114 ],
   alphaCSR[ 93 ][ 115 ],
   alphaCSR[ 93 ][ 116 ],
   alphaCSR[ 93 ][ 117 ],
   alphaCSR[ 93 ][ 118 ],
   alphaCSR[ 93 ][ 119 ],
   alphaCSR[ 93 ][ 120 ],
   alphaCSR[ 93 ][ 121 ],
   alphaCSR[ 93 ][ 122 ],
   alphaCSR[ 93 ][ 123 ],
   alphaCSR[ 93 ][ 124 ],
   alphaCSR[ 93 ][ 125 ],
   alphaCSR[ 93 ][ 126 ],
   alphaCSR[ 93 ][ 127 ],
   alphaCSR[ 93 ][ 128 ],
   alphaCSR[ 93 ][ 129 ],
   alphaCSR[ 93 ][ 130 ],
   alphaCSR[ 93 ][ 131 ],
   alphaCSR[ 93 ][ 132 ],
   alphaCSR[ 93 ][ 133 ],
   alphaCSR[ 93 ][ 134 ],
   alphaCSR[ 93 ][ 135 ],
   alphaCSR[ 93 ][ 136 ],
   alphaCSR[ 93 ][ 137 ],
   alphaCSR[ 93 ][ 138 ],
   alphaCSR[ 93 ][ 139 ],
   alphaCSR[ 93 ][ 140 ],
   alphaCSR[ 93 ][ 141 ],
   alphaCSR[ 93 ][ 142 ],
   alphaCSR[ 93 ][ 143 ],
   alphaCSR[ 93 ][ 144 ],
   alphaCSR[ 93 ][ 145 ],
   alphaCSR[ 93 ][ 146 ],
   alphaCSR[ 93 ][ 147 ],
   alphaCSR[ 93 ][ 148 ],
   alphaCSR[ 93 ][ 149 ],
   alphaCSR[ 93 ][ 150 ],
   alphaCSR[ 93 ][ 151 ],
   alphaCSR[ 93 ][ 152 ],
   alphaCSR[ 93 ][ 153 ],
   alphaCSR[ 93 ][ 154 ],
   alphaCSR[ 93 ][ 155 ],
   alphaCSR[ 93 ][ 156 ],
   alphaCSR[ 93 ][ 157 ],
   alphaCSR[ 93 ][ 158 ],
   alphaCSR[ 93 ][ 159 ],
   alphaCSR[ 93 ][ 160 ],
   alphaCSR[ 93 ][ 161 ],
   alphaCSR[ 93 ][ 162 ],
   alphaCSR[ 93 ][ 163 ],
   alphaCSR[ 93 ][ 164 ],
   alphaCSR[ 93 ][ 165 ],
   alphaCSR[ 93 ][ 166 ],
   alphaCSR[ 93 ][ 167 ],
   alphaCSR[ 93 ][ 168 ],
   alphaCSR[ 93 ][ 169 ],
   alphaCSR[ 93 ][ 170 ],
   alphaCSR[ 93 ][ 171 ],
   alphaCSR[ 93 ][ 172 ],
   alphaCSR[ 93 ][ 173 ],
   alphaCSR[ 93 ][ 174 ],
   alphaCSR[ 93 ][ 175 ],
   alphaCSR[ 93 ][ 176 ],
   alphaCSR[ 93 ][ 177 ],
   alphaCSR[ 93 ][ 178 ],
   alphaCSR[ 93 ][ 179 ],
   alphaCSR[ 93 ][ 180 ],
   alphaCSR[ 93 ][ 181 ],
   alphaCSR[ 93 ][ 182 ],
   alphaCSR[ 93 ][ 183 ],
   alphaCSR[ 93 ][ 184 ],
   alphaCSR[ 93 ][ 185 ],
   alphaCSR[ 93 ][ 186 ],
   alphaCSR[ 93 ][ 187 ],
   alphaCSR[ 93 ][ 188 ],
   alphaCSR[ 93 ][ 189 ],
   alphaCSR[ 93 ][ 190 ],
   alphaCSR[ 93 ][ 191 ],
   alphaCSR[ 93 ][ 192 ],
   alphaCSR[ 93 ][ 193 ],
   alphaCSR[ 93 ][ 194 ],
   alphaCSR[ 93 ][ 195 ],
   alphaCSR[ 93 ][ 196 ],
   alphaCSR[ 93 ][ 197 ],
   alphaCSR[ 93 ][ 198 ],
   alphaCSR[ 93 ][ 199 ],
   alphaCSR[ 93 ][ 200 ],
   alphaCSR[ 93 ][ 201 ],
   alphaCSR[ 93 ][ 202 ],
   alphaCSR[ 93 ][ 203 ],
   alphaCSR[ 93 ][ 204 ],
   alphaCSR[ 93 ][ 205 ],
   alphaCSR[ 93 ][ 206 ],
   alphaCSR[ 93 ][ 207 ],
   alphaCSR[ 93 ][ 208 ],
   alphaCSR[ 93 ][ 209 ],
   alphaCSR[ 93 ][ 210 ],
   alphaCSR[ 93 ][ 211 ],
   alphaCSR[ 93 ][ 212 ],
   alphaCSR[ 93 ][ 213 ],
   alphaCSR[ 93 ][ 214 ],
   alphaCSR[ 93 ][ 215 ],
   alphaCSR[ 93 ][ 216 ],
   alphaCSR[ 93 ][ 217 ],
   alphaCSR[ 93 ][ 218 ],
   alphaCSR[ 93 ][ 219 ],
   alphaCSR[ 93 ][ 220 ],
   alphaCSR[ 93 ][ 221 ],
   alphaCSR[ 93 ][ 222 ],
   alphaCSR[ 93 ][ 223 ],
   alphaCSR[ 93 ][ 224 ],
   alphaCSR[ 93 ][ 225 ],
   alphaCSR[ 93 ][ 226 ],
   alphaCSR[ 93 ][ 227 ],
   alphaCSR[ 93 ][ 228 ],
   alphaCSR[ 93 ][ 229 ],
   alphaCSR[ 93 ][ 230 ],
   alphaCSR[ 93 ][ 231 ],
   alphaCSR[ 93 ][ 232 ],
   alphaCSR[ 93 ][ 233 ],
   alphaCSR[ 93 ][ 234 ],
   alphaCSR[ 93 ][ 235 ],
   alphaCSR[ 93 ][ 236 ],
   alphaCSR[ 93 ][ 237 ],
   alphaCSR[ 93 ][ 238 ],
   alphaCSR[ 93 ][ 239 ],
   alphaCSR[ 93 ][ 240 ],
   alphaCSR[ 93 ][ 241 ],
   alphaCSR[ 93 ][ 242 ],
   alphaCSR[ 93 ][ 243 ],
   alphaCSR[ 93 ][ 244 ],
   alphaCSR[ 93 ][ 245 ],
   alphaCSR[ 93 ][ 246 ],
   alphaCSR[ 93 ][ 247 ],
   alphaCSR[ 93 ][ 248 ],
   alphaCSR[ 93 ][ 249 ],
   alphaCSR[ 93 ][ 250 ],
   alphaCSR[ 93 ][ 251 ],
   alphaCSR[ 93 ][ 252 ],
   alphaCSR[ 93 ][ 253 ],
   alphaCSR[ 93 ][ 254 ],
   alphaCSR[ 93 ][ 255 ],
   alphaCSR[ 93 ][ 256 ],
   alphaCSR[ 93 ][ 257 ],
   alphaCSR[ 93 ][ 258 ],
   alphaCSR[ 93 ][ 259 ],
   alphaCSR[ 93 ][ 260 ],
   alphaCSR[ 93 ][ 261 ],
   alphaCSR[ 93 ][ 262 ],
   alphaCSR[ 93 ][ 263 ],
   alphaCSR[ 93 ][ 264 ],
   alphaCSR[ 93 ][ 265 ],
   alphaCSR[ 93 ][ 266 ],
   alphaCSR[ 93 ][ 267 ],
   alphaCSR[ 93 ][ 268 ],
   alphaCSR[ 93 ][ 269 ],
   alphaCSR[ 93 ][ 270 ],
   alphaCSR[ 93 ][ 271 ],
   alphaCSR[ 93 ][ 272 ],
   alphaCSR[ 93 ][ 273 ],
   alphaCSR[ 93 ][ 274 ],
   alphaCSR[ 93 ][ 275 ],
   alphaCSR[ 93 ][ 276 ],
   alphaCSR[ 93 ][ 277 ],
   alphaCSR[ 93 ][ 278 ],
   alphaCSR[ 93 ][ 279 ],
   alphaCSR[ 93 ][ 280 ],
   alphaCSR[ 93 ][ 281 ],
   alphaCSR[ 93 ][ 282 ],
   alphaCSR[ 93 ][ 283 ],
   alphaCSR[ 93 ][ 284 ],
   alphaCSR[ 93 ][ 285 ],
   alphaCSR[ 93 ][ 286 ],
   alphaCSR[ 93 ][ 287 ],
   alphaCSR[ 93 ][ 288 ],
   alphaCSR[ 93 ][ 289 ],
   alphaCSR[ 93 ][ 290 ],
   alphaCSR[ 93 ][ 291 ],
   alphaCSR[ 93 ][ 292 ],
   alphaCSR[ 93 ][ 293 ],
   alphaCSR[ 93 ][ 294 ],
   alphaCSR[ 93 ][ 295 ],
   alphaCSR[ 93 ][ 296 ],
   alphaCSR[ 93 ][ 297 ],
   alphaCSR[ 93 ][ 298 ],
   alphaCSR[ 93 ][ 299 ],
   alphaCSR[ 93 ][ 300 ],
   alphaCSR[ 93 ][ 301 ],
   alphaCSR[ 93 ][ 302 ],
   alphaCSR[ 93 ][ 303 ],
   alphaCSR[ 93 ][ 304 ],
   alphaCSR[ 93 ][ 305 ],
   alphaCSR[ 93 ][ 306 ],
   alphaCSR[ 93 ][ 307 ],
   alphaCSR[ 93 ][ 308 ],
   alphaCSR[ 93 ][ 309 ],
   alphaCSR[ 93 ][ 310 ],
   alphaCSR[ 93 ][ 311 ],
   alphaCSR[ 93 ][ 312 ],
   alphaCSR[ 93 ][ 313 ],
   alphaCSR[ 93 ][ 314 ],
   alphaCSR[ 93 ][ 315 ],
   alphaCSR[ 93 ][ 316 ],
   alphaCSR[ 93 ][ 317 ],
   alphaCSR[ 93 ][ 318 ],
   alphaCSR[ 93 ][ 319 ],
   alphaCSR[ 93 ][ 320 ],
   alphaCSR[ 93 ][ 321 ],
   alphaCSR[ 93 ][ 322 ],
   alphaCSR[ 93 ][ 323 ],
   alphaCSR[ 93 ][ 324 ],
   alphaCSR[ 93 ][ 325 ],
   alphaCSR[ 93 ][ 326 ],
   alphaCSR[ 93 ][ 327 ],
   alphaCSR[ 93 ][ 328 ],
   alphaCSR[ 93 ][ 329 ],
   alphaCSR[ 93 ][ 330 ],
   alphaCSR[ 93 ][ 331 ],
   alphaCSR[ 93 ][ 332 ],
   alphaCSR[ 93 ][ 333 ],
   alphaCSR[ 93 ][ 334 ],
   alphaCSR[ 93 ][ 335 ],
   alphaCSR[ 93 ][ 336 ],
   alphaCSR[ 93 ][ 337 ],
   alphaCSR[ 93 ][ 338 ],
   alphaCSR[ 93 ][ 339 ],
   alphaCSR[ 93 ][ 340 ],
   alphaCSR[ 93 ][ 341 ],
   alphaCSR[ 93 ][ 342 ],
   alphaCSR[ 93 ][ 343 ],
   alphaCSR[ 93 ][ 344 ],
   alphaCSR[ 93 ][ 345 ],
   alphaCSR[ 93 ][ 346 ],
   alphaCSR[ 93 ][ 347 ],
   alphaCSR[ 93 ][ 348 ],
   alphaCSR[ 93 ][ 349 ],
   alphaCSR[ 93 ][ 350 ],
   alphaCSR[ 93 ][ 351 ],
   alphaCSR[ 93 ][ 352 ],
   alphaCSR[ 93 ][ 353 ],
   alphaCSR[ 93 ][ 354 ],
   alphaCSR[ 93 ][ 355 ],
   alphaCSR[ 93 ][ 356 ],
   alphaCSR[ 93 ][ 357 ],
   alphaCSR[ 93 ][ 358 ],
   alphaCSR[ 93 ][ 359 ],
   alphaCSR[ 93 ][ 360 ],
   alphaCSR[ 93 ][ 361 ],
   alphaCSR[ 93 ][ 362 ],
   alphaCSR[ 93 ][ 363 ],
   alphaCSR[ 93 ][ 364 ],
   alphaCSR[ 93 ][ 365 ],
   alphaCSR[ 93 ][ 366 ],
   alphaCSR[ 93 ][ 367 ],
   alphaCSR[ 93 ][ 368 ],
   alphaCSR[ 93 ][ 369 ],
   alphaCSR[ 93 ][ 370 ],
   alphaCSR[ 93 ][ 371 ],
   alphaCSR[ 93 ][ 372 ],
   alphaCSR[ 93 ][ 373 ],
   alphaCSR[ 93 ][ 374 ],
   alphaCSR[ 93 ][ 375 ],
   alphaCSR[ 93 ][ 376 ],
   alphaCSR[ 93 ][ 377 ],
   alphaCSR[ 93 ][ 378 ],
   alphaCSR[ 93 ][ 379 ],
   alphaCSR[ 93 ][ 380 ],
   alphaCSR[ 93 ][ 381 ],
   alphaCSR[ 93 ][ 382 ],
   alphaCSR[ 93 ][ 383 ],
   alphaCSR[ 94 ][ 0 ],
   alphaCSR[ 94 ][ 1 ],
   alphaCSR[ 94 ][ 2 ],
   alphaCSR[ 94 ][ 3 ],
   alphaCSR[ 94 ][ 4 ],
   alphaCSR[ 94 ][ 5 ],
   alphaCSR[ 94 ][ 6 ],
   alphaCSR[ 94 ][ 7 ],
   alphaCSR[ 94 ][ 8 ],
   alphaCSR[ 94 ][ 9 ],
   alphaCSR[ 94 ][ 10 ],
   alphaCSR[ 94 ][ 11 ],
   alphaCSR[ 94 ][ 12 ],
   alphaCSR[ 94 ][ 13 ],
   alphaCSR[ 94 ][ 14 ],
   alphaCSR[ 94 ][ 15 ],
   alphaCSR[ 94 ][ 16 ],
   alphaCSR[ 94 ][ 17 ],
   alphaCSR[ 94 ][ 18 ],
   alphaCSR[ 94 ][ 19 ],
   alphaCSR[ 94 ][ 20 ],
   alphaCSR[ 94 ][ 21 ],
   alphaCSR[ 94 ][ 22 ],
   alphaCSR[ 94 ][ 23 ],
   alphaCSR[ 94 ][ 24 ],
   alphaCSR[ 94 ][ 25 ],
   alphaCSR[ 94 ][ 26 ],
   alphaCSR[ 94 ][ 27 ],
   alphaCSR[ 94 ][ 28 ],
   alphaCSR[ 94 ][ 29 ],
   alphaCSR[ 94 ][ 30 ],
   alphaCSR[ 94 ][ 31 ],
   alphaCSR[ 94 ][ 32 ],
   alphaCSR[ 94 ][ 33 ],
   alphaCSR[ 94 ][ 34 ],
   alphaCSR[ 94 ][ 35 ],
   alphaCSR[ 94 ][ 36 ],
   alphaCSR[ 94 ][ 37 ],
   alphaCSR[ 94 ][ 38 ],
   alphaCSR[ 94 ][ 39 ],
   alphaCSR[ 94 ][ 40 ],
   alphaCSR[ 94 ][ 41 ],
   alphaCSR[ 94 ][ 42 ],
   alphaCSR[ 94 ][ 43 ],
   alphaCSR[ 94 ][ 44 ],
   alphaCSR[ 94 ][ 45 ],
   alphaCSR[ 94 ][ 46 ],
   alphaCSR[ 94 ][ 47 ],
   alphaCSR[ 94 ][ 48 ],
   alphaCSR[ 94 ][ 49 ],
   alphaCSR[ 94 ][ 50 ],
   alphaCSR[ 94 ][ 51 ],
   alphaCSR[ 94 ][ 52 ],
   alphaCSR[ 94 ][ 53 ],
   alphaCSR[ 94 ][ 54 ],
   alphaCSR[ 94 ][ 55 ],
   alphaCSR[ 94 ][ 56 ],
   alphaCSR[ 94 ][ 57 ],
   alphaCSR[ 94 ][ 58 ],
   alphaCSR[ 94 ][ 59 ],
   alphaCSR[ 94 ][ 60 ],
   alphaCSR[ 94 ][ 61 ],
   alphaCSR[ 94 ][ 62 ],
   alphaCSR[ 94 ][ 63 ],
   alphaCSR[ 94 ][ 64 ],
   alphaCSR[ 94 ][ 65 ],
   alphaCSR[ 94 ][ 66 ],
   alphaCSR[ 94 ][ 67 ],
   alphaCSR[ 94 ][ 68 ],
   alphaCSR[ 94 ][ 69 ],
   alphaCSR[ 94 ][ 70 ],
   alphaCSR[ 94 ][ 71 ],
   alphaCSR[ 94 ][ 72 ],
   alphaCSR[ 94 ][ 73 ],
   alphaCSR[ 94 ][ 74 ],
   alphaCSR[ 94 ][ 75 ],
   alphaCSR[ 94 ][ 76 ],
   alphaCSR[ 94 ][ 77 ],
   alphaCSR[ 94 ][ 78 ],
   alphaCSR[ 94 ][ 79 ],
   alphaCSR[ 94 ][ 80 ],
   alphaCSR[ 94 ][ 81 ],
   alphaCSR[ 94 ][ 82 ],
   alphaCSR[ 94 ][ 83 ],
   alphaCSR[ 94 ][ 84 ],
   alphaCSR[ 94 ][ 85 ],
   alphaCSR[ 94 ][ 86 ],
   alphaCSR[ 94 ][ 87 ],
   alphaCSR[ 94 ][ 88 ],
   alphaCSR[ 94 ][ 89 ],
   alphaCSR[ 94 ][ 90 ],
   alphaCSR[ 94 ][ 91 ],
   alphaCSR[ 94 ][ 92 ],
   alphaCSR[ 94 ][ 93 ],
   alphaCSR[ 94 ][ 94 ],
   alphaCSR[ 94 ][ 95 ],
   alphaCSR[ 94 ][ 96 ],
   alphaCSR[ 94 ][ 97 ],
   alphaCSR[ 94 ][ 98 ],
   alphaCSR[ 94 ][ 99 ],
   alphaCSR[ 94 ][ 100 ],
   alphaCSR[ 94 ][ 101 ],
   alphaCSR[ 94 ][ 102 ],
   alphaCSR[ 94 ][ 103 ],
   alphaCSR[ 94 ][ 104 ],
   alphaCSR[ 94 ][ 105 ],
   alphaCSR[ 94 ][ 106 ],
   alphaCSR[ 94 ][ 107 ],
   alphaCSR[ 94 ][ 108 ],
   alphaCSR[ 94 ][ 109 ],
   alphaCSR[ 94 ][ 110 ],
   alphaCSR[ 94 ][ 111 ],
   alphaCSR[ 94 ][ 112 ],
   alphaCSR[ 94 ][ 113 ],
   alphaCSR[ 94 ][ 114 ],
   alphaCSR[ 94 ][ 115 ],
   alphaCSR[ 94 ][ 116 ],
   alphaCSR[ 94 ][ 117 ],
   alphaCSR[ 94 ][ 118 ],
   alphaCSR[ 94 ][ 119 ],
   alphaCSR[ 94 ][ 120 ],
   alphaCSR[ 94 ][ 121 ],
   alphaCSR[ 94 ][ 122 ],
   alphaCSR[ 94 ][ 123 ],
   alphaCSR[ 94 ][ 124 ],
   alphaCSR[ 94 ][ 125 ],
   alphaCSR[ 94 ][ 126 ],
   alphaCSR[ 94 ][ 127 ],
   alphaCSR[ 94 ][ 128 ],
   alphaCSR[ 94 ][ 129 ],
   alphaCSR[ 94 ][ 130 ],
   alphaCSR[ 94 ][ 131 ],
   alphaCSR[ 94 ][ 132 ],
   alphaCSR[ 94 ][ 133 ],
   alphaCSR[ 94 ][ 134 ],
   alphaCSR[ 94 ][ 135 ],
   alphaCSR[ 94 ][ 136 ],
   alphaCSR[ 94 ][ 137 ],
   alphaCSR[ 94 ][ 138 ],
   alphaCSR[ 94 ][ 139 ],
   alphaCSR[ 94 ][ 140 ],
   alphaCSR[ 94 ][ 141 ],
   alphaCSR[ 94 ][ 142 ],
   alphaCSR[ 94 ][ 143 ],
   alphaCSR[ 94 ][ 144 ],
   alphaCSR[ 94 ][ 145 ],
   alphaCSR[ 94 ][ 146 ],
   alphaCSR[ 94 ][ 147 ],
   alphaCSR[ 94 ][ 148 ],
   alphaCSR[ 94 ][ 149 ],
   alphaCSR[ 94 ][ 150 ],
   alphaCSR[ 94 ][ 151 ],
   alphaCSR[ 94 ][ 152 ],
   alphaCSR[ 94 ][ 153 ],
   alphaCSR[ 94 ][ 154 ],
   alphaCSR[ 94 ][ 155 ],
   alphaCSR[ 94 ][ 156 ],
   alphaCSR[ 94 ][ 157 ],
   alphaCSR[ 94 ][ 158 ],
   alphaCSR[ 94 ][ 159 ],
   alphaCSR[ 94 ][ 160 ],
   alphaCSR[ 94 ][ 161 ],
   alphaCSR[ 94 ][ 162 ],
   alphaCSR[ 94 ][ 163 ],
   alphaCSR[ 94 ][ 164 ],
   alphaCSR[ 94 ][ 165 ],
   alphaCSR[ 94 ][ 166 ],
   alphaCSR[ 94 ][ 167 ],
   alphaCSR[ 94 ][ 168 ],
   alphaCSR[ 94 ][ 169 ],
   alphaCSR[ 94 ][ 170 ],
   alphaCSR[ 94 ][ 171 ],
   alphaCSR[ 94 ][ 172 ],
   alphaCSR[ 94 ][ 173 ],
   alphaCSR[ 94 ][ 174 ],
   alphaCSR[ 94 ][ 175 ],
   alphaCSR[ 94 ][ 176 ],
   alphaCSR[ 94 ][ 177 ],
   alphaCSR[ 94 ][ 178 ],
   alphaCSR[ 94 ][ 179 ],
   alphaCSR[ 94 ][ 180 ],
   alphaCSR[ 94 ][ 181 ],
   alphaCSR[ 94 ][ 182 ],
   alphaCSR[ 94 ][ 183 ],
   alphaCSR[ 94 ][ 184 ],
   alphaCSR[ 94 ][ 185 ],
   alphaCSR[ 94 ][ 186 ],
   alphaCSR[ 94 ][ 187 ],
   alphaCSR[ 94 ][ 188 ],
   alphaCSR[ 94 ][ 189 ],
   alphaCSR[ 94 ][ 190 ],
   alphaCSR[ 94 ][ 191 ],
   alphaCSR[ 94 ][ 192 ],
   alphaCSR[ 94 ][ 193 ],
   alphaCSR[ 94 ][ 194 ],
   alphaCSR[ 94 ][ 195 ],
   alphaCSR[ 94 ][ 196 ],
   alphaCSR[ 94 ][ 197 ],
   alphaCSR[ 94 ][ 198 ],
   alphaCSR[ 94 ][ 199 ],
   alphaCSR[ 94 ][ 200 ],
   alphaCSR[ 94 ][ 201 ],
   alphaCSR[ 94 ][ 202 ],
   alphaCSR[ 94 ][ 203 ],
   alphaCSR[ 94 ][ 204 ],
   alphaCSR[ 94 ][ 205 ],
   alphaCSR[ 94 ][ 206 ],
   alphaCSR[ 94 ][ 207 ],
   alphaCSR[ 94 ][ 208 ],
   alphaCSR[ 94 ][ 209 ],
   alphaCSR[ 94 ][ 210 ],
   alphaCSR[ 94 ][ 211 ],
   alphaCSR[ 94 ][ 212 ],
   alphaCSR[ 94 ][ 213 ],
   alphaCSR[ 94 ][ 214 ],
   alphaCSR[ 94 ][ 215 ],
   alphaCSR[ 94 ][ 216 ],
   alphaCSR[ 94 ][ 217 ],
   alphaCSR[ 94 ][ 218 ],
   alphaCSR[ 94 ][ 219 ],
   alphaCSR[ 94 ][ 220 ],
   alphaCSR[ 94 ][ 221 ],
   alphaCSR[ 94 ][ 222 ],
   alphaCSR[ 94 ][ 223 ],
   alphaCSR[ 94 ][ 224 ],
   alphaCSR[ 94 ][ 225 ],
   alphaCSR[ 94 ][ 226 ],
   alphaCSR[ 94 ][ 227 ],
   alphaCSR[ 94 ][ 228 ],
   alphaCSR[ 94 ][ 229 ],
   alphaCSR[ 94 ][ 230 ],
   alphaCSR[ 94 ][ 231 ],
   alphaCSR[ 94 ][ 232 ],
   alphaCSR[ 94 ][ 233 ],
   alphaCSR[ 94 ][ 234 ],
   alphaCSR[ 94 ][ 235 ],
   alphaCSR[ 94 ][ 236 ],
   alphaCSR[ 94 ][ 237 ],
   alphaCSR[ 94 ][ 238 ],
   alphaCSR[ 94 ][ 239 ],
   alphaCSR[ 94 ][ 240 ],
   alphaCSR[ 94 ][ 241 ],
   alphaCSR[ 94 ][ 242 ],
   alphaCSR[ 94 ][ 243 ],
   alphaCSR[ 94 ][ 244 ],
   alphaCSR[ 94 ][ 245 ],
   alphaCSR[ 94 ][ 246 ],
   alphaCSR[ 94 ][ 247 ],
   alphaCSR[ 94 ][ 248 ],
   alphaCSR[ 94 ][ 249 ],
   alphaCSR[ 94 ][ 250 ],
   alphaCSR[ 94 ][ 251 ],
   alphaCSR[ 94 ][ 252 ],
   alphaCSR[ 94 ][ 253 ],
   alphaCSR[ 94 ][ 254 ],
   alphaCSR[ 94 ][ 255 ],
   alphaCSR[ 94 ][ 256 ],
   alphaCSR[ 94 ][ 257 ],
   alphaCSR[ 94 ][ 258 ],
   alphaCSR[ 94 ][ 259 ],
   alphaCSR[ 94 ][ 260 ],
   alphaCSR[ 94 ][ 261 ],
   alphaCSR[ 94 ][ 262 ],
   alphaCSR[ 94 ][ 263 ],
   alphaCSR[ 94 ][ 264 ],
   alphaCSR[ 94 ][ 265 ],
   alphaCSR[ 94 ][ 266 ],
   alphaCSR[ 94 ][ 267 ],
   alphaCSR[ 94 ][ 268 ],
   alphaCSR[ 94 ][ 269 ],
   alphaCSR[ 94 ][ 270 ],
   alphaCSR[ 94 ][ 271 ],
   alphaCSR[ 94 ][ 272 ],
   alphaCSR[ 94 ][ 273 ],
   alphaCSR[ 94 ][ 274 ],
   alphaCSR[ 94 ][ 275 ],
   alphaCSR[ 94 ][ 276 ],
   alphaCSR[ 94 ][ 277 ],
   alphaCSR[ 94 ][ 278 ],
   alphaCSR[ 94 ][ 279 ],
   alphaCSR[ 94 ][ 280 ],
   alphaCSR[ 94 ][ 281 ],
   alphaCSR[ 94 ][ 282 ],
   alphaCSR[ 94 ][ 283 ],
   alphaCSR[ 94 ][ 284 ],
   alphaCSR[ 94 ][ 285 ],
   alphaCSR[ 94 ][ 286 ],
   alphaCSR[ 94 ][ 287 ],
   alphaCSR[ 94 ][ 288 ],
   alphaCSR[ 94 ][ 289 ],
   alphaCSR[ 94 ][ 290 ],
   alphaCSR[ 94 ][ 291 ],
   alphaCSR[ 94 ][ 292 ],
   alphaCSR[ 94 ][ 293 ],
   alphaCSR[ 94 ][ 294 ],
   alphaCSR[ 94 ][ 295 ],
   alphaCSR[ 94 ][ 296 ],
   alphaCSR[ 94 ][ 297 ],
   alphaCSR[ 94 ][ 298 ],
   alphaCSR[ 94 ][ 299 ],
   alphaCSR[ 94 ][ 300 ],
   alphaCSR[ 94 ][ 301 ],
   alphaCSR[ 94 ][ 302 ],
   alphaCSR[ 94 ][ 303 ],
   alphaCSR[ 94 ][ 304 ],
   alphaCSR[ 94 ][ 305 ],
   alphaCSR[ 94 ][ 306 ],
   alphaCSR[ 94 ][ 307 ],
   alphaCSR[ 94 ][ 308 ],
   alphaCSR[ 94 ][ 309 ],
   alphaCSR[ 94 ][ 310 ],
   alphaCSR[ 94 ][ 311 ],
   alphaCSR[ 94 ][ 312 ],
   alphaCSR[ 94 ][ 313 ],
   alphaCSR[ 94 ][ 314 ],
   alphaCSR[ 94 ][ 315 ],
   alphaCSR[ 94 ][ 316 ],
   alphaCSR[ 94 ][ 317 ],
   alphaCSR[ 94 ][ 318 ],
   alphaCSR[ 94 ][ 319 ],
   alphaCSR[ 94 ][ 320 ],
   alphaCSR[ 94 ][ 321 ],
   alphaCSR[ 94 ][ 322 ],
   alphaCSR[ 94 ][ 323 ],
   alphaCSR[ 94 ][ 324 ],
   alphaCSR[ 94 ][ 325 ],
   alphaCSR[ 94 ][ 326 ],
   alphaCSR[ 94 ][ 327 ],
   alphaCSR[ 94 ][ 328 ],
   alphaCSR[ 94 ][ 329 ],
   alphaCSR[ 94 ][ 330 ],
   alphaCSR[ 94 ][ 331 ],
   alphaCSR[ 94 ][ 332 ],
   alphaCSR[ 94 ][ 333 ],
   alphaCSR[ 94 ][ 334 ],
   alphaCSR[ 94 ][ 335 ],
   alphaCSR[ 94 ][ 336 ],
   alphaCSR[ 94 ][ 337 ],
   alphaCSR[ 94 ][ 338 ],
   alphaCSR[ 94 ][ 339 ],
   alphaCSR[ 94 ][ 340 ],
   alphaCSR[ 94 ][ 341 ],
   alphaCSR[ 94 ][ 342 ],
   alphaCSR[ 94 ][ 343 ],
   alphaCSR[ 94 ][ 344 ],
   alphaCSR[ 94 ][ 345 ],
   alphaCSR[ 94 ][ 346 ],
   alphaCSR[ 94 ][ 347 ],
   alphaCSR[ 94 ][ 348 ],
   alphaCSR[ 94 ][ 349 ],
   alphaCSR[ 94 ][ 350 ],
   alphaCSR[ 94 ][ 351 ],
   alphaCSR[ 94 ][ 352 ],
   alphaCSR[ 94 ][ 353 ],
   alphaCSR[ 94 ][ 354 ],
   alphaCSR[ 94 ][ 355 ],
   alphaCSR[ 94 ][ 356 ],
   alphaCSR[ 94 ][ 357 ],
   alphaCSR[ 94 ][ 358 ],
   alphaCSR[ 94 ][ 359 ],
   alphaCSR[ 94 ][ 360 ],
   alphaCSR[ 94 ][ 361 ],
   alphaCSR[ 94 ][ 362 ],
   alphaCSR[ 94 ][ 363 ],
   alphaCSR[ 94 ][ 364 ],
   alphaCSR[ 94 ][ 365 ],
   alphaCSR[ 94 ][ 366 ],
   alphaCSR[ 94 ][ 367 ],
   alphaCSR[ 94 ][ 368 ],
   alphaCSR[ 94 ][ 369 ],
   alphaCSR[ 94 ][ 370 ],
   alphaCSR[ 94 ][ 371 ],
   alphaCSR[ 94 ][ 372 ],
   alphaCSR[ 94 ][ 373 ],
   alphaCSR[ 94 ][ 374 ],
   alphaCSR[ 94 ][ 375 ],
   alphaCSR[ 94 ][ 376 ],
   alphaCSR[ 94 ][ 377 ],
   alphaCSR[ 94 ][ 378 ],
   alphaCSR[ 94 ][ 379 ],
   alphaCSR[ 94 ][ 380 ],
   alphaCSR[ 94 ][ 381 ],
   alphaCSR[ 94 ][ 382 ],
   alphaCSR[ 94 ][ 383 ],
   alphaCSR[ 95 ][ 0 ],
   alphaCSR[ 95 ][ 1 ],
   alphaCSR[ 95 ][ 2 ],
   alphaCSR[ 95 ][ 3 ],
   alphaCSR[ 95 ][ 4 ],
   alphaCSR[ 95 ][ 5 ],
   alphaCSR[ 95 ][ 6 ],
   alphaCSR[ 95 ][ 7 ],
   alphaCSR[ 95 ][ 8 ],
   alphaCSR[ 95 ][ 9 ],
   alphaCSR[ 95 ][ 10 ],
   alphaCSR[ 95 ][ 11 ],
   alphaCSR[ 95 ][ 12 ],
   alphaCSR[ 95 ][ 13 ],
   alphaCSR[ 95 ][ 14 ],
   alphaCSR[ 95 ][ 15 ],
   alphaCSR[ 95 ][ 16 ],
   alphaCSR[ 95 ][ 17 ],
   alphaCSR[ 95 ][ 18 ],
   alphaCSR[ 95 ][ 19 ],
   alphaCSR[ 95 ][ 20 ],
   alphaCSR[ 95 ][ 21 ],
   alphaCSR[ 95 ][ 22 ],
   alphaCSR[ 95 ][ 23 ],
   alphaCSR[ 95 ][ 24 ],
   alphaCSR[ 95 ][ 25 ],
   alphaCSR[ 95 ][ 26 ],
   alphaCSR[ 95 ][ 27 ],
   alphaCSR[ 95 ][ 28 ],
   alphaCSR[ 95 ][ 29 ],
   alphaCSR[ 95 ][ 30 ],
   alphaCSR[ 95 ][ 31 ],
   alphaCSR[ 95 ][ 32 ],
   alphaCSR[ 95 ][ 33 ],
   alphaCSR[ 95 ][ 34 ],
   alphaCSR[ 95 ][ 35 ],
   alphaCSR[ 95 ][ 36 ],
   alphaCSR[ 95 ][ 37 ],
   alphaCSR[ 95 ][ 38 ],
   alphaCSR[ 95 ][ 39 ],
   alphaCSR[ 95 ][ 40 ],
   alphaCSR[ 95 ][ 41 ],
   alphaCSR[ 95 ][ 42 ],
   alphaCSR[ 95 ][ 43 ],
   alphaCSR[ 95 ][ 44 ],
   alphaCSR[ 95 ][ 45 ],
   alphaCSR[ 95 ][ 46 ],
   alphaCSR[ 95 ][ 47 ],
   alphaCSR[ 95 ][ 48 ],
   alphaCSR[ 95 ][ 49 ],
   alphaCSR[ 95 ][ 50 ],
   alphaCSR[ 95 ][ 51 ],
   alphaCSR[ 95 ][ 52 ],
   alphaCSR[ 95 ][ 53 ],
   alphaCSR[ 95 ][ 54 ],
   alphaCSR[ 95 ][ 55 ],
   alphaCSR[ 95 ][ 56 ],
   alphaCSR[ 95 ][ 57 ],
   alphaCSR[ 95 ][ 58 ],
   alphaCSR[ 95 ][ 59 ],
   alphaCSR[ 95 ][ 60 ],
   alphaCSR[ 95 ][ 61 ],
   alphaCSR[ 95 ][ 62 ],
   alphaCSR[ 95 ][ 63 ],
   alphaCSR[ 95 ][ 64 ],
   alphaCSR[ 95 ][ 65 ],
   alphaCSR[ 95 ][ 66 ],
   alphaCSR[ 95 ][ 67 ],
   alphaCSR[ 95 ][ 68 ],
   alphaCSR[ 95 ][ 69 ],
   alphaCSR[ 95 ][ 70 ],
   alphaCSR[ 95 ][ 71 ],
   alphaCSR[ 95 ][ 72 ],
   alphaCSR[ 95 ][ 73 ],
   alphaCSR[ 95 ][ 74 ],
   alphaCSR[ 95 ][ 75 ],
   alphaCSR[ 95 ][ 76 ],
   alphaCSR[ 95 ][ 77 ],
   alphaCSR[ 95 ][ 78 ],
   alphaCSR[ 95 ][ 79 ],
   alphaCSR[ 95 ][ 80 ],
   alphaCSR[ 95 ][ 81 ],
   alphaCSR[ 95 ][ 82 ],
   alphaCSR[ 95 ][ 83 ],
   alphaCSR[ 95 ][ 84 ],
   alphaCSR[ 95 ][ 85 ],
   alphaCSR[ 95 ][ 86 ],
   alphaCSR[ 95 ][ 87 ],
   alphaCSR[ 95 ][ 88 ],
   alphaCSR[ 95 ][ 89 ],
   alphaCSR[ 95 ][ 90 ],
   alphaCSR[ 95 ][ 91 ],
   alphaCSR[ 95 ][ 92 ],
   alphaCSR[ 95 ][ 93 ],
   alphaCSR[ 95 ][ 94 ],
   alphaCSR[ 95 ][ 95 ],
   alphaCSR[ 95 ][ 96 ],
   alphaCSR[ 95 ][ 97 ],
   alphaCSR[ 95 ][ 98 ],
   alphaCSR[ 95 ][ 99 ],
   alphaCSR[ 95 ][ 100 ],
   alphaCSR[ 95 ][ 101 ],
   alphaCSR[ 95 ][ 102 ],
   alphaCSR[ 95 ][ 103 ],
   alphaCSR[ 95 ][ 104 ],
   alphaCSR[ 95 ][ 105 ],
   alphaCSR[ 95 ][ 106 ],
   alphaCSR[ 95 ][ 107 ],
   alphaCSR[ 95 ][ 108 ],
   alphaCSR[ 95 ][ 109 ],
   alphaCSR[ 95 ][ 110 ],
   alphaCSR[ 95 ][ 111 ],
   alphaCSR[ 95 ][ 112 ],
   alphaCSR[ 95 ][ 113 ],
   alphaCSR[ 95 ][ 114 ],
   alphaCSR[ 95 ][ 115 ],
   alphaCSR[ 95 ][ 116 ],
   alphaCSR[ 95 ][ 117 ],
   alphaCSR[ 95 ][ 118 ],
   alphaCSR[ 95 ][ 119 ],
   alphaCSR[ 95 ][ 120 ],
   alphaCSR[ 95 ][ 121 ],
   alphaCSR[ 95 ][ 122 ],
   alphaCSR[ 95 ][ 123 ],
   alphaCSR[ 95 ][ 124 ],
   alphaCSR[ 95 ][ 125 ],
   alphaCSR[ 95 ][ 126 ],
   alphaCSR[ 95 ][ 127 ],
   alphaCSR[ 95 ][ 128 ],
   alphaCSR[ 95 ][ 129 ],
   alphaCSR[ 95 ][ 130 ],
   alphaCSR[ 95 ][ 131 ],
   alphaCSR[ 95 ][ 132 ],
   alphaCSR[ 95 ][ 133 ],
   alphaCSR[ 95 ][ 134 ],
   alphaCSR[ 95 ][ 135 ],
   alphaCSR[ 95 ][ 136 ],
   alphaCSR[ 95 ][ 137 ],
   alphaCSR[ 95 ][ 138 ],
   alphaCSR[ 95 ][ 139 ],
   alphaCSR[ 95 ][ 140 ],
   alphaCSR[ 95 ][ 141 ],
   alphaCSR[ 95 ][ 142 ],
   alphaCSR[ 95 ][ 143 ],
   alphaCSR[ 95 ][ 144 ],
   alphaCSR[ 95 ][ 145 ],
   alphaCSR[ 95 ][ 146 ],
   alphaCSR[ 95 ][ 147 ],
   alphaCSR[ 95 ][ 148 ],
   alphaCSR[ 95 ][ 149 ],
   alphaCSR[ 95 ][ 150 ],
   alphaCSR[ 95 ][ 151 ],
   alphaCSR[ 95 ][ 152 ],
   alphaCSR[ 95 ][ 153 ],
   alphaCSR[ 95 ][ 154 ],
   alphaCSR[ 95 ][ 155 ],
   alphaCSR[ 95 ][ 156 ],
   alphaCSR[ 95 ][ 157 ],
   alphaCSR[ 95 ][ 158 ],
   alphaCSR[ 95 ][ 159 ],
   alphaCSR[ 95 ][ 160 ],
   alphaCSR[ 95 ][ 161 ],
   alphaCSR[ 95 ][ 162 ],
   alphaCSR[ 95 ][ 163 ],
   alphaCSR[ 95 ][ 164 ],
   alphaCSR[ 95 ][ 165 ],
   alphaCSR[ 95 ][ 166 ],
   alphaCSR[ 95 ][ 167 ],
   alphaCSR[ 95 ][ 168 ],
   alphaCSR[ 95 ][ 169 ],
   alphaCSR[ 95 ][ 170 ],
   alphaCSR[ 95 ][ 171 ],
   alphaCSR[ 95 ][ 172 ],
   alphaCSR[ 95 ][ 173 ],
   alphaCSR[ 95 ][ 174 ],
   alphaCSR[ 95 ][ 175 ],
   alphaCSR[ 95 ][ 176 ],
   alphaCSR[ 95 ][ 177 ],
   alphaCSR[ 95 ][ 178 ],
   alphaCSR[ 95 ][ 179 ],
   alphaCSR[ 95 ][ 180 ],
   alphaCSR[ 95 ][ 181 ],
   alphaCSR[ 95 ][ 182 ],
   alphaCSR[ 95 ][ 183 ],
   alphaCSR[ 95 ][ 184 ],
   alphaCSR[ 95 ][ 185 ],
   alphaCSR[ 95 ][ 186 ],
   alphaCSR[ 95 ][ 187 ],
   alphaCSR[ 95 ][ 188 ],
   alphaCSR[ 95 ][ 189 ],
   alphaCSR[ 95 ][ 190 ],
   alphaCSR[ 95 ][ 191 ],
   alphaCSR[ 95 ][ 192 ],
   alphaCSR[ 95 ][ 193 ],
   alphaCSR[ 95 ][ 194 ],
   alphaCSR[ 95 ][ 195 ],
   alphaCSR[ 95 ][ 196 ],
   alphaCSR[ 95 ][ 197 ],
   alphaCSR[ 95 ][ 198 ],
   alphaCSR[ 95 ][ 199 ],
   alphaCSR[ 95 ][ 200 ],
   alphaCSR[ 95 ][ 201 ],
   alphaCSR[ 95 ][ 202 ],
   alphaCSR[ 95 ][ 203 ],
   alphaCSR[ 95 ][ 204 ],
   alphaCSR[ 95 ][ 205 ],
   alphaCSR[ 95 ][ 206 ],
   alphaCSR[ 95 ][ 207 ],
   alphaCSR[ 95 ][ 208 ],
   alphaCSR[ 95 ][ 209 ],
   alphaCSR[ 95 ][ 210 ],
   alphaCSR[ 95 ][ 211 ],
   alphaCSR[ 95 ][ 212 ],
   alphaCSR[ 95 ][ 213 ],
   alphaCSR[ 95 ][ 214 ],
   alphaCSR[ 95 ][ 215 ],
   alphaCSR[ 95 ][ 216 ],
   alphaCSR[ 95 ][ 217 ],
   alphaCSR[ 95 ][ 218 ],
   alphaCSR[ 95 ][ 219 ],
   alphaCSR[ 95 ][ 220 ],
   alphaCSR[ 95 ][ 221 ],
   alphaCSR[ 95 ][ 222 ],
   alphaCSR[ 95 ][ 223 ],
   alphaCSR[ 95 ][ 224 ],
   alphaCSR[ 95 ][ 225 ],
   alphaCSR[ 95 ][ 226 ],
   alphaCSR[ 95 ][ 227 ],
   alphaCSR[ 95 ][ 228 ],
   alphaCSR[ 95 ][ 229 ],
   alphaCSR[ 95 ][ 230 ],
   alphaCSR[ 95 ][ 231 ],
   alphaCSR[ 95 ][ 232 ],
   alphaCSR[ 95 ][ 233 ],
   alphaCSR[ 95 ][ 234 ],
   alphaCSR[ 95 ][ 235 ],
   alphaCSR[ 95 ][ 236 ],
   alphaCSR[ 95 ][ 237 ],
   alphaCSR[ 95 ][ 238 ],
   alphaCSR[ 95 ][ 239 ],
   alphaCSR[ 95 ][ 240 ],
   alphaCSR[ 95 ][ 241 ],
   alphaCSR[ 95 ][ 242 ],
   alphaCSR[ 95 ][ 243 ],
   alphaCSR[ 95 ][ 244 ],
   alphaCSR[ 95 ][ 245 ],
   alphaCSR[ 95 ][ 246 ],
   alphaCSR[ 95 ][ 247 ],
   alphaCSR[ 95 ][ 248 ],
   alphaCSR[ 95 ][ 249 ],
   alphaCSR[ 95 ][ 250 ],
   alphaCSR[ 95 ][ 251 ],
   alphaCSR[ 95 ][ 252 ],
   alphaCSR[ 95 ][ 253 ],
   alphaCSR[ 95 ][ 254 ],
   alphaCSR[ 95 ][ 255 ],
   alphaCSR[ 95 ][ 256 ],
   alphaCSR[ 95 ][ 257 ],
   alphaCSR[ 95 ][ 258 ],
   alphaCSR[ 95 ][ 259 ],
   alphaCSR[ 95 ][ 260 ],
   alphaCSR[ 95 ][ 261 ],
   alphaCSR[ 95 ][ 262 ],
   alphaCSR[ 95 ][ 263 ],
   alphaCSR[ 95 ][ 264 ],
   alphaCSR[ 95 ][ 265 ],
   alphaCSR[ 95 ][ 266 ],
   alphaCSR[ 95 ][ 267 ],
   alphaCSR[ 95 ][ 268 ],
   alphaCSR[ 95 ][ 269 ],
   alphaCSR[ 95 ][ 270 ],
   alphaCSR[ 95 ][ 271 ],
   alphaCSR[ 95 ][ 272 ],
   alphaCSR[ 95 ][ 273 ],
   alphaCSR[ 95 ][ 274 ],
   alphaCSR[ 95 ][ 275 ],
   alphaCSR[ 95 ][ 276 ],
   alphaCSR[ 95 ][ 277 ],
   alphaCSR[ 95 ][ 278 ],
   alphaCSR[ 95 ][ 279 ],
   alphaCSR[ 95 ][ 280 ],
   alphaCSR[ 95 ][ 281 ],
   alphaCSR[ 95 ][ 282 ],
   alphaCSR[ 95 ][ 283 ],
   alphaCSR[ 95 ][ 284 ],
   alphaCSR[ 95 ][ 285 ],
   alphaCSR[ 95 ][ 286 ],
   alphaCSR[ 95 ][ 287 ],
   alphaCSR[ 95 ][ 288 ],
   alphaCSR[ 95 ][ 289 ],
   alphaCSR[ 95 ][ 290 ],
   alphaCSR[ 95 ][ 291 ],
   alphaCSR[ 95 ][ 292 ],
   alphaCSR[ 95 ][ 293 ],
   alphaCSR[ 95 ][ 294 ],
   alphaCSR[ 95 ][ 295 ],
   alphaCSR[ 95 ][ 296 ],
   alphaCSR[ 95 ][ 297 ],
   alphaCSR[ 95 ][ 298 ],
   alphaCSR[ 95 ][ 299 ],
   alphaCSR[ 95 ][ 300 ],
   alphaCSR[ 95 ][ 301 ],
   alphaCSR[ 95 ][ 302 ],
   alphaCSR[ 95 ][ 303 ],
   alphaCSR[ 95 ][ 304 ],
   alphaCSR[ 95 ][ 305 ],
   alphaCSR[ 95 ][ 306 ],
   alphaCSR[ 95 ][ 307 ],
   alphaCSR[ 95 ][ 308 ],
   alphaCSR[ 95 ][ 309 ],
   alphaCSR[ 95 ][ 310 ],
   alphaCSR[ 95 ][ 311 ],
   alphaCSR[ 95 ][ 312 ],
   alphaCSR[ 95 ][ 313 ],
   alphaCSR[ 95 ][ 314 ],
   alphaCSR[ 95 ][ 315 ],
   alphaCSR[ 95 ][ 316 ],
   alphaCSR[ 95 ][ 317 ],
   alphaCSR[ 95 ][ 318 ],
   alphaCSR[ 95 ][ 319 ],
   alphaCSR[ 95 ][ 320 ],
   alphaCSR[ 95 ][ 321 ],
   alphaCSR[ 95 ][ 322 ],
   alphaCSR[ 95 ][ 323 ],
   alphaCSR[ 95 ][ 324 ],
   alphaCSR[ 95 ][ 325 ],
   alphaCSR[ 95 ][ 326 ],
   alphaCSR[ 95 ][ 327 ],
   alphaCSR[ 95 ][ 328 ],
   alphaCSR[ 95 ][ 329 ],
   alphaCSR[ 95 ][ 330 ],
   alphaCSR[ 95 ][ 331 ],
   alphaCSR[ 95 ][ 332 ],
   alphaCSR[ 95 ][ 333 ],
   alphaCSR[ 95 ][ 334 ],
   alphaCSR[ 95 ][ 335 ],
   alphaCSR[ 95 ][ 336 ],
   alphaCSR[ 95 ][ 337 ],
   alphaCSR[ 95 ][ 338 ],
   alphaCSR[ 95 ][ 339 ],
   alphaCSR[ 95 ][ 340 ],
   alphaCSR[ 95 ][ 341 ],
   alphaCSR[ 95 ][ 342 ],
   alphaCSR[ 95 ][ 343 ],
   alphaCSR[ 95 ][ 344 ],
   alphaCSR[ 95 ][ 345 ],
   alphaCSR[ 95 ][ 346 ],
   alphaCSR[ 95 ][ 347 ],
   alphaCSR[ 95 ][ 348 ],
   alphaCSR[ 95 ][ 349 ],
   alphaCSR[ 95 ][ 350 ],
   alphaCSR[ 95 ][ 351 ],
   alphaCSR[ 95 ][ 352 ],
   alphaCSR[ 95 ][ 353 ],
   alphaCSR[ 95 ][ 354 ],
   alphaCSR[ 95 ][ 355 ],
   alphaCSR[ 95 ][ 356 ],
   alphaCSR[ 95 ][ 357 ],
   alphaCSR[ 95 ][ 358 ],
   alphaCSR[ 95 ][ 359 ],
   alphaCSR[ 95 ][ 360 ],
   alphaCSR[ 95 ][ 361 ],
   alphaCSR[ 95 ][ 362 ],
   alphaCSR[ 95 ][ 363 ],
   alphaCSR[ 95 ][ 364 ],
   alphaCSR[ 95 ][ 365 ],
   alphaCSR[ 95 ][ 366 ],
   alphaCSR[ 95 ][ 367 ],
   alphaCSR[ 95 ][ 368 ],
   alphaCSR[ 95 ][ 369 ],
   alphaCSR[ 95 ][ 370 ],
   alphaCSR[ 95 ][ 371 ],
   alphaCSR[ 95 ][ 372 ],
   alphaCSR[ 95 ][ 373 ],
   alphaCSR[ 95 ][ 374 ],
   alphaCSR[ 95 ][ 375 ],
   alphaCSR[ 95 ][ 376 ],
   alphaCSR[ 95 ][ 377 ],
   alphaCSR[ 95 ][ 378 ],
   alphaCSR[ 95 ][ 379 ],
   alphaCSR[ 95 ][ 380 ],
   alphaCSR[ 95 ][ 381 ],
   alphaCSR[ 95 ][ 382 ],
   alphaCSR[ 95 ][ 383 ],
   alphaCSR[ 96 ][ 0 ],
   alphaCSR[ 96 ][ 1 ],
   alphaCSR[ 96 ][ 2 ],
   alphaCSR[ 96 ][ 3 ],
   alphaCSR[ 96 ][ 4 ],
   alphaCSR[ 96 ][ 5 ],
   alphaCSR[ 96 ][ 6 ],
   alphaCSR[ 96 ][ 7 ],
   alphaCSR[ 96 ][ 8 ],
   alphaCSR[ 96 ][ 9 ],
   alphaCSR[ 96 ][ 10 ],
   alphaCSR[ 96 ][ 11 ],
   alphaCSR[ 96 ][ 12 ],
   alphaCSR[ 96 ][ 13 ],
   alphaCSR[ 96 ][ 14 ],
   alphaCSR[ 96 ][ 15 ],
   alphaCSR[ 96 ][ 16 ],
   alphaCSR[ 96 ][ 17 ],
   alphaCSR[ 96 ][ 18 ],
   alphaCSR[ 96 ][ 19 ],
   alphaCSR[ 96 ][ 20 ],
   alphaCSR[ 96 ][ 21 ],
   alphaCSR[ 96 ][ 22 ],
   alphaCSR[ 96 ][ 23 ],
   alphaCSR[ 96 ][ 24 ],
   alphaCSR[ 96 ][ 25 ],
   alphaCSR[ 96 ][ 26 ],
   alphaCSR[ 96 ][ 27 ],
   alphaCSR[ 96 ][ 28 ],
   alphaCSR[ 96 ][ 29 ],
   alphaCSR[ 96 ][ 30 ],
   alphaCSR[ 96 ][ 31 ],
   alphaCSR[ 96 ][ 32 ],
   alphaCSR[ 96 ][ 33 ],
   alphaCSR[ 96 ][ 34 ],
   alphaCSR[ 96 ][ 35 ],
   alphaCSR[ 96 ][ 36 ],
   alphaCSR[ 96 ][ 37 ],
   alphaCSR[ 96 ][ 38 ],
   alphaCSR[ 96 ][ 39 ],
   alphaCSR[ 96 ][ 40 ],
   alphaCSR[ 96 ][ 41 ],
   alphaCSR[ 96 ][ 42 ],
   alphaCSR[ 96 ][ 43 ],
   alphaCSR[ 96 ][ 44 ],
   alphaCSR[ 96 ][ 45 ],
   alphaCSR[ 96 ][ 46 ],
   alphaCSR[ 96 ][ 47 ],
   alphaCSR[ 96 ][ 48 ],
   alphaCSR[ 96 ][ 49 ],
   alphaCSR[ 96 ][ 50 ],
   alphaCSR[ 96 ][ 51 ],
   alphaCSR[ 96 ][ 52 ],
   alphaCSR[ 96 ][ 53 ],
   alphaCSR[ 96 ][ 54 ],
   alphaCSR[ 96 ][ 55 ],
   alphaCSR[ 96 ][ 56 ],
   alphaCSR[ 96 ][ 57 ],
   alphaCSR[ 96 ][ 58 ],
   alphaCSR[ 96 ][ 59 ],
   alphaCSR[ 96 ][ 60 ],
   alphaCSR[ 96 ][ 61 ],
   alphaCSR[ 96 ][ 62 ],
   alphaCSR[ 96 ][ 63 ],
   alphaCSR[ 96 ][ 64 ],
   alphaCSR[ 96 ][ 65 ],
   alphaCSR[ 96 ][ 66 ],
   alphaCSR[ 96 ][ 67 ],
   alphaCSR[ 96 ][ 68 ],
   alphaCSR[ 96 ][ 69 ],
   alphaCSR[ 96 ][ 70 ],
   alphaCSR[ 96 ][ 71 ],
   alphaCSR[ 96 ][ 72 ],
   alphaCSR[ 96 ][ 73 ],
   alphaCSR[ 96 ][ 74 ],
   alphaCSR[ 96 ][ 75 ],
   alphaCSR[ 96 ][ 76 ],
   alphaCSR[ 96 ][ 77 ],
   alphaCSR[ 96 ][ 78 ],
   alphaCSR[ 96 ][ 79 ],
   alphaCSR[ 96 ][ 80 ],
   alphaCSR[ 96 ][ 81 ],
   alphaCSR[ 96 ][ 82 ],
   alphaCSR[ 96 ][ 83 ],
   alphaCSR[ 96 ][ 84 ],
   alphaCSR[ 96 ][ 85 ],
   alphaCSR[ 96 ][ 86 ],
   alphaCSR[ 96 ][ 87 ],
   alphaCSR[ 96 ][ 88 ],
   alphaCSR[ 96 ][ 89 ],
   alphaCSR[ 96 ][ 90 ],
   alphaCSR[ 96 ][ 91 ],
   alphaCSR[ 96 ][ 92 ],
   alphaCSR[ 96 ][ 93 ],
   alphaCSR[ 96 ][ 94 ],
   alphaCSR[ 96 ][ 95 ],
   alphaCSR[ 96 ][ 96 ],
   alphaCSR[ 96 ][ 97 ],
   alphaCSR[ 96 ][ 98 ],
   alphaCSR[ 96 ][ 99 ],
   alphaCSR[ 96 ][ 100 ],
   alphaCSR[ 96 ][ 101 ],
   alphaCSR[ 96 ][ 102 ],
   alphaCSR[ 96 ][ 103 ],
   alphaCSR[ 96 ][ 104 ],
   alphaCSR[ 96 ][ 105 ],
   alphaCSR[ 96 ][ 106 ],
   alphaCSR[ 96 ][ 107 ],
   alphaCSR[ 96 ][ 108 ],
   alphaCSR[ 96 ][ 109 ],
   alphaCSR[ 96 ][ 110 ],
   alphaCSR[ 96 ][ 111 ],
   alphaCSR[ 96 ][ 112 ],
   alphaCSR[ 96 ][ 113 ],
   alphaCSR[ 96 ][ 114 ],
   alphaCSR[ 96 ][ 115 ],
   alphaCSR[ 96 ][ 116 ],
   alphaCSR[ 96 ][ 117 ],
   alphaCSR[ 96 ][ 118 ],
   alphaCSR[ 96 ][ 119 ],
   alphaCSR[ 96 ][ 120 ],
   alphaCSR[ 96 ][ 121 ],
   alphaCSR[ 96 ][ 122 ],
   alphaCSR[ 96 ][ 123 ],
   alphaCSR[ 96 ][ 124 ],
   alphaCSR[ 96 ][ 125 ],
   alphaCSR[ 96 ][ 126 ],
   alphaCSR[ 96 ][ 127 ],
   alphaCSR[ 96 ][ 128 ],
   alphaCSR[ 96 ][ 129 ],
   alphaCSR[ 96 ][ 130 ],
   alphaCSR[ 96 ][ 131 ],
   alphaCSR[ 96 ][ 132 ],
   alphaCSR[ 96 ][ 133 ],
   alphaCSR[ 96 ][ 134 ],
   alphaCSR[ 96 ][ 135 ],
   alphaCSR[ 96 ][ 136 ],
   alphaCSR[ 96 ][ 137 ],
   alphaCSR[ 96 ][ 138 ],
   alphaCSR[ 96 ][ 139 ],
   alphaCSR[ 96 ][ 140 ],
   alphaCSR[ 96 ][ 141 ],
   alphaCSR[ 96 ][ 142 ],
   alphaCSR[ 96 ][ 143 ],
   alphaCSR[ 96 ][ 144 ],
   alphaCSR[ 96 ][ 145 ],
   alphaCSR[ 96 ][ 146 ],
   alphaCSR[ 96 ][ 147 ],
   alphaCSR[ 96 ][ 148 ],
   alphaCSR[ 96 ][ 149 ],
   alphaCSR[ 96 ][ 150 ],
   alphaCSR[ 96 ][ 151 ],
   alphaCSR[ 96 ][ 152 ],
   alphaCSR[ 96 ][ 153 ],
   alphaCSR[ 96 ][ 154 ],
   alphaCSR[ 96 ][ 155 ],
   alphaCSR[ 96 ][ 156 ],
   alphaCSR[ 96 ][ 157 ],
   alphaCSR[ 96 ][ 158 ],
   alphaCSR[ 96 ][ 159 ],
   alphaCSR[ 96 ][ 160 ],
   alphaCSR[ 96 ][ 161 ],
   alphaCSR[ 96 ][ 162 ],
   alphaCSR[ 96 ][ 163 ],
   alphaCSR[ 96 ][ 164 ],
   alphaCSR[ 96 ][ 165 ],
   alphaCSR[ 96 ][ 166 ],
   alphaCSR[ 96 ][ 167 ],
   alphaCSR[ 96 ][ 168 ],
   alphaCSR[ 96 ][ 169 ],
   alphaCSR[ 96 ][ 170 ],
   alphaCSR[ 96 ][ 171 ],
   alphaCSR[ 96 ][ 172 ],
   alphaCSR[ 96 ][ 173 ],
   alphaCSR[ 96 ][ 174 ],
   alphaCSR[ 96 ][ 175 ],
   alphaCSR[ 96 ][ 176 ],
   alphaCSR[ 96 ][ 177 ],
   alphaCSR[ 96 ][ 178 ],
   alphaCSR[ 96 ][ 179 ],
   alphaCSR[ 96 ][ 180 ],
   alphaCSR[ 96 ][ 181 ],
   alphaCSR[ 96 ][ 182 ],
   alphaCSR[ 96 ][ 183 ],
   alphaCSR[ 96 ][ 184 ],
   alphaCSR[ 96 ][ 185 ],
   alphaCSR[ 96 ][ 186 ],
   alphaCSR[ 96 ][ 187 ],
   alphaCSR[ 96 ][ 188 ],
   alphaCSR[ 96 ][ 189 ],
   alphaCSR[ 96 ][ 190 ],
   alphaCSR[ 96 ][ 191 ],
   alphaCSR[ 96 ][ 192 ],
   alphaCSR[ 96 ][ 193 ],
   alphaCSR[ 96 ][ 194 ],
   alphaCSR[ 96 ][ 195 ],
   alphaCSR[ 96 ][ 196 ],
   alphaCSR[ 96 ][ 197 ],
   alphaCSR[ 96 ][ 198 ],
   alphaCSR[ 96 ][ 199 ],
   alphaCSR[ 96 ][ 200 ],
   alphaCSR[ 96 ][ 201 ],
   alphaCSR[ 96 ][ 202 ],
   alphaCSR[ 96 ][ 203 ],
   alphaCSR[ 96 ][ 204 ],
   alphaCSR[ 96 ][ 205 ],
   alphaCSR[ 96 ][ 206 ],
   alphaCSR[ 96 ][ 207 ],
   alphaCSR[ 96 ][ 208 ],
   alphaCSR[ 96 ][ 209 ],
   alphaCSR[ 96 ][ 210 ],
   alphaCSR[ 96 ][ 211 ],
   alphaCSR[ 96 ][ 212 ],
   alphaCSR[ 96 ][ 213 ],
   alphaCSR[ 96 ][ 214 ],
   alphaCSR[ 96 ][ 215 ],
   alphaCSR[ 96 ][ 216 ],
   alphaCSR[ 96 ][ 217 ],
   alphaCSR[ 96 ][ 218 ],
   alphaCSR[ 96 ][ 219 ],
   alphaCSR[ 96 ][ 220 ],
   alphaCSR[ 96 ][ 221 ],
   alphaCSR[ 96 ][ 222 ],
   alphaCSR[ 96 ][ 223 ],
   alphaCSR[ 96 ][ 224 ],
   alphaCSR[ 96 ][ 225 ],
   alphaCSR[ 96 ][ 226 ],
   alphaCSR[ 96 ][ 227 ],
   alphaCSR[ 96 ][ 228 ],
   alphaCSR[ 96 ][ 229 ],
   alphaCSR[ 96 ][ 230 ],
   alphaCSR[ 96 ][ 231 ],
   alphaCSR[ 96 ][ 232 ],
   alphaCSR[ 96 ][ 233 ],
   alphaCSR[ 96 ][ 234 ],
   alphaCSR[ 96 ][ 235 ],
   alphaCSR[ 96 ][ 236 ],
   alphaCSR[ 96 ][ 237 ],
   alphaCSR[ 96 ][ 238 ],
   alphaCSR[ 96 ][ 239 ],
   alphaCSR[ 96 ][ 240 ],
   alphaCSR[ 96 ][ 241 ],
   alphaCSR[ 96 ][ 242 ],
   alphaCSR[ 96 ][ 243 ],
   alphaCSR[ 96 ][ 244 ],
   alphaCSR[ 96 ][ 245 ],
   alphaCSR[ 96 ][ 246 ],
   alphaCSR[ 96 ][ 247 ],
   alphaCSR[ 96 ][ 248 ],
   alphaCSR[ 96 ][ 249 ],
   alphaCSR[ 96 ][ 250 ],
   alphaCSR[ 96 ][ 251 ],
   alphaCSR[ 96 ][ 252 ],
   alphaCSR[ 96 ][ 253 ],
   alphaCSR[ 96 ][ 254 ],
   alphaCSR[ 96 ][ 255 ],
   alphaCSR[ 96 ][ 256 ],
   alphaCSR[ 96 ][ 257 ],
   alphaCSR[ 96 ][ 258 ],
   alphaCSR[ 96 ][ 259 ],
   alphaCSR[ 96 ][ 260 ],
   alphaCSR[ 96 ][ 261 ],
   alphaCSR[ 96 ][ 262 ],
   alphaCSR[ 96 ][ 263 ],
   alphaCSR[ 96 ][ 264 ],
   alphaCSR[ 96 ][ 265 ],
   alphaCSR[ 96 ][ 266 ],
   alphaCSR[ 96 ][ 267 ],
   alphaCSR[ 96 ][ 268 ],
   alphaCSR[ 96 ][ 269 ],
   alphaCSR[ 96 ][ 270 ],
   alphaCSR[ 96 ][ 271 ],
   alphaCSR[ 96 ][ 272 ],
   alphaCSR[ 96 ][ 273 ],
   alphaCSR[ 96 ][ 274 ],
   alphaCSR[ 96 ][ 275 ],
   alphaCSR[ 96 ][ 276 ],
   alphaCSR[ 96 ][ 277 ],
   alphaCSR[ 96 ][ 278 ],
   alphaCSR[ 96 ][ 279 ],
   alphaCSR[ 96 ][ 280 ],
   alphaCSR[ 96 ][ 281 ],
   alphaCSR[ 96 ][ 282 ],
   alphaCSR[ 96 ][ 283 ],
   alphaCSR[ 96 ][ 284 ],
   alphaCSR[ 96 ][ 285 ],
   alphaCSR[ 96 ][ 286 ],
   alphaCSR[ 96 ][ 287 ],
   alphaCSR[ 96 ][ 288 ],
   alphaCSR[ 96 ][ 289 ],
   alphaCSR[ 96 ][ 290 ],
   alphaCSR[ 96 ][ 291 ],
   alphaCSR[ 96 ][ 292 ],
   alphaCSR[ 96 ][ 293 ],
   alphaCSR[ 96 ][ 294 ],
   alphaCSR[ 96 ][ 295 ],
   alphaCSR[ 96 ][ 296 ],
   alphaCSR[ 96 ][ 297 ],
   alphaCSR[ 96 ][ 298 ],
   alphaCSR[ 96 ][ 299 ],
   alphaCSR[ 96 ][ 300 ],
   alphaCSR[ 96 ][ 301 ],
   alphaCSR[ 96 ][ 302 ],
   alphaCSR[ 96 ][ 303 ],
   alphaCSR[ 96 ][ 304 ],
   alphaCSR[ 96 ][ 305 ],
   alphaCSR[ 96 ][ 306 ],
   alphaCSR[ 96 ][ 307 ],
   alphaCSR[ 96 ][ 308 ],
   alphaCSR[ 96 ][ 309 ],
   alphaCSR[ 96 ][ 310 ],
   alphaCSR[ 96 ][ 311 ],
   alphaCSR[ 96 ][ 312 ],
   alphaCSR[ 96 ][ 313 ],
   alphaCSR[ 96 ][ 314 ],
   alphaCSR[ 96 ][ 315 ],
   alphaCSR[ 96 ][ 316 ],
   alphaCSR[ 96 ][ 317 ],
   alphaCSR[ 96 ][ 318 ],
   alphaCSR[ 96 ][ 319 ],
   alphaCSR[ 96 ][ 320 ],
   alphaCSR[ 96 ][ 321 ],
   alphaCSR[ 96 ][ 322 ],
   alphaCSR[ 96 ][ 323 ],
   alphaCSR[ 96 ][ 324 ],
   alphaCSR[ 96 ][ 325 ],
   alphaCSR[ 96 ][ 326 ],
   alphaCSR[ 96 ][ 327 ],
   alphaCSR[ 96 ][ 328 ],
   alphaCSR[ 96 ][ 329 ],
   alphaCSR[ 96 ][ 330 ],
   alphaCSR[ 96 ][ 331 ],
   alphaCSR[ 96 ][ 332 ],
   alphaCSR[ 96 ][ 333 ],
   alphaCSR[ 96 ][ 334 ],
   alphaCSR[ 96 ][ 335 ],
   alphaCSR[ 96 ][ 336 ],
   alphaCSR[ 96 ][ 337 ],
   alphaCSR[ 96 ][ 338 ],
   alphaCSR[ 96 ][ 339 ],
   alphaCSR[ 96 ][ 340 ],
   alphaCSR[ 96 ][ 341 ],
   alphaCSR[ 96 ][ 342 ],
   alphaCSR[ 96 ][ 343 ],
   alphaCSR[ 96 ][ 344 ],
   alphaCSR[ 96 ][ 345 ],
   alphaCSR[ 96 ][ 346 ],
   alphaCSR[ 96 ][ 347 ],
   alphaCSR[ 96 ][ 348 ],
   alphaCSR[ 96 ][ 349 ],
   alphaCSR[ 96 ][ 350 ],
   alphaCSR[ 96 ][ 351 ],
   alphaCSR[ 96 ][ 352 ],
   alphaCSR[ 96 ][ 353 ],
   alphaCSR[ 96 ][ 354 ],
   alphaCSR[ 96 ][ 355 ],
   alphaCSR[ 96 ][ 356 ],
   alphaCSR[ 96 ][ 357 ],
   alphaCSR[ 96 ][ 358 ],
   alphaCSR[ 96 ][ 359 ],
   alphaCSR[ 96 ][ 360 ],
   alphaCSR[ 96 ][ 361 ],
   alphaCSR[ 96 ][ 362 ],
   alphaCSR[ 96 ][ 363 ],
   alphaCSR[ 96 ][ 364 ],
   alphaCSR[ 96 ][ 365 ],
   alphaCSR[ 96 ][ 366 ],
   alphaCSR[ 96 ][ 367 ],
   alphaCSR[ 96 ][ 368 ],
   alphaCSR[ 96 ][ 369 ],
   alphaCSR[ 96 ][ 370 ],
   alphaCSR[ 96 ][ 371 ],
   alphaCSR[ 96 ][ 372 ],
   alphaCSR[ 96 ][ 373 ],
   alphaCSR[ 96 ][ 374 ],
   alphaCSR[ 96 ][ 375 ],
   alphaCSR[ 96 ][ 376 ],
   alphaCSR[ 96 ][ 377 ],
   alphaCSR[ 96 ][ 378 ],
   alphaCSR[ 96 ][ 379 ],
   alphaCSR[ 96 ][ 380 ],
   alphaCSR[ 96 ][ 381 ],
   alphaCSR[ 96 ][ 382 ],
   alphaCSR[ 96 ][ 383 ],
   alphaCSR[ 97 ][ 0 ],
   alphaCSR[ 97 ][ 1 ],
   alphaCSR[ 97 ][ 2 ],
   alphaCSR[ 97 ][ 3 ],
   alphaCSR[ 97 ][ 4 ],
   alphaCSR[ 97 ][ 5 ],
   alphaCSR[ 97 ][ 6 ],
   alphaCSR[ 97 ][ 7 ],
   alphaCSR[ 97 ][ 8 ],
   alphaCSR[ 97 ][ 9 ],
   alphaCSR[ 97 ][ 10 ],
   alphaCSR[ 97 ][ 11 ],
   alphaCSR[ 97 ][ 12 ],
   alphaCSR[ 97 ][ 13 ],
   alphaCSR[ 97 ][ 14 ],
   alphaCSR[ 97 ][ 15 ],
   alphaCSR[ 97 ][ 16 ],
   alphaCSR[ 97 ][ 17 ],
   alphaCSR[ 97 ][ 18 ],
   alphaCSR[ 97 ][ 19 ],
   alphaCSR[ 97 ][ 20 ],
   alphaCSR[ 97 ][ 21 ],
   alphaCSR[ 97 ][ 22 ],
   alphaCSR[ 97 ][ 23 ],
   alphaCSR[ 97 ][ 24 ],
   alphaCSR[ 97 ][ 25 ],
   alphaCSR[ 97 ][ 26 ],
   alphaCSR[ 97 ][ 27 ],
   alphaCSR[ 97 ][ 28 ],
   alphaCSR[ 97 ][ 29 ],
   alphaCSR[ 97 ][ 30 ],
   alphaCSR[ 97 ][ 31 ],
   alphaCSR[ 97 ][ 32 ],
   alphaCSR[ 97 ][ 33 ],
   alphaCSR[ 97 ][ 34 ],
   alphaCSR[ 97 ][ 35 ],
   alphaCSR[ 97 ][ 36 ],
   alphaCSR[ 97 ][ 37 ],
   alphaCSR[ 97 ][ 38 ],
   alphaCSR[ 97 ][ 39 ],
   alphaCSR[ 97 ][ 40 ],
   alphaCSR[ 97 ][ 41 ],
   alphaCSR[ 97 ][ 42 ],
   alphaCSR[ 97 ][ 43 ],
   alphaCSR[ 97 ][ 44 ],
   alphaCSR[ 97 ][ 45 ],
   alphaCSR[ 97 ][ 46 ],
   alphaCSR[ 97 ][ 47 ],
   alphaCSR[ 97 ][ 48 ],
   alphaCSR[ 97 ][ 49 ],
   alphaCSR[ 97 ][ 50 ],
   alphaCSR[ 97 ][ 51 ],
   alphaCSR[ 97 ][ 52 ],
   alphaCSR[ 97 ][ 53 ],
   alphaCSR[ 97 ][ 54 ],
   alphaCSR[ 97 ][ 55 ],
   alphaCSR[ 97 ][ 56 ],
   alphaCSR[ 97 ][ 57 ],
   alphaCSR[ 97 ][ 58 ],
   alphaCSR[ 97 ][ 59 ],
   alphaCSR[ 97 ][ 60 ],
   alphaCSR[ 97 ][ 61 ],
   alphaCSR[ 97 ][ 62 ],
   alphaCSR[ 97 ][ 63 ],
   alphaCSR[ 97 ][ 64 ],
   alphaCSR[ 97 ][ 65 ],
   alphaCSR[ 97 ][ 66 ],
   alphaCSR[ 97 ][ 67 ],
   alphaCSR[ 97 ][ 68 ],
   alphaCSR[ 97 ][ 69 ],
   alphaCSR[ 97 ][ 70 ],
   alphaCSR[ 97 ][ 71 ],
   alphaCSR[ 97 ][ 72 ],
   alphaCSR[ 97 ][ 73 ],
   alphaCSR[ 97 ][ 74 ],
   alphaCSR[ 97 ][ 75 ],
   alphaCSR[ 97 ][ 76 ],
   alphaCSR[ 97 ][ 77 ],
   alphaCSR[ 97 ][ 78 ],
   alphaCSR[ 97 ][ 79 ],
   alphaCSR[ 97 ][ 80 ],
   alphaCSR[ 97 ][ 81 ],
   alphaCSR[ 97 ][ 82 ],
   alphaCSR[ 97 ][ 83 ],
   alphaCSR[ 97 ][ 84 ],
   alphaCSR[ 97 ][ 85 ],
   alphaCSR[ 97 ][ 86 ],
   alphaCSR[ 97 ][ 87 ],
   alphaCSR[ 97 ][ 88 ],
   alphaCSR[ 97 ][ 89 ],
   alphaCSR[ 97 ][ 90 ],
   alphaCSR[ 97 ][ 91 ],
   alphaCSR[ 97 ][ 92 ],
   alphaCSR[ 97 ][ 93 ],
   alphaCSR[ 97 ][ 94 ],
   alphaCSR[ 97 ][ 95 ],
   alphaCSR[ 97 ][ 96 ],
   alphaCSR[ 97 ][ 97 ],
   alphaCSR[ 97 ][ 98 ],
   alphaCSR[ 97 ][ 99 ],
   alphaCSR[ 97 ][ 100 ],
   alphaCSR[ 97 ][ 101 ],
   alphaCSR[ 97 ][ 102 ],
   alphaCSR[ 97 ][ 103 ],
   alphaCSR[ 97 ][ 104 ],
   alphaCSR[ 97 ][ 105 ],
   alphaCSR[ 97 ][ 106 ],
   alphaCSR[ 97 ][ 107 ],
   alphaCSR[ 97 ][ 108 ],
   alphaCSR[ 97 ][ 109 ],
   alphaCSR[ 97 ][ 110 ],
   alphaCSR[ 97 ][ 111 ],
   alphaCSR[ 97 ][ 112 ],
   alphaCSR[ 97 ][ 113 ],
   alphaCSR[ 97 ][ 114 ],
   alphaCSR[ 97 ][ 115 ],
   alphaCSR[ 97 ][ 116 ],
   alphaCSR[ 97 ][ 117 ],
   alphaCSR[ 97 ][ 118 ],
   alphaCSR[ 97 ][ 119 ],
   alphaCSR[ 97 ][ 120 ],
   alphaCSR[ 97 ][ 121 ],
   alphaCSR[ 97 ][ 122 ],
   alphaCSR[ 97 ][ 123 ],
   alphaCSR[ 97 ][ 124 ],
   alphaCSR[ 97 ][ 125 ],
   alphaCSR[ 97 ][ 126 ],
   alphaCSR[ 97 ][ 127 ],
   alphaCSR[ 97 ][ 128 ],
   alphaCSR[ 97 ][ 129 ],
   alphaCSR[ 97 ][ 130 ],
   alphaCSR[ 97 ][ 131 ],
   alphaCSR[ 97 ][ 132 ],
   alphaCSR[ 97 ][ 133 ],
   alphaCSR[ 97 ][ 134 ],
   alphaCSR[ 97 ][ 135 ],
   alphaCSR[ 97 ][ 136 ],
   alphaCSR[ 97 ][ 137 ],
   alphaCSR[ 97 ][ 138 ],
   alphaCSR[ 97 ][ 139 ],
   alphaCSR[ 97 ][ 140 ],
   alphaCSR[ 97 ][ 141 ],
   alphaCSR[ 97 ][ 142 ],
   alphaCSR[ 97 ][ 143 ],
   alphaCSR[ 97 ][ 144 ],
   alphaCSR[ 97 ][ 145 ],
   alphaCSR[ 97 ][ 146 ],
   alphaCSR[ 97 ][ 147 ],
   alphaCSR[ 97 ][ 148 ],
   alphaCSR[ 97 ][ 149 ],
   alphaCSR[ 97 ][ 150 ],
   alphaCSR[ 97 ][ 151 ],
   alphaCSR[ 97 ][ 152 ],
   alphaCSR[ 97 ][ 153 ],
   alphaCSR[ 97 ][ 154 ],
   alphaCSR[ 97 ][ 155 ],
   alphaCSR[ 97 ][ 156 ],
   alphaCSR[ 97 ][ 157 ],
   alphaCSR[ 97 ][ 158 ],
   alphaCSR[ 97 ][ 159 ],
   alphaCSR[ 97 ][ 160 ],
   alphaCSR[ 97 ][ 161 ],
   alphaCSR[ 97 ][ 162 ],
   alphaCSR[ 97 ][ 163 ],
   alphaCSR[ 97 ][ 164 ],
   alphaCSR[ 97 ][ 165 ],
   alphaCSR[ 97 ][ 166 ],
   alphaCSR[ 97 ][ 167 ],
   alphaCSR[ 97 ][ 168 ],
   alphaCSR[ 97 ][ 169 ],
   alphaCSR[ 97 ][ 170 ],
   alphaCSR[ 97 ][ 171 ],
   alphaCSR[ 97 ][ 172 ],
   alphaCSR[ 97 ][ 173 ],
   alphaCSR[ 97 ][ 174 ],
   alphaCSR[ 97 ][ 175 ],
   alphaCSR[ 97 ][ 176 ],
   alphaCSR[ 97 ][ 177 ],
   alphaCSR[ 97 ][ 178 ],
   alphaCSR[ 97 ][ 179 ],
   alphaCSR[ 97 ][ 180 ],
   alphaCSR[ 97 ][ 181 ],
   alphaCSR[ 97 ][ 182 ],
   alphaCSR[ 97 ][ 183 ],
   alphaCSR[ 97 ][ 184 ],
   alphaCSR[ 97 ][ 185 ],
   alphaCSR[ 97 ][ 186 ],
   alphaCSR[ 97 ][ 187 ],
   alphaCSR[ 97 ][ 188 ],
   alphaCSR[ 97 ][ 189 ],
   alphaCSR[ 97 ][ 190 ],
   alphaCSR[ 97 ][ 191 ],
   alphaCSR[ 97 ][ 192 ],
   alphaCSR[ 97 ][ 193 ],
   alphaCSR[ 97 ][ 194 ],
   alphaCSR[ 97 ][ 195 ],
   alphaCSR[ 97 ][ 196 ],
   alphaCSR[ 97 ][ 197 ],
   alphaCSR[ 97 ][ 198 ],
   alphaCSR[ 97 ][ 199 ],
   alphaCSR[ 97 ][ 200 ],
   alphaCSR[ 97 ][ 201 ],
   alphaCSR[ 97 ][ 202 ],
   alphaCSR[ 97 ][ 203 ],
   alphaCSR[ 97 ][ 204 ],
   alphaCSR[ 97 ][ 205 ],
   alphaCSR[ 97 ][ 206 ],
   alphaCSR[ 97 ][ 207 ],
   alphaCSR[ 97 ][ 208 ],
   alphaCSR[ 97 ][ 209 ],
   alphaCSR[ 97 ][ 210 ],
   alphaCSR[ 97 ][ 211 ],
   alphaCSR[ 97 ][ 212 ],
   alphaCSR[ 97 ][ 213 ],
   alphaCSR[ 97 ][ 214 ],
   alphaCSR[ 97 ][ 215 ],
   alphaCSR[ 97 ][ 216 ],
   alphaCSR[ 97 ][ 217 ],
   alphaCSR[ 97 ][ 218 ],
   alphaCSR[ 97 ][ 219 ],
   alphaCSR[ 97 ][ 220 ],
   alphaCSR[ 97 ][ 221 ],
   alphaCSR[ 97 ][ 222 ],
   alphaCSR[ 97 ][ 223 ],
   alphaCSR[ 97 ][ 224 ],
   alphaCSR[ 97 ][ 225 ],
   alphaCSR[ 97 ][ 226 ],
   alphaCSR[ 97 ][ 227 ],
   alphaCSR[ 97 ][ 228 ],
   alphaCSR[ 97 ][ 229 ],
   alphaCSR[ 97 ][ 230 ],
   alphaCSR[ 97 ][ 231 ],
   alphaCSR[ 97 ][ 232 ],
   alphaCSR[ 97 ][ 233 ],
   alphaCSR[ 97 ][ 234 ],
   alphaCSR[ 97 ][ 235 ],
   alphaCSR[ 97 ][ 236 ],
   alphaCSR[ 97 ][ 237 ],
   alphaCSR[ 97 ][ 238 ],
   alphaCSR[ 97 ][ 239 ],
   alphaCSR[ 97 ][ 240 ],
   alphaCSR[ 97 ][ 241 ],
   alphaCSR[ 97 ][ 242 ],
   alphaCSR[ 97 ][ 243 ],
   alphaCSR[ 97 ][ 244 ],
   alphaCSR[ 97 ][ 245 ],
   alphaCSR[ 97 ][ 246 ],
   alphaCSR[ 97 ][ 247 ],
   alphaCSR[ 97 ][ 248 ],
   alphaCSR[ 97 ][ 249 ],
   alphaCSR[ 97 ][ 250 ],
   alphaCSR[ 97 ][ 251 ],
   alphaCSR[ 97 ][ 252 ],
   alphaCSR[ 97 ][ 253 ],
   alphaCSR[ 97 ][ 254 ],
   alphaCSR[ 97 ][ 255 ],
   alphaCSR[ 97 ][ 256 ],
   alphaCSR[ 97 ][ 257 ],
   alphaCSR[ 97 ][ 258 ],
   alphaCSR[ 97 ][ 259 ],
   alphaCSR[ 97 ][ 260 ],
   alphaCSR[ 97 ][ 261 ],
   alphaCSR[ 97 ][ 262 ],
   alphaCSR[ 97 ][ 263 ],
   alphaCSR[ 97 ][ 264 ],
   alphaCSR[ 97 ][ 265 ],
   alphaCSR[ 97 ][ 266 ],
   alphaCSR[ 97 ][ 267 ],
   alphaCSR[ 97 ][ 268 ],
   alphaCSR[ 97 ][ 269 ],
   alphaCSR[ 97 ][ 270 ],
   alphaCSR[ 97 ][ 271 ],
   alphaCSR[ 97 ][ 272 ],
   alphaCSR[ 97 ][ 273 ],
   alphaCSR[ 97 ][ 274 ],
   alphaCSR[ 97 ][ 275 ],
   alphaCSR[ 97 ][ 276 ],
   alphaCSR[ 97 ][ 277 ],
   alphaCSR[ 97 ][ 278 ],
   alphaCSR[ 97 ][ 279 ],
   alphaCSR[ 97 ][ 280 ],
   alphaCSR[ 97 ][ 281 ],
   alphaCSR[ 97 ][ 282 ],
   alphaCSR[ 97 ][ 283 ],
   alphaCSR[ 97 ][ 284 ],
   alphaCSR[ 97 ][ 285 ],
   alphaCSR[ 97 ][ 286 ],
   alphaCSR[ 97 ][ 287 ],
   alphaCSR[ 97 ][ 288 ],
   alphaCSR[ 97 ][ 289 ],
   alphaCSR[ 97 ][ 290 ],
   alphaCSR[ 97 ][ 291 ],
   alphaCSR[ 97 ][ 292 ],
   alphaCSR[ 97 ][ 293 ],
   alphaCSR[ 97 ][ 294 ],
   alphaCSR[ 97 ][ 295 ],
   alphaCSR[ 97 ][ 296 ],
   alphaCSR[ 97 ][ 297 ],
   alphaCSR[ 97 ][ 298 ],
   alphaCSR[ 97 ][ 299 ],
   alphaCSR[ 97 ][ 300 ],
   alphaCSR[ 97 ][ 301 ],
   alphaCSR[ 97 ][ 302 ],
   alphaCSR[ 97 ][ 303 ],
   alphaCSR[ 97 ][ 304 ],
   alphaCSR[ 97 ][ 305 ],
   alphaCSR[ 97 ][ 306 ],
   alphaCSR[ 97 ][ 307 ],
   alphaCSR[ 97 ][ 308 ],
   alphaCSR[ 97 ][ 309 ],
   alphaCSR[ 97 ][ 310 ],
   alphaCSR[ 97 ][ 311 ],
   alphaCSR[ 97 ][ 312 ],
   alphaCSR[ 97 ][ 313 ],
   alphaCSR[ 97 ][ 314 ],
   alphaCSR[ 97 ][ 315 ],
   alphaCSR[ 97 ][ 316 ],
   alphaCSR[ 97 ][ 317 ],
   alphaCSR[ 97 ][ 318 ],
   alphaCSR[ 97 ][ 319 ],
   alphaCSR[ 97 ][ 320 ],
   alphaCSR[ 97 ][ 321 ],
   alphaCSR[ 97 ][ 322 ],
   alphaCSR[ 97 ][ 323 ],
   alphaCSR[ 97 ][ 324 ],
   alphaCSR[ 97 ][ 325 ],
   alphaCSR[ 97 ][ 326 ],
   alphaCSR[ 97 ][ 327 ],
   alphaCSR[ 97 ][ 328 ],
   alphaCSR[ 97 ][ 329 ],
   alphaCSR[ 97 ][ 330 ],
   alphaCSR[ 97 ][ 331 ],
   alphaCSR[ 97 ][ 332 ],
   alphaCSR[ 97 ][ 333 ],
   alphaCSR[ 97 ][ 334 ],
   alphaCSR[ 97 ][ 335 ],
   alphaCSR[ 97 ][ 336 ],
   alphaCSR[ 97 ][ 337 ],
   alphaCSR[ 97 ][ 338 ],
   alphaCSR[ 97 ][ 339 ],
   alphaCSR[ 97 ][ 340 ],
   alphaCSR[ 97 ][ 341 ],
   alphaCSR[ 97 ][ 342 ],
   alphaCSR[ 97 ][ 343 ],
   alphaCSR[ 97 ][ 344 ],
   alphaCSR[ 97 ][ 345 ],
   alphaCSR[ 97 ][ 346 ],
   alphaCSR[ 97 ][ 347 ],
   alphaCSR[ 97 ][ 348 ],
   alphaCSR[ 97 ][ 349 ],
   alphaCSR[ 97 ][ 350 ],
   alphaCSR[ 97 ][ 351 ],
   alphaCSR[ 97 ][ 352 ],
   alphaCSR[ 97 ][ 353 ],
   alphaCSR[ 97 ][ 354 ],
   alphaCSR[ 97 ][ 355 ],
   alphaCSR[ 97 ][ 356 ],
   alphaCSR[ 97 ][ 357 ],
   alphaCSR[ 97 ][ 358 ],
   alphaCSR[ 97 ][ 359 ],
   alphaCSR[ 97 ][ 360 ],
   alphaCSR[ 97 ][ 361 ],
   alphaCSR[ 97 ][ 362 ],
   alphaCSR[ 97 ][ 363 ],
   alphaCSR[ 97 ][ 364 ],
   alphaCSR[ 97 ][ 365 ],
   alphaCSR[ 97 ][ 366 ],
   alphaCSR[ 97 ][ 367 ],
   alphaCSR[ 97 ][ 368 ],
   alphaCSR[ 97 ][ 369 ],
   alphaCSR[ 97 ][ 370 ],
   alphaCSR[ 97 ][ 371 ],
   alphaCSR[ 97 ][ 372 ],
   alphaCSR[ 97 ][ 373 ],
   alphaCSR[ 97 ][ 374 ],
   alphaCSR[ 97 ][ 375 ],
   alphaCSR[ 97 ][ 376 ],
   alphaCSR[ 97 ][ 377 ],
   alphaCSR[ 97 ][ 378 ],
   alphaCSR[ 97 ][ 379 ],
   alphaCSR[ 97 ][ 380 ],
   alphaCSR[ 97 ][ 381 ],
   alphaCSR[ 97 ][ 382 ],
   alphaCSR[ 97 ][ 383 ],
   alphaCSR[ 98 ][ 0 ],
   alphaCSR[ 98 ][ 1 ],
   alphaCSR[ 98 ][ 2 ],
   alphaCSR[ 98 ][ 3 ],
   alphaCSR[ 98 ][ 4 ],
   alphaCSR[ 98 ][ 5 ],
   alphaCSR[ 98 ][ 6 ],
   alphaCSR[ 98 ][ 7 ],
   alphaCSR[ 98 ][ 8 ],
   alphaCSR[ 98 ][ 9 ],
   alphaCSR[ 98 ][ 10 ],
   alphaCSR[ 98 ][ 11 ],
   alphaCSR[ 98 ][ 12 ],
   alphaCSR[ 98 ][ 13 ],
   alphaCSR[ 98 ][ 14 ],
   alphaCSR[ 98 ][ 15 ],
   alphaCSR[ 98 ][ 16 ],
   alphaCSR[ 98 ][ 17 ],
   alphaCSR[ 98 ][ 18 ],
   alphaCSR[ 98 ][ 19 ],
   alphaCSR[ 98 ][ 20 ],
   alphaCSR[ 98 ][ 21 ],
   alphaCSR[ 98 ][ 22 ],
   alphaCSR[ 98 ][ 23 ],
   alphaCSR[ 98 ][ 24 ],
   alphaCSR[ 98 ][ 25 ],
   alphaCSR[ 98 ][ 26 ],
   alphaCSR[ 98 ][ 27 ],
   alphaCSR[ 98 ][ 28 ],
   alphaCSR[ 98 ][ 29 ],
   alphaCSR[ 98 ][ 30 ],
   alphaCSR[ 98 ][ 31 ],
   alphaCSR[ 98 ][ 32 ],
   alphaCSR[ 98 ][ 33 ],
   alphaCSR[ 98 ][ 34 ],
   alphaCSR[ 98 ][ 35 ],
   alphaCSR[ 98 ][ 36 ],
   alphaCSR[ 98 ][ 37 ],
   alphaCSR[ 98 ][ 38 ],
   alphaCSR[ 98 ][ 39 ],
   alphaCSR[ 98 ][ 40 ],
   alphaCSR[ 98 ][ 41 ],
   alphaCSR[ 98 ][ 42 ],
   alphaCSR[ 98 ][ 43 ],
   alphaCSR[ 98 ][ 44 ],
   alphaCSR[ 98 ][ 45 ],
   alphaCSR[ 98 ][ 46 ],
   alphaCSR[ 98 ][ 47 ],
   alphaCSR[ 98 ][ 48 ],
   alphaCSR[ 98 ][ 49 ],
   alphaCSR[ 98 ][ 50 ],
   alphaCSR[ 98 ][ 51 ],
   alphaCSR[ 98 ][ 52 ],
   alphaCSR[ 98 ][ 53 ],
   alphaCSR[ 98 ][ 54 ],
   alphaCSR[ 98 ][ 55 ],
   alphaCSR[ 98 ][ 56 ],
   alphaCSR[ 98 ][ 57 ],
   alphaCSR[ 98 ][ 58 ],
   alphaCSR[ 98 ][ 59 ],
   alphaCSR[ 98 ][ 60 ],
   alphaCSR[ 98 ][ 61 ],
   alphaCSR[ 98 ][ 62 ],
   alphaCSR[ 98 ][ 63 ],
   alphaCSR[ 98 ][ 64 ],
   alphaCSR[ 98 ][ 65 ],
   alphaCSR[ 98 ][ 66 ],
   alphaCSR[ 98 ][ 67 ],
   alphaCSR[ 98 ][ 68 ],
   alphaCSR[ 98 ][ 69 ],
   alphaCSR[ 98 ][ 70 ],
   alphaCSR[ 98 ][ 71 ],
   alphaCSR[ 98 ][ 72 ],
   alphaCSR[ 98 ][ 73 ],
   alphaCSR[ 98 ][ 74 ],
   alphaCSR[ 98 ][ 75 ],
   alphaCSR[ 98 ][ 76 ],
   alphaCSR[ 98 ][ 77 ],
   alphaCSR[ 98 ][ 78 ],
   alphaCSR[ 98 ][ 79 ],
   alphaCSR[ 98 ][ 80 ],
   alphaCSR[ 98 ][ 81 ],
   alphaCSR[ 98 ][ 82 ],
   alphaCSR[ 98 ][ 83 ],
   alphaCSR[ 98 ][ 84 ],
   alphaCSR[ 98 ][ 85 ],
   alphaCSR[ 98 ][ 86 ],
   alphaCSR[ 98 ][ 87 ],
   alphaCSR[ 98 ][ 88 ],
   alphaCSR[ 98 ][ 89 ],
   alphaCSR[ 98 ][ 90 ],
   alphaCSR[ 98 ][ 91 ],
   alphaCSR[ 98 ][ 92 ],
   alphaCSR[ 98 ][ 93 ],
   alphaCSR[ 98 ][ 94 ],
   alphaCSR[ 98 ][ 95 ],
   alphaCSR[ 98 ][ 96 ],
   alphaCSR[ 98 ][ 97 ],
   alphaCSR[ 98 ][ 98 ],
   alphaCSR[ 98 ][ 99 ],
   alphaCSR[ 98 ][ 100 ],
   alphaCSR[ 98 ][ 101 ],
   alphaCSR[ 98 ][ 102 ],
   alphaCSR[ 98 ][ 103 ],
   alphaCSR[ 98 ][ 104 ],
   alphaCSR[ 98 ][ 105 ],
   alphaCSR[ 98 ][ 106 ],
   alphaCSR[ 98 ][ 107 ],
   alphaCSR[ 98 ][ 108 ],
   alphaCSR[ 98 ][ 109 ],
   alphaCSR[ 98 ][ 110 ],
   alphaCSR[ 98 ][ 111 ],
   alphaCSR[ 98 ][ 112 ],
   alphaCSR[ 98 ][ 113 ],
   alphaCSR[ 98 ][ 114 ],
   alphaCSR[ 98 ][ 115 ],
   alphaCSR[ 98 ][ 116 ],
   alphaCSR[ 98 ][ 117 ],
   alphaCSR[ 98 ][ 118 ],
   alphaCSR[ 98 ][ 119 ],
   alphaCSR[ 98 ][ 120 ],
   alphaCSR[ 98 ][ 121 ],
   alphaCSR[ 98 ][ 122 ],
   alphaCSR[ 98 ][ 123 ],
   alphaCSR[ 98 ][ 124 ],
   alphaCSR[ 98 ][ 125 ],
   alphaCSR[ 98 ][ 126 ],
   alphaCSR[ 98 ][ 127 ],
   alphaCSR[ 98 ][ 128 ],
   alphaCSR[ 98 ][ 129 ],
   alphaCSR[ 98 ][ 130 ],
   alphaCSR[ 98 ][ 131 ],
   alphaCSR[ 98 ][ 132 ],
   alphaCSR[ 98 ][ 133 ],
   alphaCSR[ 98 ][ 134 ],
   alphaCSR[ 98 ][ 135 ],
   alphaCSR[ 98 ][ 136 ],
   alphaCSR[ 98 ][ 137 ],
   alphaCSR[ 98 ][ 138 ],
   alphaCSR[ 98 ][ 139 ],
   alphaCSR[ 98 ][ 140 ],
   alphaCSR[ 98 ][ 141 ],
   alphaCSR[ 98 ][ 142 ],
   alphaCSR[ 98 ][ 143 ],
   alphaCSR[ 98 ][ 144 ],
   alphaCSR[ 98 ][ 145 ],
   alphaCSR[ 98 ][ 146 ],
   alphaCSR[ 98 ][ 147 ],
   alphaCSR[ 98 ][ 148 ],
   alphaCSR[ 98 ][ 149 ],
   alphaCSR[ 98 ][ 150 ],
   alphaCSR[ 98 ][ 151 ],
   alphaCSR[ 98 ][ 152 ],
   alphaCSR[ 98 ][ 153 ],
   alphaCSR[ 98 ][ 154 ],
   alphaCSR[ 98 ][ 155 ],
   alphaCSR[ 98 ][ 156 ],
   alphaCSR[ 98 ][ 157 ],
   alphaCSR[ 98 ][ 158 ],
   alphaCSR[ 98 ][ 159 ],
   alphaCSR[ 98 ][ 160 ],
   alphaCSR[ 98 ][ 161 ],
   alphaCSR[ 98 ][ 162 ],
   alphaCSR[ 98 ][ 163 ],
   alphaCSR[ 98 ][ 164 ],
   alphaCSR[ 98 ][ 165 ],
   alphaCSR[ 98 ][ 166 ],
   alphaCSR[ 98 ][ 167 ],
   alphaCSR[ 98 ][ 168 ],
   alphaCSR[ 98 ][ 169 ],
   alphaCSR[ 98 ][ 170 ],
   alphaCSR[ 98 ][ 171 ],
   alphaCSR[ 98 ][ 172 ],
   alphaCSR[ 98 ][ 173 ],
   alphaCSR[ 98 ][ 174 ],
   alphaCSR[ 98 ][ 175 ],
   alphaCSR[ 98 ][ 176 ],
   alphaCSR[ 98 ][ 177 ],
   alphaCSR[ 98 ][ 178 ],
   alphaCSR[ 98 ][ 179 ],
   alphaCSR[ 98 ][ 180 ],
   alphaCSR[ 98 ][ 181 ],
   alphaCSR[ 98 ][ 182 ],
   alphaCSR[ 98 ][ 183 ],
   alphaCSR[ 98 ][ 184 ],
   alphaCSR[ 98 ][ 185 ],
   alphaCSR[ 98 ][ 186 ],
   alphaCSR[ 98 ][ 187 ],
   alphaCSR[ 98 ][ 188 ],
   alphaCSR[ 98 ][ 189 ],
   alphaCSR[ 98 ][ 190 ],
   alphaCSR[ 98 ][ 191 ],
   alphaCSR[ 98 ][ 192 ],
   alphaCSR[ 98 ][ 193 ],
   alphaCSR[ 98 ][ 194 ],
   alphaCSR[ 98 ][ 195 ],
   alphaCSR[ 98 ][ 196 ],
   alphaCSR[ 98 ][ 197 ],
   alphaCSR[ 98 ][ 198 ],
   alphaCSR[ 98 ][ 199 ],
   alphaCSR[ 98 ][ 200 ],
   alphaCSR[ 98 ][ 201 ],
   alphaCSR[ 98 ][ 202 ],
   alphaCSR[ 98 ][ 203 ],
   alphaCSR[ 98 ][ 204 ],
   alphaCSR[ 98 ][ 205 ],
   alphaCSR[ 98 ][ 206 ],
   alphaCSR[ 98 ][ 207 ],
   alphaCSR[ 98 ][ 208 ],
   alphaCSR[ 98 ][ 209 ],
   alphaCSR[ 98 ][ 210 ],
   alphaCSR[ 98 ][ 211 ],
   alphaCSR[ 98 ][ 212 ],
   alphaCSR[ 98 ][ 213 ],
   alphaCSR[ 98 ][ 214 ],
   alphaCSR[ 98 ][ 215 ],
   alphaCSR[ 98 ][ 216 ],
   alphaCSR[ 98 ][ 217 ],
   alphaCSR[ 98 ][ 218 ],
   alphaCSR[ 98 ][ 219 ],
   alphaCSR[ 98 ][ 220 ],
   alphaCSR[ 98 ][ 221 ],
   alphaCSR[ 98 ][ 222 ],
   alphaCSR[ 98 ][ 223 ],
   alphaCSR[ 98 ][ 224 ],
   alphaCSR[ 98 ][ 225 ],
   alphaCSR[ 98 ][ 226 ],
   alphaCSR[ 98 ][ 227 ],
   alphaCSR[ 98 ][ 228 ],
   alphaCSR[ 98 ][ 229 ],
   alphaCSR[ 98 ][ 230 ],
   alphaCSR[ 98 ][ 231 ],
   alphaCSR[ 98 ][ 232 ],
   alphaCSR[ 98 ][ 233 ],
   alphaCSR[ 98 ][ 234 ],
   alphaCSR[ 98 ][ 235 ],
   alphaCSR[ 98 ][ 236 ],
   alphaCSR[ 98 ][ 237 ],
   alphaCSR[ 98 ][ 238 ],
   alphaCSR[ 98 ][ 239 ],
   alphaCSR[ 98 ][ 240 ],
   alphaCSR[ 98 ][ 241 ],
   alphaCSR[ 98 ][ 242 ],
   alphaCSR[ 98 ][ 243 ],
   alphaCSR[ 98 ][ 244 ],
   alphaCSR[ 98 ][ 245 ],
   alphaCSR[ 98 ][ 246 ],
   alphaCSR[ 98 ][ 247 ],
   alphaCSR[ 98 ][ 248 ],
   alphaCSR[ 98 ][ 249 ],
   alphaCSR[ 98 ][ 250 ],
   alphaCSR[ 98 ][ 251 ],
   alphaCSR[ 98 ][ 252 ],
   alphaCSR[ 98 ][ 253 ],
   alphaCSR[ 98 ][ 254 ],
   alphaCSR[ 98 ][ 255 ],
   alphaCSR[ 98 ][ 256 ],
   alphaCSR[ 98 ][ 257 ],
   alphaCSR[ 98 ][ 258 ],
   alphaCSR[ 98 ][ 259 ],
   alphaCSR[ 98 ][ 260 ],
   alphaCSR[ 98 ][ 261 ],
   alphaCSR[ 98 ][ 262 ],
   alphaCSR[ 98 ][ 263 ],
   alphaCSR[ 98 ][ 264 ],
   alphaCSR[ 98 ][ 265 ],
   alphaCSR[ 98 ][ 266 ],
   alphaCSR[ 98 ][ 267 ],
   alphaCSR[ 98 ][ 268 ],
   alphaCSR[ 98 ][ 269 ],
   alphaCSR[ 98 ][ 270 ],
   alphaCSR[ 98 ][ 271 ],
   alphaCSR[ 98 ][ 272 ],
   alphaCSR[ 98 ][ 273 ],
   alphaCSR[ 98 ][ 274 ],
   alphaCSR[ 98 ][ 275 ],
   alphaCSR[ 98 ][ 276 ],
   alphaCSR[ 98 ][ 277 ],
   alphaCSR[ 98 ][ 278 ],
   alphaCSR[ 98 ][ 279 ],
   alphaCSR[ 98 ][ 280 ],
   alphaCSR[ 98 ][ 281 ],
   alphaCSR[ 98 ][ 282 ],
   alphaCSR[ 98 ][ 283 ],
   alphaCSR[ 98 ][ 284 ],
   alphaCSR[ 98 ][ 285 ],
   alphaCSR[ 98 ][ 286 ],
   alphaCSR[ 98 ][ 287 ],
   alphaCSR[ 98 ][ 288 ],
   alphaCSR[ 98 ][ 289 ],
   alphaCSR[ 98 ][ 290 ],
   alphaCSR[ 98 ][ 291 ],
   alphaCSR[ 98 ][ 292 ],
   alphaCSR[ 98 ][ 293 ],
   alphaCSR[ 98 ][ 294 ],
   alphaCSR[ 98 ][ 295 ],
   alphaCSR[ 98 ][ 296 ],
   alphaCSR[ 98 ][ 297 ],
   alphaCSR[ 98 ][ 298 ],
   alphaCSR[ 98 ][ 299 ],
   alphaCSR[ 98 ][ 300 ],
   alphaCSR[ 98 ][ 301 ],
   alphaCSR[ 98 ][ 302 ],
   alphaCSR[ 98 ][ 303 ],
   alphaCSR[ 98 ][ 304 ],
   alphaCSR[ 98 ][ 305 ],
   alphaCSR[ 98 ][ 306 ],
   alphaCSR[ 98 ][ 307 ],
   alphaCSR[ 98 ][ 308 ],
   alphaCSR[ 98 ][ 309 ],
   alphaCSR[ 98 ][ 310 ],
   alphaCSR[ 98 ][ 311 ],
   alphaCSR[ 98 ][ 312 ],
   alphaCSR[ 98 ][ 313 ],
   alphaCSR[ 98 ][ 314 ],
   alphaCSR[ 98 ][ 315 ],
   alphaCSR[ 98 ][ 316 ],
   alphaCSR[ 98 ][ 317 ],
   alphaCSR[ 98 ][ 318 ],
   alphaCSR[ 98 ][ 319 ],
   alphaCSR[ 98 ][ 320 ],
   alphaCSR[ 98 ][ 321 ],
   alphaCSR[ 98 ][ 322 ],
   alphaCSR[ 98 ][ 323 ],
   alphaCSR[ 98 ][ 324 ],
   alphaCSR[ 98 ][ 325 ],
   alphaCSR[ 98 ][ 326 ],
   alphaCSR[ 98 ][ 327 ],
   alphaCSR[ 98 ][ 328 ],
   alphaCSR[ 98 ][ 329 ],
   alphaCSR[ 98 ][ 330 ],
   alphaCSR[ 98 ][ 331 ],
   alphaCSR[ 98 ][ 332 ],
   alphaCSR[ 98 ][ 333 ],
   alphaCSR[ 98 ][ 334 ],
   alphaCSR[ 98 ][ 335 ],
   alphaCSR[ 98 ][ 336 ],
   alphaCSR[ 98 ][ 337 ],
   alphaCSR[ 98 ][ 338 ],
   alphaCSR[ 98 ][ 339 ],
   alphaCSR[ 98 ][ 340 ],
   alphaCSR[ 98 ][ 341 ],
   alphaCSR[ 98 ][ 342 ],
   alphaCSR[ 98 ][ 343 ],
   alphaCSR[ 98 ][ 344 ],
   alphaCSR[ 98 ][ 345 ],
   alphaCSR[ 98 ][ 346 ],
   alphaCSR[ 98 ][ 347 ],
   alphaCSR[ 98 ][ 348 ],
   alphaCSR[ 98 ][ 349 ],
   alphaCSR[ 98 ][ 350 ],
   alphaCSR[ 98 ][ 351 ],
   alphaCSR[ 98 ][ 352 ],
   alphaCSR[ 98 ][ 353 ],
   alphaCSR[ 98 ][ 354 ],
   alphaCSR[ 98 ][ 355 ],
   alphaCSR[ 98 ][ 356 ],
   alphaCSR[ 98 ][ 357 ],
   alphaCSR[ 98 ][ 358 ],
   alphaCSR[ 98 ][ 359 ],
   alphaCSR[ 98 ][ 360 ],
   alphaCSR[ 98 ][ 361 ],
   alphaCSR[ 98 ][ 362 ],
   alphaCSR[ 98 ][ 363 ],
   alphaCSR[ 98 ][ 364 ],
   alphaCSR[ 98 ][ 365 ],
   alphaCSR[ 98 ][ 366 ],
   alphaCSR[ 98 ][ 367 ],
   alphaCSR[ 98 ][ 368 ],
   alphaCSR[ 98 ][ 369 ],
   alphaCSR[ 98 ][ 370 ],
   alphaCSR[ 98 ][ 371 ],
   alphaCSR[ 98 ][ 372 ],
   alphaCSR[ 98 ][ 373 ],
   alphaCSR[ 98 ][ 374 ],
   alphaCSR[ 98 ][ 375 ],
   alphaCSR[ 98 ][ 376 ],
   alphaCSR[ 98 ][ 377 ],
   alphaCSR[ 98 ][ 378 ],
   alphaCSR[ 98 ][ 379 ],
   alphaCSR[ 98 ][ 380 ],
   alphaCSR[ 98 ][ 381 ],
   alphaCSR[ 98 ][ 382 ],
   alphaCSR[ 98 ][ 383 ],
   alphaCSR[ 99 ][ 0 ],
   alphaCSR[ 99 ][ 1 ],
   alphaCSR[ 99 ][ 2 ],
   alphaCSR[ 99 ][ 3 ],
   alphaCSR[ 99 ][ 4 ],
   alphaCSR[ 99 ][ 5 ],
   alphaCSR[ 99 ][ 6 ],
   alphaCSR[ 99 ][ 7 ],
   alphaCSR[ 99 ][ 8 ],
   alphaCSR[ 99 ][ 9 ],
   alphaCSR[ 99 ][ 10 ],
   alphaCSR[ 99 ][ 11 ],
   alphaCSR[ 99 ][ 12 ],
   alphaCSR[ 99 ][ 13 ],
   alphaCSR[ 99 ][ 14 ],
   alphaCSR[ 99 ][ 15 ],
   alphaCSR[ 99 ][ 16 ],
   alphaCSR[ 99 ][ 17 ],
   alphaCSR[ 99 ][ 18 ],
   alphaCSR[ 99 ][ 19 ],
   alphaCSR[ 99 ][ 20 ],
   alphaCSR[ 99 ][ 21 ],
   alphaCSR[ 99 ][ 22 ],
   alphaCSR[ 99 ][ 23 ],
   alphaCSR[ 99 ][ 24 ],
   alphaCSR[ 99 ][ 25 ],
   alphaCSR[ 99 ][ 26 ],
   alphaCSR[ 99 ][ 27 ],
   alphaCSR[ 99 ][ 28 ],
   alphaCSR[ 99 ][ 29 ],
   alphaCSR[ 99 ][ 30 ],
   alphaCSR[ 99 ][ 31 ],
   alphaCSR[ 99 ][ 32 ],
   alphaCSR[ 99 ][ 33 ],
   alphaCSR[ 99 ][ 34 ],
   alphaCSR[ 99 ][ 35 ],
   alphaCSR[ 99 ][ 36 ],
   alphaCSR[ 99 ][ 37 ],
   alphaCSR[ 99 ][ 38 ],
   alphaCSR[ 99 ][ 39 ],
   alphaCSR[ 99 ][ 40 ],
   alphaCSR[ 99 ][ 41 ],
   alphaCSR[ 99 ][ 42 ],
   alphaCSR[ 99 ][ 43 ],
   alphaCSR[ 99 ][ 44 ],
   alphaCSR[ 99 ][ 45 ],
   alphaCSR[ 99 ][ 46 ],
   alphaCSR[ 99 ][ 47 ],
   alphaCSR[ 99 ][ 48 ],
   alphaCSR[ 99 ][ 49 ],
   alphaCSR[ 99 ][ 50 ],
   alphaCSR[ 99 ][ 51 ],
   alphaCSR[ 99 ][ 52 ],
   alphaCSR[ 99 ][ 53 ],
   alphaCSR[ 99 ][ 54 ],
   alphaCSR[ 99 ][ 55 ],
   alphaCSR[ 99 ][ 56 ],
   alphaCSR[ 99 ][ 57 ],
   alphaCSR[ 99 ][ 58 ],
   alphaCSR[ 99 ][ 59 ],
   alphaCSR[ 99 ][ 60 ],
   alphaCSR[ 99 ][ 61 ],
   alphaCSR[ 99 ][ 62 ],
   alphaCSR[ 99 ][ 63 ],
   alphaCSR[ 99 ][ 64 ],
   alphaCSR[ 99 ][ 65 ],
   alphaCSR[ 99 ][ 66 ],
   alphaCSR[ 99 ][ 67 ],
   alphaCSR[ 99 ][ 68 ],
   alphaCSR[ 99 ][ 69 ],
   alphaCSR[ 99 ][ 70 ],
   alphaCSR[ 99 ][ 71 ],
   alphaCSR[ 99 ][ 72 ],
   alphaCSR[ 99 ][ 73 ],
   alphaCSR[ 99 ][ 74 ],
   alphaCSR[ 99 ][ 75 ],
   alphaCSR[ 99 ][ 76 ],
   alphaCSR[ 99 ][ 77 ],
   alphaCSR[ 99 ][ 78 ],
   alphaCSR[ 99 ][ 79 ],
   alphaCSR[ 99 ][ 80 ],
   alphaCSR[ 99 ][ 81 ],
   alphaCSR[ 99 ][ 82 ],
   alphaCSR[ 99 ][ 83 ],
   alphaCSR[ 99 ][ 84 ],
   alphaCSR[ 99 ][ 85 ],
   alphaCSR[ 99 ][ 86 ],
   alphaCSR[ 99 ][ 87 ],
   alphaCSR[ 99 ][ 88 ],
   alphaCSR[ 99 ][ 89 ],
   alphaCSR[ 99 ][ 90 ],
   alphaCSR[ 99 ][ 91 ],
   alphaCSR[ 99 ][ 92 ],
   alphaCSR[ 99 ][ 93 ],
   alphaCSR[ 99 ][ 94 ],
   alphaCSR[ 99 ][ 95 ],
   alphaCSR[ 99 ][ 96 ],
   alphaCSR[ 99 ][ 97 ],
   alphaCSR[ 99 ][ 98 ],
   alphaCSR[ 99 ][ 99 ],
   alphaCSR[ 99 ][ 100 ],
   alphaCSR[ 99 ][ 101 ],
   alphaCSR[ 99 ][ 102 ],
   alphaCSR[ 99 ][ 103 ],
   alphaCSR[ 99 ][ 104 ],
   alphaCSR[ 99 ][ 105 ],
   alphaCSR[ 99 ][ 106 ],
   alphaCSR[ 99 ][ 107 ],
   alphaCSR[ 99 ][ 108 ],
   alphaCSR[ 99 ][ 109 ],
   alphaCSR[ 99 ][ 110 ],
   alphaCSR[ 99 ][ 111 ],
   alphaCSR[ 99 ][ 112 ],
   alphaCSR[ 99 ][ 113 ],
   alphaCSR[ 99 ][ 114 ],
   alphaCSR[ 99 ][ 115 ],
   alphaCSR[ 99 ][ 116 ],
   alphaCSR[ 99 ][ 117 ],
   alphaCSR[ 99 ][ 118 ],
   alphaCSR[ 99 ][ 119 ],
   alphaCSR[ 99 ][ 120 ],
   alphaCSR[ 99 ][ 121 ],
   alphaCSR[ 99 ][ 122 ],
   alphaCSR[ 99 ][ 123 ],
   alphaCSR[ 99 ][ 124 ],
   alphaCSR[ 99 ][ 125 ],
   alphaCSR[ 99 ][ 126 ],
   alphaCSR[ 99 ][ 127 ],
   alphaCSR[ 99 ][ 128 ],
   alphaCSR[ 99 ][ 129 ],
   alphaCSR[ 99 ][ 130 ],
   alphaCSR[ 99 ][ 131 ],
   alphaCSR[ 99 ][ 132 ],
   alphaCSR[ 99 ][ 133 ],
   alphaCSR[ 99 ][ 134 ],
   alphaCSR[ 99 ][ 135 ],
   alphaCSR[ 99 ][ 136 ],
   alphaCSR[ 99 ][ 137 ],
   alphaCSR[ 99 ][ 138 ],
   alphaCSR[ 99 ][ 139 ],
   alphaCSR[ 99 ][ 140 ],
   alphaCSR[ 99 ][ 141 ],
   alphaCSR[ 99 ][ 142 ],
   alphaCSR[ 99 ][ 143 ],
   alphaCSR[ 99 ][ 144 ],
   alphaCSR[ 99 ][ 145 ],
   alphaCSR[ 99 ][ 146 ],
   alphaCSR[ 99 ][ 147 ],
   alphaCSR[ 99 ][ 148 ],
   alphaCSR[ 99 ][ 149 ],
   alphaCSR[ 99 ][ 150 ],
   alphaCSR[ 99 ][ 151 ],
   alphaCSR[ 99 ][ 152 ],
   alphaCSR[ 99 ][ 153 ],
   alphaCSR[ 99 ][ 154 ],
   alphaCSR[ 99 ][ 155 ],
   alphaCSR[ 99 ][ 156 ],
   alphaCSR[ 99 ][ 157 ],
   alphaCSR[ 99 ][ 158 ],
   alphaCSR[ 99 ][ 159 ],
   alphaCSR[ 99 ][ 160 ],
   alphaCSR[ 99 ][ 161 ],
   alphaCSR[ 99 ][ 162 ],
   alphaCSR[ 99 ][ 163 ],
   alphaCSR[ 99 ][ 164 ],
   alphaCSR[ 99 ][ 165 ],
   alphaCSR[ 99 ][ 166 ],
   alphaCSR[ 99 ][ 167 ],
   alphaCSR[ 99 ][ 168 ],
   alphaCSR[ 99 ][ 169 ],
   alphaCSR[ 99 ][ 170 ],
   alphaCSR[ 99 ][ 171 ],
   alphaCSR[ 99 ][ 172 ],
   alphaCSR[ 99 ][ 173 ],
   alphaCSR[ 99 ][ 174 ],
   alphaCSR[ 99 ][ 175 ],
   alphaCSR[ 99 ][ 176 ],
   alphaCSR[ 99 ][ 177 ],
   alphaCSR[ 99 ][ 178 ],
   alphaCSR[ 99 ][ 179 ],
   alphaCSR[ 99 ][ 180 ],
   alphaCSR[ 99 ][ 181 ],
   alphaCSR[ 99 ][ 182 ],
   alphaCSR[ 99 ][ 183 ],
   alphaCSR[ 99 ][ 184 ],
   alphaCSR[ 99 ][ 185 ],
   alphaCSR[ 99 ][ 186 ],
   alphaCSR[ 99 ][ 187 ],
   alphaCSR[ 99 ][ 188 ],
   alphaCSR[ 99 ][ 189 ],
   alphaCSR[ 99 ][ 190 ],
   alphaCSR[ 99 ][ 191 ],
   alphaCSR[ 99 ][ 192 ],
   alphaCSR[ 99 ][ 193 ],
   alphaCSR[ 99 ][ 194 ],
   alphaCSR[ 99 ][ 195 ],
   alphaCSR[ 99 ][ 196 ],
   alphaCSR[ 99 ][ 197 ],
   alphaCSR[ 99 ][ 198 ],
   alphaCSR[ 99 ][ 199 ],
   alphaCSR[ 99 ][ 200 ],
   alphaCSR[ 99 ][ 201 ],
   alphaCSR[ 99 ][ 202 ],
   alphaCSR[ 99 ][ 203 ],
   alphaCSR[ 99 ][ 204 ],
   alphaCSR[ 99 ][ 205 ],
   alphaCSR[ 99 ][ 206 ],
   alphaCSR[ 99 ][ 207 ],
   alphaCSR[ 99 ][ 208 ],
   alphaCSR[ 99 ][ 209 ],
   alphaCSR[ 99 ][ 210 ],
   alphaCSR[ 99 ][ 211 ],
   alphaCSR[ 99 ][ 212 ],
   alphaCSR[ 99 ][ 213 ],
   alphaCSR[ 99 ][ 214 ],
   alphaCSR[ 99 ][ 215 ],
   alphaCSR[ 99 ][ 216 ],
   alphaCSR[ 99 ][ 217 ],
   alphaCSR[ 99 ][ 218 ],
   alphaCSR[ 99 ][ 219 ],
   alphaCSR[ 99 ][ 220 ],
   alphaCSR[ 99 ][ 221 ],
   alphaCSR[ 99 ][ 222 ],
   alphaCSR[ 99 ][ 223 ],
   alphaCSR[ 99 ][ 224 ],
   alphaCSR[ 99 ][ 225 ],
   alphaCSR[ 99 ][ 226 ],
   alphaCSR[ 99 ][ 227 ],
   alphaCSR[ 99 ][ 228 ],
   alphaCSR[ 99 ][ 229 ],
   alphaCSR[ 99 ][ 230 ],
   alphaCSR[ 99 ][ 231 ],
   alphaCSR[ 99 ][ 232 ],
   alphaCSR[ 99 ][ 233 ],
   alphaCSR[ 99 ][ 234 ],
   alphaCSR[ 99 ][ 235 ],
   alphaCSR[ 99 ][ 236 ],
   alphaCSR[ 99 ][ 237 ],
   alphaCSR[ 99 ][ 238 ],
   alphaCSR[ 99 ][ 239 ],
   alphaCSR[ 99 ][ 240 ],
   alphaCSR[ 99 ][ 241 ],
   alphaCSR[ 99 ][ 242 ],
   alphaCSR[ 99 ][ 243 ],
   alphaCSR[ 99 ][ 244 ],
   alphaCSR[ 99 ][ 245 ],
   alphaCSR[ 99 ][ 246 ],
   alphaCSR[ 99 ][ 247 ],
   alphaCSR[ 99 ][ 248 ],
   alphaCSR[ 99 ][ 249 ],
   alphaCSR[ 99 ][ 250 ],
   alphaCSR[ 99 ][ 251 ],
   alphaCSR[ 99 ][ 252 ],
   alphaCSR[ 99 ][ 253 ],
   alphaCSR[ 99 ][ 254 ],
   alphaCSR[ 99 ][ 255 ],
   alphaCSR[ 99 ][ 256 ],
   alphaCSR[ 99 ][ 257 ],
   alphaCSR[ 99 ][ 258 ],
   alphaCSR[ 99 ][ 259 ],
   alphaCSR[ 99 ][ 260 ],
   alphaCSR[ 99 ][ 261 ],
   alphaCSR[ 99 ][ 262 ],
   alphaCSR[ 99 ][ 263 ],
   alphaCSR[ 99 ][ 264 ],
   alphaCSR[ 99 ][ 265 ],
   alphaCSR[ 99 ][ 266 ],
   alphaCSR[ 99 ][ 267 ],
   alphaCSR[ 99 ][ 268 ],
   alphaCSR[ 99 ][ 269 ],
   alphaCSR[ 99 ][ 270 ],
   alphaCSR[ 99 ][ 271 ],
   alphaCSR[ 99 ][ 272 ],
   alphaCSR[ 99 ][ 273 ],
   alphaCSR[ 99 ][ 274 ],
   alphaCSR[ 99 ][ 275 ],
   alphaCSR[ 99 ][ 276 ],
   alphaCSR[ 99 ][ 277 ],
   alphaCSR[ 99 ][ 278 ],
   alphaCSR[ 99 ][ 279 ],
   alphaCSR[ 99 ][ 280 ],
   alphaCSR[ 99 ][ 281 ],
   alphaCSR[ 99 ][ 282 ],
   alphaCSR[ 99 ][ 283 ],
   alphaCSR[ 99 ][ 284 ],
   alphaCSR[ 99 ][ 285 ],
   alphaCSR[ 99 ][ 286 ],
   alphaCSR[ 99 ][ 287 ],
   alphaCSR[ 99 ][ 288 ],
   alphaCSR[ 99 ][ 289 ],
   alphaCSR[ 99 ][ 290 ],
   alphaCSR[ 99 ][ 291 ],
   alphaCSR[ 99 ][ 292 ],
   alphaCSR[ 99 ][ 293 ],
   alphaCSR[ 99 ][ 294 ],
   alphaCSR[ 99 ][ 295 ],
   alphaCSR[ 99 ][ 296 ],
   alphaCSR[ 99 ][ 297 ],
   alphaCSR[ 99 ][ 298 ],
   alphaCSR[ 99 ][ 299 ],
   alphaCSR[ 99 ][ 300 ],
   alphaCSR[ 99 ][ 301 ],
   alphaCSR[ 99 ][ 302 ],
   alphaCSR[ 99 ][ 303 ],
   alphaCSR[ 99 ][ 304 ],
   alphaCSR[ 99 ][ 305 ],
   alphaCSR[ 99 ][ 306 ],
   alphaCSR[ 99 ][ 307 ],
   alphaCSR[ 99 ][ 308 ],
   alphaCSR[ 99 ][ 309 ],
   alphaCSR[ 99 ][ 310 ],
   alphaCSR[ 99 ][ 311 ],
   alphaCSR[ 99 ][ 312 ],
   alphaCSR[ 99 ][ 313 ],
   alphaCSR[ 99 ][ 314 ],
   alphaCSR[ 99 ][ 315 ],
   alphaCSR[ 99 ][ 316 ],
   alphaCSR[ 99 ][ 317 ],
   alphaCSR[ 99 ][ 318 ],
   alphaCSR[ 99 ][ 319 ],
   alphaCSR[ 99 ][ 320 ],
   alphaCSR[ 99 ][ 321 ],
   alphaCSR[ 99 ][ 322 ],
   alphaCSR[ 99 ][ 323 ],
   alphaCSR[ 99 ][ 324 ],
   alphaCSR[ 99 ][ 325 ],
   alphaCSR[ 99 ][ 326 ],
   alphaCSR[ 99 ][ 327 ],
   alphaCSR[ 99 ][ 328 ],
   alphaCSR[ 99 ][ 329 ],
   alphaCSR[ 99 ][ 330 ],
   alphaCSR[ 99 ][ 331 ],
   alphaCSR[ 99 ][ 332 ],
   alphaCSR[ 99 ][ 333 ],
   alphaCSR[ 99 ][ 334 ],
   alphaCSR[ 99 ][ 335 ],
   alphaCSR[ 99 ][ 336 ],
   alphaCSR[ 99 ][ 337 ],
   alphaCSR[ 99 ][ 338 ],
   alphaCSR[ 99 ][ 339 ],
   alphaCSR[ 99 ][ 340 ],
   alphaCSR[ 99 ][ 341 ],
   alphaCSR[ 99 ][ 342 ],
   alphaCSR[ 99 ][ 343 ],
   alphaCSR[ 99 ][ 344 ],
   alphaCSR[ 99 ][ 345 ],
   alphaCSR[ 99 ][ 346 ],
   alphaCSR[ 99 ][ 347 ],
   alphaCSR[ 99 ][ 348 ],
   alphaCSR[ 99 ][ 349 ],
   alphaCSR[ 99 ][ 350 ],
   alphaCSR[ 99 ][ 351 ],
   alphaCSR[ 99 ][ 352 ],
   alphaCSR[ 99 ][ 353 ],
   alphaCSR[ 99 ][ 354 ],
   alphaCSR[ 99 ][ 355 ],
   alphaCSR[ 99 ][ 356 ],
   alphaCSR[ 99 ][ 357 ],
   alphaCSR[ 99 ][ 358 ],
   alphaCSR[ 99 ][ 359 ],
   alphaCSR[ 99 ][ 360 ],
   alphaCSR[ 99 ][ 361 ],
   alphaCSR[ 99 ][ 362 ],
   alphaCSR[ 99 ][ 363 ],
   alphaCSR[ 99 ][ 364 ],
   alphaCSR[ 99 ][ 365 ],
   alphaCSR[ 99 ][ 366 ],
   alphaCSR[ 99 ][ 367 ],
   alphaCSR[ 99 ][ 368 ],
   alphaCSR[ 99 ][ 369 ],
   alphaCSR[ 99 ][ 370 ],
   alphaCSR[ 99 ][ 371 ],
   alphaCSR[ 99 ][ 372 ],
   alphaCSR[ 99 ][ 373 ],
   alphaCSR[ 99 ][ 374 ],
   alphaCSR[ 99 ][ 375 ],
   alphaCSR[ 99 ][ 376 ],
   alphaCSR[ 99 ][ 377 ],
   alphaCSR[ 99 ][ 378 ],
   alphaCSR[ 99 ][ 379 ],
   alphaCSR[ 99 ][ 380 ],
   alphaCSR[ 99 ][ 381 ],
   alphaCSR[ 99 ][ 382 ],
   alphaCSR[ 99 ][ 383 ],
   alphaCSR[ 100 ][ 0 ],
   alphaCSR[ 100 ][ 1 ],
   alphaCSR[ 100 ][ 2 ],
   alphaCSR[ 100 ][ 3 ],
   alphaCSR[ 100 ][ 4 ],
   alphaCSR[ 100 ][ 5 ],
   alphaCSR[ 100 ][ 6 ],
   alphaCSR[ 100 ][ 7 ],
   alphaCSR[ 100 ][ 8 ],
   alphaCSR[ 100 ][ 9 ],
   alphaCSR[ 100 ][ 10 ],
   alphaCSR[ 100 ][ 11 ],
   alphaCSR[ 100 ][ 12 ],
   alphaCSR[ 100 ][ 13 ],
   alphaCSR[ 100 ][ 14 ],
   alphaCSR[ 100 ][ 15 ],
   alphaCSR[ 100 ][ 16 ],
   alphaCSR[ 100 ][ 17 ],
   alphaCSR[ 100 ][ 18 ],
   alphaCSR[ 100 ][ 19 ],
   alphaCSR[ 100 ][ 20 ],
   alphaCSR[ 100 ][ 21 ],
   alphaCSR[ 100 ][ 22 ],
   alphaCSR[ 100 ][ 23 ],
   alphaCSR[ 100 ][ 24 ],
   alphaCSR[ 100 ][ 25 ],
   alphaCSR[ 100 ][ 26 ],
   alphaCSR[ 100 ][ 27 ],
   alphaCSR[ 100 ][ 28 ],
   alphaCSR[ 100 ][ 29 ],
   alphaCSR[ 100 ][ 30 ],
   alphaCSR[ 100 ][ 31 ],
   alphaCSR[ 100 ][ 32 ],
   alphaCSR[ 100 ][ 33 ],
   alphaCSR[ 100 ][ 34 ],
   alphaCSR[ 100 ][ 35 ],
   alphaCSR[ 100 ][ 36 ],
   alphaCSR[ 100 ][ 37 ],
   alphaCSR[ 100 ][ 38 ],
   alphaCSR[ 100 ][ 39 ],
   alphaCSR[ 100 ][ 40 ],
   alphaCSR[ 100 ][ 41 ],
   alphaCSR[ 100 ][ 42 ],
   alphaCSR[ 100 ][ 43 ],
   alphaCSR[ 100 ][ 44 ],
   alphaCSR[ 100 ][ 45 ],
   alphaCSR[ 100 ][ 46 ],
   alphaCSR[ 100 ][ 47 ],
   alphaCSR[ 100 ][ 48 ],
   alphaCSR[ 100 ][ 49 ],
   alphaCSR[ 100 ][ 50 ],
   alphaCSR[ 100 ][ 51 ],
   alphaCSR[ 100 ][ 52 ],
   alphaCSR[ 100 ][ 53 ],
   alphaCSR[ 100 ][ 54 ],
   alphaCSR[ 100 ][ 55 ],
   alphaCSR[ 100 ][ 56 ],
   alphaCSR[ 100 ][ 57 ],
   alphaCSR[ 100 ][ 58 ],
   alphaCSR[ 100 ][ 59 ],
   alphaCSR[ 100 ][ 60 ],
   alphaCSR[ 100 ][ 61 ],
   alphaCSR[ 100 ][ 62 ],
   alphaCSR[ 100 ][ 63 ],
   alphaCSR[ 100 ][ 64 ],
   alphaCSR[ 100 ][ 65 ],
   alphaCSR[ 100 ][ 66 ],
   alphaCSR[ 100 ][ 67 ],
   alphaCSR[ 100 ][ 68 ],
   alphaCSR[ 100 ][ 69 ],
   alphaCSR[ 100 ][ 70 ],
   alphaCSR[ 100 ][ 71 ],
   alphaCSR[ 100 ][ 72 ],
   alphaCSR[ 100 ][ 73 ],
   alphaCSR[ 100 ][ 74 ],
   alphaCSR[ 100 ][ 75 ],
   alphaCSR[ 100 ][ 76 ],
   alphaCSR[ 100 ][ 77 ],
   alphaCSR[ 100 ][ 78 ],
   alphaCSR[ 100 ][ 79 ],
   alphaCSR[ 100 ][ 80 ],
   alphaCSR[ 100 ][ 81 ],
   alphaCSR[ 100 ][ 82 ],
   alphaCSR[ 100 ][ 83 ],
   alphaCSR[ 100 ][ 84 ],
   alphaCSR[ 100 ][ 85 ],
   alphaCSR[ 100 ][ 86 ],
   alphaCSR[ 100 ][ 87 ],
   alphaCSR[ 100 ][ 88 ],
   alphaCSR[ 100 ][ 89 ],
   alphaCSR[ 100 ][ 90 ],
   alphaCSR[ 100 ][ 91 ],
   alphaCSR[ 100 ][ 92 ],
   alphaCSR[ 100 ][ 93 ],
   alphaCSR[ 100 ][ 94 ],
   alphaCSR[ 100 ][ 95 ],
   alphaCSR[ 100 ][ 96 ],
   alphaCSR[ 100 ][ 97 ],
   alphaCSR[ 100 ][ 98 ],
   alphaCSR[ 100 ][ 99 ],
   alphaCSR[ 100 ][ 100 ],
   alphaCSR[ 100 ][ 101 ],
   alphaCSR[ 100 ][ 102 ],
   alphaCSR[ 100 ][ 103 ],
   alphaCSR[ 100 ][ 104 ],
   alphaCSR[ 100 ][ 105 ],
   alphaCSR[ 100 ][ 106 ],
   alphaCSR[ 100 ][ 107 ],
   alphaCSR[ 100 ][ 108 ],
   alphaCSR[ 100 ][ 109 ],
   alphaCSR[ 100 ][ 110 ],
   alphaCSR[ 100 ][ 111 ],
   alphaCSR[ 100 ][ 112 ],
   alphaCSR[ 100 ][ 113 ],
   alphaCSR[ 100 ][ 114 ],
   alphaCSR[ 100 ][ 115 ],
   alphaCSR[ 100 ][ 116 ],
   alphaCSR[ 100 ][ 117 ],
   alphaCSR[ 100 ][ 118 ],
   alphaCSR[ 100 ][ 119 ],
   alphaCSR[ 100 ][ 120 ],
   alphaCSR[ 100 ][ 121 ],
   alphaCSR[ 100 ][ 122 ],
   alphaCSR[ 100 ][ 123 ],
   alphaCSR[ 100 ][ 124 ],
   alphaCSR[ 100 ][ 125 ],
   alphaCSR[ 100 ][ 126 ],
   alphaCSR[ 100 ][ 127 ],
   alphaCSR[ 100 ][ 128 ],
   alphaCSR[ 100 ][ 129 ],
   alphaCSR[ 100 ][ 130 ],
   alphaCSR[ 100 ][ 131 ],
   alphaCSR[ 100 ][ 132 ],
   alphaCSR[ 100 ][ 133 ],
   alphaCSR[ 100 ][ 134 ],
   alphaCSR[ 100 ][ 135 ],
   alphaCSR[ 100 ][ 136 ],
   alphaCSR[ 100 ][ 137 ],
   alphaCSR[ 100 ][ 138 ],
   alphaCSR[ 100 ][ 139 ],
   alphaCSR[ 100 ][ 140 ],
   alphaCSR[ 100 ][ 141 ],
   alphaCSR[ 100 ][ 142 ],
   alphaCSR[ 100 ][ 143 ],
   alphaCSR[ 100 ][ 144 ],
   alphaCSR[ 100 ][ 145 ],
   alphaCSR[ 100 ][ 146 ],
   alphaCSR[ 100 ][ 147 ],
   alphaCSR[ 100 ][ 148 ],
   alphaCSR[ 100 ][ 149 ],
   alphaCSR[ 100 ][ 150 ],
   alphaCSR[ 100 ][ 151 ],
   alphaCSR[ 100 ][ 152 ],
   alphaCSR[ 100 ][ 153 ],
   alphaCSR[ 100 ][ 154 ],
   alphaCSR[ 100 ][ 155 ],
   alphaCSR[ 100 ][ 156 ],
   alphaCSR[ 100 ][ 157 ],
   alphaCSR[ 100 ][ 158 ],
   alphaCSR[ 100 ][ 159 ],
   alphaCSR[ 100 ][ 160 ],
   alphaCSR[ 100 ][ 161 ],
   alphaCSR[ 100 ][ 162 ],
   alphaCSR[ 100 ][ 163 ],
   alphaCSR[ 100 ][ 164 ],
   alphaCSR[ 100 ][ 165 ],
   alphaCSR[ 100 ][ 166 ],
   alphaCSR[ 100 ][ 167 ],
   alphaCSR[ 100 ][ 168 ],
   alphaCSR[ 100 ][ 169 ],
   alphaCSR[ 100 ][ 170 ],
   alphaCSR[ 100 ][ 171 ],
   alphaCSR[ 100 ][ 172 ],
   alphaCSR[ 100 ][ 173 ],
   alphaCSR[ 100 ][ 174 ],
   alphaCSR[ 100 ][ 175 ],
   alphaCSR[ 100 ][ 176 ],
   alphaCSR[ 100 ][ 177 ],
   alphaCSR[ 100 ][ 178 ],
   alphaCSR[ 100 ][ 179 ],
   alphaCSR[ 100 ][ 180 ],
   alphaCSR[ 100 ][ 181 ],
   alphaCSR[ 100 ][ 182 ],
   alphaCSR[ 100 ][ 183 ],
   alphaCSR[ 100 ][ 184 ],
   alphaCSR[ 100 ][ 185 ],
   alphaCSR[ 100 ][ 186 ],
   alphaCSR[ 100 ][ 187 ],
   alphaCSR[ 100 ][ 188 ],
   alphaCSR[ 100 ][ 189 ],
   alphaCSR[ 100 ][ 190 ],
   alphaCSR[ 100 ][ 191 ],
   alphaCSR[ 100 ][ 192 ],
   alphaCSR[ 100 ][ 193 ],
   alphaCSR[ 100 ][ 194 ],
   alphaCSR[ 100 ][ 195 ],
   alphaCSR[ 100 ][ 196 ],
   alphaCSR[ 100 ][ 197 ],
   alphaCSR[ 100 ][ 198 ],
   alphaCSR[ 100 ][ 199 ],
   alphaCSR[ 100 ][ 200 ],
   alphaCSR[ 100 ][ 201 ],
   alphaCSR[ 100 ][ 202 ],
   alphaCSR[ 100 ][ 203 ],
   alphaCSR[ 100 ][ 204 ],
   alphaCSR[ 100 ][ 205 ],
   alphaCSR[ 100 ][ 206 ],
   alphaCSR[ 100 ][ 207 ],
   alphaCSR[ 100 ][ 208 ],
   alphaCSR[ 100 ][ 209 ],
   alphaCSR[ 100 ][ 210 ],
   alphaCSR[ 100 ][ 211 ],
   alphaCSR[ 100 ][ 212 ],
   alphaCSR[ 100 ][ 213 ],
   alphaCSR[ 100 ][ 214 ],
   alphaCSR[ 100 ][ 215 ],
   alphaCSR[ 100 ][ 216 ],
   alphaCSR[ 100 ][ 217 ],
   alphaCSR[ 100 ][ 218 ],
   alphaCSR[ 100 ][ 219 ],
   alphaCSR[ 100 ][ 220 ],
   alphaCSR[ 100 ][ 221 ],
   alphaCSR[ 100 ][ 222 ],
   alphaCSR[ 100 ][ 223 ],
   alphaCSR[ 100 ][ 224 ],
   alphaCSR[ 100 ][ 225 ],
   alphaCSR[ 100 ][ 226 ],
   alphaCSR[ 100 ][ 227 ],
   alphaCSR[ 100 ][ 228 ],
   alphaCSR[ 100 ][ 229 ],
   alphaCSR[ 100 ][ 230 ],
   alphaCSR[ 100 ][ 231 ],
   alphaCSR[ 100 ][ 232 ],
   alphaCSR[ 100 ][ 233 ],
   alphaCSR[ 100 ][ 234 ],
   alphaCSR[ 100 ][ 235 ],
   alphaCSR[ 100 ][ 236 ],
   alphaCSR[ 100 ][ 237 ],
   alphaCSR[ 100 ][ 238 ],
   alphaCSR[ 100 ][ 239 ],
   alphaCSR[ 100 ][ 240 ],
   alphaCSR[ 100 ][ 241 ],
   alphaCSR[ 100 ][ 242 ],
   alphaCSR[ 100 ][ 243 ],
   alphaCSR[ 100 ][ 244 ],
   alphaCSR[ 100 ][ 245 ],
   alphaCSR[ 100 ][ 246 ],
   alphaCSR[ 100 ][ 247 ],
   alphaCSR[ 100 ][ 248 ],
   alphaCSR[ 100 ][ 249 ],
   alphaCSR[ 100 ][ 250 ],
   alphaCSR[ 100 ][ 251 ],
   alphaCSR[ 100 ][ 252 ],
   alphaCSR[ 100 ][ 253 ],
   alphaCSR[ 100 ][ 254 ],
   alphaCSR[ 100 ][ 255 ],
   alphaCSR[ 100 ][ 256 ],
   alphaCSR[ 100 ][ 257 ],
   alphaCSR[ 100 ][ 258 ],
   alphaCSR[ 100 ][ 259 ],
   alphaCSR[ 100 ][ 260 ],
   alphaCSR[ 100 ][ 261 ],
   alphaCSR[ 100 ][ 262 ],
   alphaCSR[ 100 ][ 263 ],
   alphaCSR[ 100 ][ 264 ],
   alphaCSR[ 100 ][ 265 ],
   alphaCSR[ 100 ][ 266 ],
   alphaCSR[ 100 ][ 267 ],
   alphaCSR[ 100 ][ 268 ],
   alphaCSR[ 100 ][ 269 ],
   alphaCSR[ 100 ][ 270 ],
   alphaCSR[ 100 ][ 271 ],
   alphaCSR[ 100 ][ 272 ],
   alphaCSR[ 100 ][ 273 ],
   alphaCSR[ 100 ][ 274 ],
   alphaCSR[ 100 ][ 275 ],
   alphaCSR[ 100 ][ 276 ],
   alphaCSR[ 100 ][ 277 ],
   alphaCSR[ 100 ][ 278 ],
   alphaCSR[ 100 ][ 279 ],
   alphaCSR[ 100 ][ 280 ],
   alphaCSR[ 100 ][ 281 ],
   alphaCSR[ 100 ][ 282 ],
   alphaCSR[ 100 ][ 283 ],
   alphaCSR[ 100 ][ 284 ],
   alphaCSR[ 100 ][ 285 ],
   alphaCSR[ 100 ][ 286 ],
   alphaCSR[ 100 ][ 287 ],
   alphaCSR[ 100 ][ 288 ],
   alphaCSR[ 100 ][ 289 ],
   alphaCSR[ 100 ][ 290 ],
   alphaCSR[ 100 ][ 291 ],
   alphaCSR[ 100 ][ 292 ],
   alphaCSR[ 100 ][ 293 ],
   alphaCSR[ 100 ][ 294 ],
   alphaCSR[ 100 ][ 295 ],
   alphaCSR[ 100 ][ 296 ],
   alphaCSR[ 100 ][ 297 ],
   alphaCSR[ 100 ][ 298 ],
   alphaCSR[ 100 ][ 299 ],
   alphaCSR[ 100 ][ 300 ],
   alphaCSR[ 100 ][ 301 ],
   alphaCSR[ 100 ][ 302 ],
   alphaCSR[ 100 ][ 303 ],
   alphaCSR[ 100 ][ 304 ],
   alphaCSR[ 100 ][ 305 ],
   alphaCSR[ 100 ][ 306 ],
   alphaCSR[ 100 ][ 307 ],
   alphaCSR[ 100 ][ 308 ],
   alphaCSR[ 100 ][ 309 ],
   alphaCSR[ 100 ][ 310 ],
   alphaCSR[ 100 ][ 311 ],
   alphaCSR[ 100 ][ 312 ],
   alphaCSR[ 100 ][ 313 ],
   alphaCSR[ 100 ][ 314 ],
   alphaCSR[ 100 ][ 315 ],
   alphaCSR[ 100 ][ 316 ],
   alphaCSR[ 100 ][ 317 ],
   alphaCSR[ 100 ][ 318 ],
   alphaCSR[ 100 ][ 319 ],
   alphaCSR[ 100 ][ 320 ],
   alphaCSR[ 100 ][ 321 ],
   alphaCSR[ 100 ][ 322 ],
   alphaCSR[ 100 ][ 323 ],
   alphaCSR[ 100 ][ 324 ],
   alphaCSR[ 100 ][ 325 ],
   alphaCSR[ 100 ][ 326 ],
   alphaCSR[ 100 ][ 327 ],
   alphaCSR[ 100 ][ 328 ],
   alphaCSR[ 100 ][ 329 ],
   alphaCSR[ 100 ][ 330 ],
   alphaCSR[ 100 ][ 331 ],
   alphaCSR[ 100 ][ 332 ],
   alphaCSR[ 100 ][ 333 ],
   alphaCSR[ 100 ][ 334 ],
   alphaCSR[ 100 ][ 335 ],
   alphaCSR[ 100 ][ 336 ],
   alphaCSR[ 100 ][ 337 ],
   alphaCSR[ 100 ][ 338 ],
   alphaCSR[ 100 ][ 339 ],
   alphaCSR[ 100 ][ 340 ],
   alphaCSR[ 100 ][ 341 ],
   alphaCSR[ 100 ][ 342 ],
   alphaCSR[ 100 ][ 343 ],
   alphaCSR[ 100 ][ 344 ],
   alphaCSR[ 100 ][ 345 ],
   alphaCSR[ 100 ][ 346 ],
   alphaCSR[ 100 ][ 347 ],
   alphaCSR[ 100 ][ 348 ],
   alphaCSR[ 100 ][ 349 ],
   alphaCSR[ 100 ][ 350 ],
   alphaCSR[ 100 ][ 351 ],
   alphaCSR[ 100 ][ 352 ],
   alphaCSR[ 100 ][ 353 ],
   alphaCSR[ 100 ][ 354 ],
   alphaCSR[ 100 ][ 355 ],
   alphaCSR[ 100 ][ 356 ],
   alphaCSR[ 100 ][ 357 ],
   alphaCSR[ 100 ][ 358 ],
   alphaCSR[ 100 ][ 359 ],
   alphaCSR[ 100 ][ 360 ],
   alphaCSR[ 100 ][ 361 ],
   alphaCSR[ 100 ][ 362 ],
   alphaCSR[ 100 ][ 363 ],
   alphaCSR[ 100 ][ 364 ],
   alphaCSR[ 100 ][ 365 ],
   alphaCSR[ 100 ][ 366 ],
   alphaCSR[ 100 ][ 367 ],
   alphaCSR[ 100 ][ 368 ],
   alphaCSR[ 100 ][ 369 ],
   alphaCSR[ 100 ][ 370 ],
   alphaCSR[ 100 ][ 371 ],
   alphaCSR[ 100 ][ 372 ],
   alphaCSR[ 100 ][ 373 ],
   alphaCSR[ 100 ][ 374 ],
   alphaCSR[ 100 ][ 375 ],
   alphaCSR[ 100 ][ 376 ],
   alphaCSR[ 100 ][ 377 ],
   alphaCSR[ 100 ][ 378 ],
   alphaCSR[ 100 ][ 379 ],
   alphaCSR[ 100 ][ 380 ],
   alphaCSR[ 100 ][ 381 ],
   alphaCSR[ 100 ][ 382 ],
   alphaCSR[ 100 ][ 383 ],
   alphaCSR[ 101 ][ 0 ],
   alphaCSR[ 101 ][ 1 ],
   alphaCSR[ 101 ][ 2 ],
   alphaCSR[ 101 ][ 3 ],
   alphaCSR[ 101 ][ 4 ],
   alphaCSR[ 101 ][ 5 ],
   alphaCSR[ 101 ][ 6 ],
   alphaCSR[ 101 ][ 7 ],
   alphaCSR[ 101 ][ 8 ],
   alphaCSR[ 101 ][ 9 ],
   alphaCSR[ 101 ][ 10 ],
   alphaCSR[ 101 ][ 11 ],
   alphaCSR[ 101 ][ 12 ],
   alphaCSR[ 101 ][ 13 ],
   alphaCSR[ 101 ][ 14 ],
   alphaCSR[ 101 ][ 15 ],
   alphaCSR[ 101 ][ 16 ],
   alphaCSR[ 101 ][ 17 ],
   alphaCSR[ 101 ][ 18 ],
   alphaCSR[ 101 ][ 19 ],
   alphaCSR[ 101 ][ 20 ],
   alphaCSR[ 101 ][ 21 ],
   alphaCSR[ 101 ][ 22 ],
   alphaCSR[ 101 ][ 23 ],
   alphaCSR[ 101 ][ 24 ],
   alphaCSR[ 101 ][ 25 ],
   alphaCSR[ 101 ][ 26 ],
   alphaCSR[ 101 ][ 27 ],
   alphaCSR[ 101 ][ 28 ],
   alphaCSR[ 101 ][ 29 ],
   alphaCSR[ 101 ][ 30 ],
   alphaCSR[ 101 ][ 31 ],
   alphaCSR[ 101 ][ 32 ],
   alphaCSR[ 101 ][ 33 ],
   alphaCSR[ 101 ][ 34 ],
   alphaCSR[ 101 ][ 35 ],
   alphaCSR[ 101 ][ 36 ],
   alphaCSR[ 101 ][ 37 ],
   alphaCSR[ 101 ][ 38 ],
   alphaCSR[ 101 ][ 39 ],
   alphaCSR[ 101 ][ 40 ],
   alphaCSR[ 101 ][ 41 ],
   alphaCSR[ 101 ][ 42 ],
   alphaCSR[ 101 ][ 43 ],
   alphaCSR[ 101 ][ 44 ],
   alphaCSR[ 101 ][ 45 ],
   alphaCSR[ 101 ][ 46 ],
   alphaCSR[ 101 ][ 47 ],
   alphaCSR[ 101 ][ 48 ],
   alphaCSR[ 101 ][ 49 ],
   alphaCSR[ 101 ][ 50 ],
   alphaCSR[ 101 ][ 51 ],
   alphaCSR[ 101 ][ 52 ],
   alphaCSR[ 101 ][ 53 ],
   alphaCSR[ 101 ][ 54 ],
   alphaCSR[ 101 ][ 55 ],
   alphaCSR[ 101 ][ 56 ],
   alphaCSR[ 101 ][ 57 ],
   alphaCSR[ 101 ][ 58 ],
   alphaCSR[ 101 ][ 59 ],
   alphaCSR[ 101 ][ 60 ],
   alphaCSR[ 101 ][ 61 ],
   alphaCSR[ 101 ][ 62 ],
   alphaCSR[ 101 ][ 63 ],
   alphaCSR[ 101 ][ 64 ],
   alphaCSR[ 101 ][ 65 ],
   alphaCSR[ 101 ][ 66 ],
   alphaCSR[ 101 ][ 67 ],
   alphaCSR[ 101 ][ 68 ],
   alphaCSR[ 101 ][ 69 ],
   alphaCSR[ 101 ][ 70 ],
   alphaCSR[ 101 ][ 71 ],
   alphaCSR[ 101 ][ 72 ],
   alphaCSR[ 101 ][ 73 ],
   alphaCSR[ 101 ][ 74 ],
   alphaCSR[ 101 ][ 75 ],
   alphaCSR[ 101 ][ 76 ],
   alphaCSR[ 101 ][ 77 ],
   alphaCSR[ 101 ][ 78 ],
   alphaCSR[ 101 ][ 79 ],
   alphaCSR[ 101 ][ 80 ],
   alphaCSR[ 101 ][ 81 ],
   alphaCSR[ 101 ][ 82 ],
   alphaCSR[ 101 ][ 83 ],
   alphaCSR[ 101 ][ 84 ],
   alphaCSR[ 101 ][ 85 ],
   alphaCSR[ 101 ][ 86 ],
   alphaCSR[ 101 ][ 87 ],
   alphaCSR[ 101 ][ 88 ],
   alphaCSR[ 101 ][ 89 ],
   alphaCSR[ 101 ][ 90 ],
   alphaCSR[ 101 ][ 91 ],
   alphaCSR[ 101 ][ 92 ],
   alphaCSR[ 101 ][ 93 ],
   alphaCSR[ 101 ][ 94 ],
   alphaCSR[ 101 ][ 95 ],
   alphaCSR[ 101 ][ 96 ],
   alphaCSR[ 101 ][ 97 ],
   alphaCSR[ 101 ][ 98 ],
   alphaCSR[ 101 ][ 99 ],
   alphaCSR[ 101 ][ 100 ],
   alphaCSR[ 101 ][ 101 ],
   alphaCSR[ 101 ][ 102 ],
   alphaCSR[ 101 ][ 103 ],
   alphaCSR[ 101 ][ 104 ],
   alphaCSR[ 101 ][ 105 ],
   alphaCSR[ 101 ][ 106 ],
   alphaCSR[ 101 ][ 107 ],
   alphaCSR[ 101 ][ 108 ],
   alphaCSR[ 101 ][ 109 ],
   alphaCSR[ 101 ][ 110 ],
   alphaCSR[ 101 ][ 111 ],
   alphaCSR[ 101 ][ 112 ],
   alphaCSR[ 101 ][ 113 ],
   alphaCSR[ 101 ][ 114 ],
   alphaCSR[ 101 ][ 115 ],
   alphaCSR[ 101 ][ 116 ],
   alphaCSR[ 101 ][ 117 ],
   alphaCSR[ 101 ][ 118 ],
   alphaCSR[ 101 ][ 119 ],
   alphaCSR[ 101 ][ 120 ],
   alphaCSR[ 101 ][ 121 ],
   alphaCSR[ 101 ][ 122 ],
   alphaCSR[ 101 ][ 123 ],
   alphaCSR[ 101 ][ 124 ],
   alphaCSR[ 101 ][ 125 ],
   alphaCSR[ 101 ][ 126 ],
   alphaCSR[ 101 ][ 127 ],
   alphaCSR[ 101 ][ 128 ],
   alphaCSR[ 101 ][ 129 ],
   alphaCSR[ 101 ][ 130 ],
   alphaCSR[ 101 ][ 131 ],
   alphaCSR[ 101 ][ 132 ],
   alphaCSR[ 101 ][ 133 ],
   alphaCSR[ 101 ][ 134 ],
   alphaCSR[ 101 ][ 135 ],
   alphaCSR[ 101 ][ 136 ],
   alphaCSR[ 101 ][ 137 ],
   alphaCSR[ 101 ][ 138 ],
   alphaCSR[ 101 ][ 139 ],
   alphaCSR[ 101 ][ 140 ],
   alphaCSR[ 101 ][ 141 ],
   alphaCSR[ 101 ][ 142 ],
   alphaCSR[ 101 ][ 143 ],
   alphaCSR[ 101 ][ 144 ],
   alphaCSR[ 101 ][ 145 ],
   alphaCSR[ 101 ][ 146 ],
   alphaCSR[ 101 ][ 147 ],
   alphaCSR[ 101 ][ 148 ],
   alphaCSR[ 101 ][ 149 ],
   alphaCSR[ 101 ][ 150 ],
   alphaCSR[ 101 ][ 151 ],
   alphaCSR[ 101 ][ 152 ],
   alphaCSR[ 101 ][ 153 ],
   alphaCSR[ 101 ][ 154 ],
   alphaCSR[ 101 ][ 155 ],
   alphaCSR[ 101 ][ 156 ],
   alphaCSR[ 101 ][ 157 ],
   alphaCSR[ 101 ][ 158 ],
   alphaCSR[ 101 ][ 159 ],
   alphaCSR[ 101 ][ 160 ],
   alphaCSR[ 101 ][ 161 ],
   alphaCSR[ 101 ][ 162 ],
   alphaCSR[ 101 ][ 163 ],
   alphaCSR[ 101 ][ 164 ],
   alphaCSR[ 101 ][ 165 ],
   alphaCSR[ 101 ][ 166 ],
   alphaCSR[ 101 ][ 167 ],
   alphaCSR[ 101 ][ 168 ],
   alphaCSR[ 101 ][ 169 ],
   alphaCSR[ 101 ][ 170 ],
   alphaCSR[ 101 ][ 171 ],
   alphaCSR[ 101 ][ 172 ],
   alphaCSR[ 101 ][ 173 ],
   alphaCSR[ 101 ][ 174 ],
   alphaCSR[ 101 ][ 175 ],
   alphaCSR[ 101 ][ 176 ],
   alphaCSR[ 101 ][ 177 ],
   alphaCSR[ 101 ][ 178 ],
   alphaCSR[ 101 ][ 179 ],
   alphaCSR[ 101 ][ 180 ],
   alphaCSR[ 101 ][ 181 ],
   alphaCSR[ 101 ][ 182 ],
   alphaCSR[ 101 ][ 183 ],
   alphaCSR[ 101 ][ 184 ],
   alphaCSR[ 101 ][ 185 ],
   alphaCSR[ 101 ][ 186 ],
   alphaCSR[ 101 ][ 187 ],
   alphaCSR[ 101 ][ 188 ],
   alphaCSR[ 101 ][ 189 ],
   alphaCSR[ 101 ][ 190 ],
   alphaCSR[ 101 ][ 191 ],
   alphaCSR[ 101 ][ 192 ],
   alphaCSR[ 101 ][ 193 ],
   alphaCSR[ 101 ][ 194 ],
   alphaCSR[ 101 ][ 195 ],
   alphaCSR[ 101 ][ 196 ],
   alphaCSR[ 101 ][ 197 ],
   alphaCSR[ 101 ][ 198 ],
   alphaCSR[ 101 ][ 199 ],
   alphaCSR[ 101 ][ 200 ],
   alphaCSR[ 101 ][ 201 ],
   alphaCSR[ 101 ][ 202 ],
   alphaCSR[ 101 ][ 203 ],
   alphaCSR[ 101 ][ 204 ],
   alphaCSR[ 101 ][ 205 ],
   alphaCSR[ 101 ][ 206 ],
   alphaCSR[ 101 ][ 207 ],
   alphaCSR[ 101 ][ 208 ],
   alphaCSR[ 101 ][ 209 ],
   alphaCSR[ 101 ][ 210 ],
   alphaCSR[ 101 ][ 211 ],
   alphaCSR[ 101 ][ 212 ],
   alphaCSR[ 101 ][ 213 ],
   alphaCSR[ 101 ][ 214 ],
   alphaCSR[ 101 ][ 215 ],
   alphaCSR[ 101 ][ 216 ],
   alphaCSR[ 101 ][ 217 ],
   alphaCSR[ 101 ][ 218 ],
   alphaCSR[ 101 ][ 219 ],
   alphaCSR[ 101 ][ 220 ],
   alphaCSR[ 101 ][ 221 ],
   alphaCSR[ 101 ][ 222 ],
   alphaCSR[ 101 ][ 223 ],
   alphaCSR[ 101 ][ 224 ],
   alphaCSR[ 101 ][ 225 ],
   alphaCSR[ 101 ][ 226 ],
   alphaCSR[ 101 ][ 227 ],
   alphaCSR[ 101 ][ 228 ],
   alphaCSR[ 101 ][ 229 ],
   alphaCSR[ 101 ][ 230 ],
   alphaCSR[ 101 ][ 231 ],
   alphaCSR[ 101 ][ 232 ],
   alphaCSR[ 101 ][ 233 ],
   alphaCSR[ 101 ][ 234 ],
   alphaCSR[ 101 ][ 235 ],
   alphaCSR[ 101 ][ 236 ],
   alphaCSR[ 101 ][ 237 ],
   alphaCSR[ 101 ][ 238 ],
   alphaCSR[ 101 ][ 239 ],
   alphaCSR[ 101 ][ 240 ],
   alphaCSR[ 101 ][ 241 ],
   alphaCSR[ 101 ][ 242 ],
   alphaCSR[ 101 ][ 243 ],
   alphaCSR[ 101 ][ 244 ],
   alphaCSR[ 101 ][ 245 ],
   alphaCSR[ 101 ][ 246 ],
   alphaCSR[ 101 ][ 247 ],
   alphaCSR[ 101 ][ 248 ],
   alphaCSR[ 101 ][ 249 ],
   alphaCSR[ 101 ][ 250 ],
   alphaCSR[ 101 ][ 251 ],
   alphaCSR[ 101 ][ 252 ],
   alphaCSR[ 101 ][ 253 ],
   alphaCSR[ 101 ][ 254 ],
   alphaCSR[ 101 ][ 255 ],
   alphaCSR[ 101 ][ 256 ],
   alphaCSR[ 101 ][ 257 ],
   alphaCSR[ 101 ][ 258 ],
   alphaCSR[ 101 ][ 259 ],
   alphaCSR[ 101 ][ 260 ],
   alphaCSR[ 101 ][ 261 ],
   alphaCSR[ 101 ][ 262 ],
   alphaCSR[ 101 ][ 263 ],
   alphaCSR[ 101 ][ 264 ],
   alphaCSR[ 101 ][ 265 ],
   alphaCSR[ 101 ][ 266 ],
   alphaCSR[ 101 ][ 267 ],
   alphaCSR[ 101 ][ 268 ],
   alphaCSR[ 101 ][ 269 ],
   alphaCSR[ 101 ][ 270 ],
   alphaCSR[ 101 ][ 271 ],
   alphaCSR[ 101 ][ 272 ],
   alphaCSR[ 101 ][ 273 ],
   alphaCSR[ 101 ][ 274 ],
   alphaCSR[ 101 ][ 275 ],
   alphaCSR[ 101 ][ 276 ],
   alphaCSR[ 101 ][ 277 ],
   alphaCSR[ 101 ][ 278 ],
   alphaCSR[ 101 ][ 279 ],
   alphaCSR[ 101 ][ 280 ],
   alphaCSR[ 101 ][ 281 ],
   alphaCSR[ 101 ][ 282 ],
   alphaCSR[ 101 ][ 283 ],
   alphaCSR[ 101 ][ 284 ],
   alphaCSR[ 101 ][ 285 ],
   alphaCSR[ 101 ][ 286 ],
   alphaCSR[ 101 ][ 287 ],
   alphaCSR[ 101 ][ 288 ],
   alphaCSR[ 101 ][ 289 ],
   alphaCSR[ 101 ][ 290 ],
   alphaCSR[ 101 ][ 291 ],
   alphaCSR[ 101 ][ 292 ],
   alphaCSR[ 101 ][ 293 ],
   alphaCSR[ 101 ][ 294 ],
   alphaCSR[ 101 ][ 295 ],
   alphaCSR[ 101 ][ 296 ],
   alphaCSR[ 101 ][ 297 ],
   alphaCSR[ 101 ][ 298 ],
   alphaCSR[ 101 ][ 299 ],
   alphaCSR[ 101 ][ 300 ],
   alphaCSR[ 101 ][ 301 ],
   alphaCSR[ 101 ][ 302 ],
   alphaCSR[ 101 ][ 303 ],
   alphaCSR[ 101 ][ 304 ],
   alphaCSR[ 101 ][ 305 ],
   alphaCSR[ 101 ][ 306 ],
   alphaCSR[ 101 ][ 307 ],
   alphaCSR[ 101 ][ 308 ],
   alphaCSR[ 101 ][ 309 ],
   alphaCSR[ 101 ][ 310 ],
   alphaCSR[ 101 ][ 311 ],
   alphaCSR[ 101 ][ 312 ],
   alphaCSR[ 101 ][ 313 ],
   alphaCSR[ 101 ][ 314 ],
   alphaCSR[ 101 ][ 315 ],
   alphaCSR[ 101 ][ 316 ],
   alphaCSR[ 101 ][ 317 ],
   alphaCSR[ 101 ][ 318 ],
   alphaCSR[ 101 ][ 319 ],
   alphaCSR[ 101 ][ 320 ],
   alphaCSR[ 101 ][ 321 ],
   alphaCSR[ 101 ][ 322 ],
   alphaCSR[ 101 ][ 323 ],
   alphaCSR[ 101 ][ 324 ],
   alphaCSR[ 101 ][ 325 ],
   alphaCSR[ 101 ][ 326 ],
   alphaCSR[ 101 ][ 327 ],
   alphaCSR[ 101 ][ 328 ],
   alphaCSR[ 101 ][ 329 ],
   alphaCSR[ 101 ][ 330 ],
   alphaCSR[ 101 ][ 331 ],
   alphaCSR[ 101 ][ 332 ],
   alphaCSR[ 101 ][ 333 ],
   alphaCSR[ 101 ][ 334 ],
   alphaCSR[ 101 ][ 335 ],
   alphaCSR[ 101 ][ 336 ],
   alphaCSR[ 101 ][ 337 ],
   alphaCSR[ 101 ][ 338 ],
   alphaCSR[ 101 ][ 339 ],
   alphaCSR[ 101 ][ 340 ],
   alphaCSR[ 101 ][ 341 ],
   alphaCSR[ 101 ][ 342 ],
   alphaCSR[ 101 ][ 343 ],
   alphaCSR[ 101 ][ 344 ],
   alphaCSR[ 101 ][ 345 ],
   alphaCSR[ 101 ][ 346 ],
   alphaCSR[ 101 ][ 347 ],
   alphaCSR[ 101 ][ 348 ],
   alphaCSR[ 101 ][ 349 ],
   alphaCSR[ 101 ][ 350 ],
   alphaCSR[ 101 ][ 351 ],
   alphaCSR[ 101 ][ 352 ],
   alphaCSR[ 101 ][ 353 ],
   alphaCSR[ 101 ][ 354 ],
   alphaCSR[ 101 ][ 355 ],
   alphaCSR[ 101 ][ 356 ],
   alphaCSR[ 101 ][ 357 ],
   alphaCSR[ 101 ][ 358 ],
   alphaCSR[ 101 ][ 359 ],
   alphaCSR[ 101 ][ 360 ],
   alphaCSR[ 101 ][ 361 ],
   alphaCSR[ 101 ][ 362 ],
   alphaCSR[ 101 ][ 363 ],
   alphaCSR[ 101 ][ 364 ],
   alphaCSR[ 101 ][ 365 ],
   alphaCSR[ 101 ][ 366 ],
   alphaCSR[ 101 ][ 367 ],
   alphaCSR[ 101 ][ 368 ],
   alphaCSR[ 101 ][ 369 ],
   alphaCSR[ 101 ][ 370 ],
   alphaCSR[ 101 ][ 371 ],
   alphaCSR[ 101 ][ 372 ],
   alphaCSR[ 101 ][ 373 ],
   alphaCSR[ 101 ][ 374 ],
   alphaCSR[ 101 ][ 375 ],
   alphaCSR[ 101 ][ 376 ],
   alphaCSR[ 101 ][ 377 ],
   alphaCSR[ 101 ][ 378 ],
   alphaCSR[ 101 ][ 379 ],
   alphaCSR[ 101 ][ 380 ],
   alphaCSR[ 101 ][ 381 ],
   alphaCSR[ 101 ][ 382 ],
   alphaCSR[ 101 ][ 383 ],
   alphaCSR[ 102 ][ 0 ],
   alphaCSR[ 102 ][ 1 ],
   alphaCSR[ 102 ][ 2 ],
   alphaCSR[ 102 ][ 3 ],
   alphaCSR[ 102 ][ 4 ],
   alphaCSR[ 102 ][ 5 ],
   alphaCSR[ 102 ][ 6 ],
   alphaCSR[ 102 ][ 7 ],
   alphaCSR[ 102 ][ 8 ],
   alphaCSR[ 102 ][ 9 ],
   alphaCSR[ 102 ][ 10 ],
   alphaCSR[ 102 ][ 11 ],
   alphaCSR[ 102 ][ 12 ],
   alphaCSR[ 102 ][ 13 ],
   alphaCSR[ 102 ][ 14 ],
   alphaCSR[ 102 ][ 15 ],
   alphaCSR[ 102 ][ 16 ],
   alphaCSR[ 102 ][ 17 ],
   alphaCSR[ 102 ][ 18 ],
   alphaCSR[ 102 ][ 19 ],
   alphaCSR[ 102 ][ 20 ],
   alphaCSR[ 102 ][ 21 ],
   alphaCSR[ 102 ][ 22 ],
   alphaCSR[ 102 ][ 23 ],
   alphaCSR[ 102 ][ 24 ],
   alphaCSR[ 102 ][ 25 ],
   alphaCSR[ 102 ][ 26 ],
   alphaCSR[ 102 ][ 27 ],
   alphaCSR[ 102 ][ 28 ],
   alphaCSR[ 102 ][ 29 ],
   alphaCSR[ 102 ][ 30 ],
   alphaCSR[ 102 ][ 31 ],
   alphaCSR[ 102 ][ 32 ],
   alphaCSR[ 102 ][ 33 ],
   alphaCSR[ 102 ][ 34 ],
   alphaCSR[ 102 ][ 35 ],
   alphaCSR[ 102 ][ 36 ],
   alphaCSR[ 102 ][ 37 ],
   alphaCSR[ 102 ][ 38 ],
   alphaCSR[ 102 ][ 39 ],
   alphaCSR[ 102 ][ 40 ],
   alphaCSR[ 102 ][ 41 ],
   alphaCSR[ 102 ][ 42 ],
   alphaCSR[ 102 ][ 43 ],
   alphaCSR[ 102 ][ 44 ],
   alphaCSR[ 102 ][ 45 ],
   alphaCSR[ 102 ][ 46 ],
   alphaCSR[ 102 ][ 47 ],
   alphaCSR[ 102 ][ 48 ],
   alphaCSR[ 102 ][ 49 ],
   alphaCSR[ 102 ][ 50 ],
   alphaCSR[ 102 ][ 51 ],
   alphaCSR[ 102 ][ 52 ],
   alphaCSR[ 102 ][ 53 ],
   alphaCSR[ 102 ][ 54 ],
   alphaCSR[ 102 ][ 55 ],
   alphaCSR[ 102 ][ 56 ],
   alphaCSR[ 102 ][ 57 ],
   alphaCSR[ 102 ][ 58 ],
   alphaCSR[ 102 ][ 59 ],
   alphaCSR[ 102 ][ 60 ],
   alphaCSR[ 102 ][ 61 ],
   alphaCSR[ 102 ][ 62 ],
   alphaCSR[ 102 ][ 63 ],
   alphaCSR[ 102 ][ 64 ],
   alphaCSR[ 102 ][ 65 ],
   alphaCSR[ 102 ][ 66 ],
   alphaCSR[ 102 ][ 67 ],
   alphaCSR[ 102 ][ 68 ],
   alphaCSR[ 102 ][ 69 ],
   alphaCSR[ 102 ][ 70 ],
   alphaCSR[ 102 ][ 71 ],
   alphaCSR[ 102 ][ 72 ],
   alphaCSR[ 102 ][ 73 ],
   alphaCSR[ 102 ][ 74 ],
   alphaCSR[ 102 ][ 75 ],
   alphaCSR[ 102 ][ 76 ],
   alphaCSR[ 102 ][ 77 ],
   alphaCSR[ 102 ][ 78 ],
   alphaCSR[ 102 ][ 79 ],
   alphaCSR[ 102 ][ 80 ],
   alphaCSR[ 102 ][ 81 ],
   alphaCSR[ 102 ][ 82 ],
   alphaCSR[ 102 ][ 83 ],
   alphaCSR[ 102 ][ 84 ],
   alphaCSR[ 102 ][ 85 ],
   alphaCSR[ 102 ][ 86 ],
   alphaCSR[ 102 ][ 87 ],
   alphaCSR[ 102 ][ 88 ],
   alphaCSR[ 102 ][ 89 ],
   alphaCSR[ 102 ][ 90 ],
   alphaCSR[ 102 ][ 91 ],
   alphaCSR[ 102 ][ 92 ],
   alphaCSR[ 102 ][ 93 ],
   alphaCSR[ 102 ][ 94 ],
   alphaCSR[ 102 ][ 95 ],
   alphaCSR[ 102 ][ 96 ],
   alphaCSR[ 102 ][ 97 ],
   alphaCSR[ 102 ][ 98 ],
   alphaCSR[ 102 ][ 99 ],
   alphaCSR[ 102 ][ 100 ],
   alphaCSR[ 102 ][ 101 ],
   alphaCSR[ 102 ][ 102 ],
   alphaCSR[ 102 ][ 103 ],
   alphaCSR[ 102 ][ 104 ],
   alphaCSR[ 102 ][ 105 ],
   alphaCSR[ 102 ][ 106 ],
   alphaCSR[ 102 ][ 107 ],
   alphaCSR[ 102 ][ 108 ],
   alphaCSR[ 102 ][ 109 ],
   alphaCSR[ 102 ][ 110 ],
   alphaCSR[ 102 ][ 111 ],
   alphaCSR[ 102 ][ 112 ],
   alphaCSR[ 102 ][ 113 ],
   alphaCSR[ 102 ][ 114 ],
   alphaCSR[ 102 ][ 115 ],
   alphaCSR[ 102 ][ 116 ],
   alphaCSR[ 102 ][ 117 ],
   alphaCSR[ 102 ][ 118 ],
   alphaCSR[ 102 ][ 119 ],
   alphaCSR[ 102 ][ 120 ],
   alphaCSR[ 102 ][ 121 ],
   alphaCSR[ 102 ][ 122 ],
   alphaCSR[ 102 ][ 123 ],
   alphaCSR[ 102 ][ 124 ],
   alphaCSR[ 102 ][ 125 ],
   alphaCSR[ 102 ][ 126 ],
   alphaCSR[ 102 ][ 127 ],
   alphaCSR[ 102 ][ 128 ],
   alphaCSR[ 102 ][ 129 ],
   alphaCSR[ 102 ][ 130 ],
   alphaCSR[ 102 ][ 131 ],
   alphaCSR[ 102 ][ 132 ],
   alphaCSR[ 102 ][ 133 ],
   alphaCSR[ 102 ][ 134 ],
   alphaCSR[ 102 ][ 135 ],
   alphaCSR[ 102 ][ 136 ],
   alphaCSR[ 102 ][ 137 ],
   alphaCSR[ 102 ][ 138 ],
   alphaCSR[ 102 ][ 139 ],
   alphaCSR[ 102 ][ 140 ],
   alphaCSR[ 102 ][ 141 ],
   alphaCSR[ 102 ][ 142 ],
   alphaCSR[ 102 ][ 143 ],
   alphaCSR[ 102 ][ 144 ],
   alphaCSR[ 102 ][ 145 ],
   alphaCSR[ 102 ][ 146 ],
   alphaCSR[ 102 ][ 147 ],
   alphaCSR[ 102 ][ 148 ],
   alphaCSR[ 102 ][ 149 ],
   alphaCSR[ 102 ][ 150 ],
   alphaCSR[ 102 ][ 151 ],
   alphaCSR[ 102 ][ 152 ],
   alphaCSR[ 102 ][ 153 ],
   alphaCSR[ 102 ][ 154 ],
   alphaCSR[ 102 ][ 155 ],
   alphaCSR[ 102 ][ 156 ],
   alphaCSR[ 102 ][ 157 ],
   alphaCSR[ 102 ][ 158 ],
   alphaCSR[ 102 ][ 159 ],
   alphaCSR[ 102 ][ 160 ],
   alphaCSR[ 102 ][ 161 ],
   alphaCSR[ 102 ][ 162 ],
   alphaCSR[ 102 ][ 163 ],
   alphaCSR[ 102 ][ 164 ],
   alphaCSR[ 102 ][ 165 ],
   alphaCSR[ 102 ][ 166 ],
   alphaCSR[ 102 ][ 167 ],
   alphaCSR[ 102 ][ 168 ],
   alphaCSR[ 102 ][ 169 ],
   alphaCSR[ 102 ][ 170 ],
   alphaCSR[ 102 ][ 171 ],
   alphaCSR[ 102 ][ 172 ],
   alphaCSR[ 102 ][ 173 ],
   alphaCSR[ 102 ][ 174 ],
   alphaCSR[ 102 ][ 175 ],
   alphaCSR[ 102 ][ 176 ],
   alphaCSR[ 102 ][ 177 ],
   alphaCSR[ 102 ][ 178 ],
   alphaCSR[ 102 ][ 179 ],
   alphaCSR[ 102 ][ 180 ],
   alphaCSR[ 102 ][ 181 ],
   alphaCSR[ 102 ][ 182 ],
   alphaCSR[ 102 ][ 183 ],
   alphaCSR[ 102 ][ 184 ],
   alphaCSR[ 102 ][ 185 ],
   alphaCSR[ 102 ][ 186 ],
   alphaCSR[ 102 ][ 187 ],
   alphaCSR[ 102 ][ 188 ],
   alphaCSR[ 102 ][ 189 ],
   alphaCSR[ 102 ][ 190 ],
   alphaCSR[ 102 ][ 191 ],
   alphaCSR[ 102 ][ 192 ],
   alphaCSR[ 102 ][ 193 ],
   alphaCSR[ 102 ][ 194 ],
   alphaCSR[ 102 ][ 195 ],
   alphaCSR[ 102 ][ 196 ],
   alphaCSR[ 102 ][ 197 ],
   alphaCSR[ 102 ][ 198 ],
   alphaCSR[ 102 ][ 199 ],
   alphaCSR[ 102 ][ 200 ],
   alphaCSR[ 102 ][ 201 ],
   alphaCSR[ 102 ][ 202 ],
   alphaCSR[ 102 ][ 203 ],
   alphaCSR[ 102 ][ 204 ],
   alphaCSR[ 102 ][ 205 ],
   alphaCSR[ 102 ][ 206 ],
   alphaCSR[ 102 ][ 207 ],
   alphaCSR[ 102 ][ 208 ],
   alphaCSR[ 102 ][ 209 ],
   alphaCSR[ 102 ][ 210 ],
   alphaCSR[ 102 ][ 211 ],
   alphaCSR[ 102 ][ 212 ],
   alphaCSR[ 102 ][ 213 ],
   alphaCSR[ 102 ][ 214 ],
   alphaCSR[ 102 ][ 215 ],
   alphaCSR[ 102 ][ 216 ],
   alphaCSR[ 102 ][ 217 ],
   alphaCSR[ 102 ][ 218 ],
   alphaCSR[ 102 ][ 219 ],
   alphaCSR[ 102 ][ 220 ],
   alphaCSR[ 102 ][ 221 ],
   alphaCSR[ 102 ][ 222 ],
   alphaCSR[ 102 ][ 223 ],
   alphaCSR[ 102 ][ 224 ],
   alphaCSR[ 102 ][ 225 ],
   alphaCSR[ 102 ][ 226 ],
   alphaCSR[ 102 ][ 227 ],
   alphaCSR[ 102 ][ 228 ],
   alphaCSR[ 102 ][ 229 ],
   alphaCSR[ 102 ][ 230 ],
   alphaCSR[ 102 ][ 231 ],
   alphaCSR[ 102 ][ 232 ],
   alphaCSR[ 102 ][ 233 ],
   alphaCSR[ 102 ][ 234 ],
   alphaCSR[ 102 ][ 235 ],
   alphaCSR[ 102 ][ 236 ],
   alphaCSR[ 102 ][ 237 ],
   alphaCSR[ 102 ][ 238 ],
   alphaCSR[ 102 ][ 239 ],
   alphaCSR[ 102 ][ 240 ],
   alphaCSR[ 102 ][ 241 ],
   alphaCSR[ 102 ][ 242 ],
   alphaCSR[ 102 ][ 243 ],
   alphaCSR[ 102 ][ 244 ],
   alphaCSR[ 102 ][ 245 ],
   alphaCSR[ 102 ][ 246 ],
   alphaCSR[ 102 ][ 247 ],
   alphaCSR[ 102 ][ 248 ],
   alphaCSR[ 102 ][ 249 ],
   alphaCSR[ 102 ][ 250 ],
   alphaCSR[ 102 ][ 251 ],
   alphaCSR[ 102 ][ 252 ],
   alphaCSR[ 102 ][ 253 ],
   alphaCSR[ 102 ][ 254 ],
   alphaCSR[ 102 ][ 255 ],
   alphaCSR[ 102 ][ 256 ],
   alphaCSR[ 102 ][ 257 ],
   alphaCSR[ 102 ][ 258 ],
   alphaCSR[ 102 ][ 259 ],
   alphaCSR[ 102 ][ 260 ],
   alphaCSR[ 102 ][ 261 ],
   alphaCSR[ 102 ][ 262 ],
   alphaCSR[ 102 ][ 263 ],
   alphaCSR[ 102 ][ 264 ],
   alphaCSR[ 102 ][ 265 ],
   alphaCSR[ 102 ][ 266 ],
   alphaCSR[ 102 ][ 267 ],
   alphaCSR[ 102 ][ 268 ],
   alphaCSR[ 102 ][ 269 ],
   alphaCSR[ 102 ][ 270 ],
   alphaCSR[ 102 ][ 271 ],
   alphaCSR[ 102 ][ 272 ],
   alphaCSR[ 102 ][ 273 ],
   alphaCSR[ 102 ][ 274 ],
   alphaCSR[ 102 ][ 275 ],
   alphaCSR[ 102 ][ 276 ],
   alphaCSR[ 102 ][ 277 ],
   alphaCSR[ 102 ][ 278 ],
   alphaCSR[ 102 ][ 279 ],
   alphaCSR[ 102 ][ 280 ],
   alphaCSR[ 102 ][ 281 ],
   alphaCSR[ 102 ][ 282 ],
   alphaCSR[ 102 ][ 283 ],
   alphaCSR[ 102 ][ 284 ],
   alphaCSR[ 102 ][ 285 ],
   alphaCSR[ 102 ][ 286 ],
   alphaCSR[ 102 ][ 287 ],
   alphaCSR[ 102 ][ 288 ],
   alphaCSR[ 102 ][ 289 ],
   alphaCSR[ 102 ][ 290 ],
   alphaCSR[ 102 ][ 291 ],
   alphaCSR[ 102 ][ 292 ],
   alphaCSR[ 102 ][ 293 ],
   alphaCSR[ 102 ][ 294 ],
   alphaCSR[ 102 ][ 295 ],
   alphaCSR[ 102 ][ 296 ],
   alphaCSR[ 102 ][ 297 ],
   alphaCSR[ 102 ][ 298 ],
   alphaCSR[ 102 ][ 299 ],
   alphaCSR[ 102 ][ 300 ],
   alphaCSR[ 102 ][ 301 ],
   alphaCSR[ 102 ][ 302 ],
   alphaCSR[ 102 ][ 303 ],
   alphaCSR[ 102 ][ 304 ],
   alphaCSR[ 102 ][ 305 ],
   alphaCSR[ 102 ][ 306 ],
   alphaCSR[ 102 ][ 307 ],
   alphaCSR[ 102 ][ 308 ],
   alphaCSR[ 102 ][ 309 ],
   alphaCSR[ 102 ][ 310 ],
   alphaCSR[ 102 ][ 311 ],
   alphaCSR[ 102 ][ 312 ],
   alphaCSR[ 102 ][ 313 ],
   alphaCSR[ 102 ][ 314 ],
   alphaCSR[ 102 ][ 315 ],
   alphaCSR[ 102 ][ 316 ],
   alphaCSR[ 102 ][ 317 ],
   alphaCSR[ 102 ][ 318 ],
   alphaCSR[ 102 ][ 319 ],
   alphaCSR[ 102 ][ 320 ],
   alphaCSR[ 102 ][ 321 ],
   alphaCSR[ 102 ][ 322 ],
   alphaCSR[ 102 ][ 323 ],
   alphaCSR[ 102 ][ 324 ],
   alphaCSR[ 102 ][ 325 ],
   alphaCSR[ 102 ][ 326 ],
   alphaCSR[ 102 ][ 327 ],
   alphaCSR[ 102 ][ 328 ],
   alphaCSR[ 102 ][ 329 ],
   alphaCSR[ 102 ][ 330 ],
   alphaCSR[ 102 ][ 331 ],
   alphaCSR[ 102 ][ 332 ],
   alphaCSR[ 102 ][ 333 ],
   alphaCSR[ 102 ][ 334 ],
   alphaCSR[ 102 ][ 335 ],
   alphaCSR[ 102 ][ 336 ],
   alphaCSR[ 102 ][ 337 ],
   alphaCSR[ 102 ][ 338 ],
   alphaCSR[ 102 ][ 339 ],
   alphaCSR[ 102 ][ 340 ],
   alphaCSR[ 102 ][ 341 ],
   alphaCSR[ 102 ][ 342 ],
   alphaCSR[ 102 ][ 343 ],
   alphaCSR[ 102 ][ 344 ],
   alphaCSR[ 102 ][ 345 ],
   alphaCSR[ 102 ][ 346 ],
   alphaCSR[ 102 ][ 347 ],
   alphaCSR[ 102 ][ 348 ],
   alphaCSR[ 102 ][ 349 ],
   alphaCSR[ 102 ][ 350 ],
   alphaCSR[ 102 ][ 351 ],
   alphaCSR[ 102 ][ 352 ],
   alphaCSR[ 102 ][ 353 ],
   alphaCSR[ 102 ][ 354 ],
   alphaCSR[ 102 ][ 355 ],
   alphaCSR[ 102 ][ 356 ],
   alphaCSR[ 102 ][ 357 ],
   alphaCSR[ 102 ][ 358 ],
   alphaCSR[ 102 ][ 359 ],
   alphaCSR[ 102 ][ 360 ],
   alphaCSR[ 102 ][ 361 ],
   alphaCSR[ 102 ][ 362 ],
   alphaCSR[ 102 ][ 363 ],
   alphaCSR[ 102 ][ 364 ],
   alphaCSR[ 102 ][ 365 ],
   alphaCSR[ 102 ][ 366 ],
   alphaCSR[ 102 ][ 367 ],
   alphaCSR[ 102 ][ 368 ],
   alphaCSR[ 102 ][ 369 ],
   alphaCSR[ 102 ][ 370 ],
   alphaCSR[ 102 ][ 371 ],
   alphaCSR[ 102 ][ 372 ],
   alphaCSR[ 102 ][ 373 ],
   alphaCSR[ 102 ][ 374 ],
   alphaCSR[ 102 ][ 375 ],
   alphaCSR[ 102 ][ 376 ],
   alphaCSR[ 102 ][ 377 ],
   alphaCSR[ 102 ][ 378 ],
   alphaCSR[ 102 ][ 379 ],
   alphaCSR[ 102 ][ 380 ],
   alphaCSR[ 102 ][ 381 ],
   alphaCSR[ 102 ][ 382 ],
   alphaCSR[ 102 ][ 383 ],
   alphaCSR[ 103 ][ 0 ],
   alphaCSR[ 103 ][ 1 ],
   alphaCSR[ 103 ][ 2 ],
   alphaCSR[ 103 ][ 3 ],
   alphaCSR[ 103 ][ 4 ],
   alphaCSR[ 103 ][ 5 ],
   alphaCSR[ 103 ][ 6 ],
   alphaCSR[ 103 ][ 7 ],
   alphaCSR[ 103 ][ 8 ],
   alphaCSR[ 103 ][ 9 ],
   alphaCSR[ 103 ][ 10 ],
   alphaCSR[ 103 ][ 11 ],
   alphaCSR[ 103 ][ 12 ],
   alphaCSR[ 103 ][ 13 ],
   alphaCSR[ 103 ][ 14 ],
   alphaCSR[ 103 ][ 15 ],
   alphaCSR[ 103 ][ 16 ],
   alphaCSR[ 103 ][ 17 ],
   alphaCSR[ 103 ][ 18 ],
   alphaCSR[ 103 ][ 19 ],
   alphaCSR[ 103 ][ 20 ],
   alphaCSR[ 103 ][ 21 ],
   alphaCSR[ 103 ][ 22 ],
   alphaCSR[ 103 ][ 23 ],
   alphaCSR[ 103 ][ 24 ],
   alphaCSR[ 103 ][ 25 ],
   alphaCSR[ 103 ][ 26 ],
   alphaCSR[ 103 ][ 27 ],
   alphaCSR[ 103 ][ 28 ],
   alphaCSR[ 103 ][ 29 ],
   alphaCSR[ 103 ][ 30 ],
   alphaCSR[ 103 ][ 31 ],
   alphaCSR[ 103 ][ 32 ],
   alphaCSR[ 103 ][ 33 ],
   alphaCSR[ 103 ][ 34 ],
   alphaCSR[ 103 ][ 35 ],
   alphaCSR[ 103 ][ 36 ],
   alphaCSR[ 103 ][ 37 ],
   alphaCSR[ 103 ][ 38 ],
   alphaCSR[ 103 ][ 39 ],
   alphaCSR[ 103 ][ 40 ],
   alphaCSR[ 103 ][ 41 ],
   alphaCSR[ 103 ][ 42 ],
   alphaCSR[ 103 ][ 43 ],
   alphaCSR[ 103 ][ 44 ],
   alphaCSR[ 103 ][ 45 ],
   alphaCSR[ 103 ][ 46 ],
   alphaCSR[ 103 ][ 47 ],
   alphaCSR[ 103 ][ 48 ],
   alphaCSR[ 103 ][ 49 ],
   alphaCSR[ 103 ][ 50 ],
   alphaCSR[ 103 ][ 51 ],
   alphaCSR[ 103 ][ 52 ],
   alphaCSR[ 103 ][ 53 ],
   alphaCSR[ 103 ][ 54 ],
   alphaCSR[ 103 ][ 55 ],
   alphaCSR[ 103 ][ 56 ],
   alphaCSR[ 103 ][ 57 ],
   alphaCSR[ 103 ][ 58 ],
   alphaCSR[ 103 ][ 59 ],
   alphaCSR[ 103 ][ 60 ],
   alphaCSR[ 103 ][ 61 ],
   alphaCSR[ 103 ][ 62 ],
   alphaCSR[ 103 ][ 63 ],
   alphaCSR[ 103 ][ 64 ],
   alphaCSR[ 103 ][ 65 ],
   alphaCSR[ 103 ][ 66 ],
   alphaCSR[ 103 ][ 67 ],
   alphaCSR[ 103 ][ 68 ],
   alphaCSR[ 103 ][ 69 ],
   alphaCSR[ 103 ][ 70 ],
   alphaCSR[ 103 ][ 71 ],
   alphaCSR[ 103 ][ 72 ],
   alphaCSR[ 103 ][ 73 ],
   alphaCSR[ 103 ][ 74 ],
   alphaCSR[ 103 ][ 75 ],
   alphaCSR[ 103 ][ 76 ],
   alphaCSR[ 103 ][ 77 ],
   alphaCSR[ 103 ][ 78 ],
   alphaCSR[ 103 ][ 79 ],
   alphaCSR[ 103 ][ 80 ],
   alphaCSR[ 103 ][ 81 ],
   alphaCSR[ 103 ][ 82 ],
   alphaCSR[ 103 ][ 83 ],
   alphaCSR[ 103 ][ 84 ],
   alphaCSR[ 103 ][ 85 ],
   alphaCSR[ 103 ][ 86 ],
   alphaCSR[ 103 ][ 87 ],
   alphaCSR[ 103 ][ 88 ],
   alphaCSR[ 103 ][ 89 ],
   alphaCSR[ 103 ][ 90 ],
   alphaCSR[ 103 ][ 91 ],
   alphaCSR[ 103 ][ 92 ],
   alphaCSR[ 103 ][ 93 ],
   alphaCSR[ 103 ][ 94 ],
   alphaCSR[ 103 ][ 95 ],
   alphaCSR[ 103 ][ 96 ],
   alphaCSR[ 103 ][ 97 ],
   alphaCSR[ 103 ][ 98 ],
   alphaCSR[ 103 ][ 99 ],
   alphaCSR[ 103 ][ 100 ],
   alphaCSR[ 103 ][ 101 ],
   alphaCSR[ 103 ][ 102 ],
   alphaCSR[ 103 ][ 103 ],
   alphaCSR[ 103 ][ 104 ],
   alphaCSR[ 103 ][ 105 ],
   alphaCSR[ 103 ][ 106 ],
   alphaCSR[ 103 ][ 107 ],
   alphaCSR[ 103 ][ 108 ],
   alphaCSR[ 103 ][ 109 ],
   alphaCSR[ 103 ][ 110 ],
   alphaCSR[ 103 ][ 111 ],
   alphaCSR[ 103 ][ 112 ],
   alphaCSR[ 103 ][ 113 ],
   alphaCSR[ 103 ][ 114 ],
   alphaCSR[ 103 ][ 115 ],
   alphaCSR[ 103 ][ 116 ],
   alphaCSR[ 103 ][ 117 ],
   alphaCSR[ 103 ][ 118 ],
   alphaCSR[ 103 ][ 119 ],
   alphaCSR[ 103 ][ 120 ],
   alphaCSR[ 103 ][ 121 ],
   alphaCSR[ 103 ][ 122 ],
   alphaCSR[ 103 ][ 123 ],
   alphaCSR[ 103 ][ 124 ],
   alphaCSR[ 103 ][ 125 ],
   alphaCSR[ 103 ][ 126 ],
   alphaCSR[ 103 ][ 127 ],
   alphaCSR[ 103 ][ 128 ],
   alphaCSR[ 103 ][ 129 ],
   alphaCSR[ 103 ][ 130 ],
   alphaCSR[ 103 ][ 131 ],
   alphaCSR[ 103 ][ 132 ],
   alphaCSR[ 103 ][ 133 ],
   alphaCSR[ 103 ][ 134 ],
   alphaCSR[ 103 ][ 135 ],
   alphaCSR[ 103 ][ 136 ],
   alphaCSR[ 103 ][ 137 ],
   alphaCSR[ 103 ][ 138 ],
   alphaCSR[ 103 ][ 139 ],
   alphaCSR[ 103 ][ 140 ],
   alphaCSR[ 103 ][ 141 ],
   alphaCSR[ 103 ][ 142 ],
   alphaCSR[ 103 ][ 143 ],
   alphaCSR[ 103 ][ 144 ],
   alphaCSR[ 103 ][ 145 ],
   alphaCSR[ 103 ][ 146 ],
   alphaCSR[ 103 ][ 147 ],
   alphaCSR[ 103 ][ 148 ],
   alphaCSR[ 103 ][ 149 ],
   alphaCSR[ 103 ][ 150 ],
   alphaCSR[ 103 ][ 151 ],
   alphaCSR[ 103 ][ 152 ],
   alphaCSR[ 103 ][ 153 ],
   alphaCSR[ 103 ][ 154 ],
   alphaCSR[ 103 ][ 155 ],
   alphaCSR[ 103 ][ 156 ],
   alphaCSR[ 103 ][ 157 ],
   alphaCSR[ 103 ][ 158 ],
   alphaCSR[ 103 ][ 159 ],
   alphaCSR[ 103 ][ 160 ],
   alphaCSR[ 103 ][ 161 ],
   alphaCSR[ 103 ][ 162 ],
   alphaCSR[ 103 ][ 163 ],
   alphaCSR[ 103 ][ 164 ],
   alphaCSR[ 103 ][ 165 ],
   alphaCSR[ 103 ][ 166 ],
   alphaCSR[ 103 ][ 167 ],
   alphaCSR[ 103 ][ 168 ],
   alphaCSR[ 103 ][ 169 ],
   alphaCSR[ 103 ][ 170 ],
   alphaCSR[ 103 ][ 171 ],
   alphaCSR[ 103 ][ 172 ],
   alphaCSR[ 103 ][ 173 ],
   alphaCSR[ 103 ][ 174 ],
   alphaCSR[ 103 ][ 175 ],
   alphaCSR[ 103 ][ 176 ],
   alphaCSR[ 103 ][ 177 ],
   alphaCSR[ 103 ][ 178 ],
   alphaCSR[ 103 ][ 179 ],
   alphaCSR[ 103 ][ 180 ],
   alphaCSR[ 103 ][ 181 ],
   alphaCSR[ 103 ][ 182 ],
   alphaCSR[ 103 ][ 183 ],
   alphaCSR[ 103 ][ 184 ],
   alphaCSR[ 103 ][ 185 ],
   alphaCSR[ 103 ][ 186 ],
   alphaCSR[ 103 ][ 187 ],
   alphaCSR[ 103 ][ 188 ],
   alphaCSR[ 103 ][ 189 ],
   alphaCSR[ 103 ][ 190 ],
   alphaCSR[ 103 ][ 191 ],
   alphaCSR[ 103 ][ 192 ],
   alphaCSR[ 103 ][ 193 ],
   alphaCSR[ 103 ][ 194 ],
   alphaCSR[ 103 ][ 195 ],
   alphaCSR[ 103 ][ 196 ],
   alphaCSR[ 103 ][ 197 ],
   alphaCSR[ 103 ][ 198 ],
   alphaCSR[ 103 ][ 199 ],
   alphaCSR[ 103 ][ 200 ],
   alphaCSR[ 103 ][ 201 ],
   alphaCSR[ 103 ][ 202 ],
   alphaCSR[ 103 ][ 203 ],
   alphaCSR[ 103 ][ 204 ],
   alphaCSR[ 103 ][ 205 ],
   alphaCSR[ 103 ][ 206 ],
   alphaCSR[ 103 ][ 207 ],
   alphaCSR[ 103 ][ 208 ],
   alphaCSR[ 103 ][ 209 ],
   alphaCSR[ 103 ][ 210 ],
   alphaCSR[ 103 ][ 211 ],
   alphaCSR[ 103 ][ 212 ],
   alphaCSR[ 103 ][ 213 ],
   alphaCSR[ 103 ][ 214 ],
   alphaCSR[ 103 ][ 215 ],
   alphaCSR[ 103 ][ 216 ],
   alphaCSR[ 103 ][ 217 ],
   alphaCSR[ 103 ][ 218 ],
   alphaCSR[ 103 ][ 219 ],
   alphaCSR[ 103 ][ 220 ],
   alphaCSR[ 103 ][ 221 ],
   alphaCSR[ 103 ][ 222 ],
   alphaCSR[ 103 ][ 223 ],
   alphaCSR[ 103 ][ 224 ],
   alphaCSR[ 103 ][ 225 ],
   alphaCSR[ 103 ][ 226 ],
   alphaCSR[ 103 ][ 227 ],
   alphaCSR[ 103 ][ 228 ],
   alphaCSR[ 103 ][ 229 ],
   alphaCSR[ 103 ][ 230 ],
   alphaCSR[ 103 ][ 231 ],
   alphaCSR[ 103 ][ 232 ],
   alphaCSR[ 103 ][ 233 ],
   alphaCSR[ 103 ][ 234 ],
   alphaCSR[ 103 ][ 235 ],
   alphaCSR[ 103 ][ 236 ],
   alphaCSR[ 103 ][ 237 ],
   alphaCSR[ 103 ][ 238 ],
   alphaCSR[ 103 ][ 239 ],
   alphaCSR[ 103 ][ 240 ],
   alphaCSR[ 103 ][ 241 ],
   alphaCSR[ 103 ][ 242 ],
   alphaCSR[ 103 ][ 243 ],
   alphaCSR[ 103 ][ 244 ],
   alphaCSR[ 103 ][ 245 ],
   alphaCSR[ 103 ][ 246 ],
   alphaCSR[ 103 ][ 247 ],
   alphaCSR[ 103 ][ 248 ],
   alphaCSR[ 103 ][ 249 ],
   alphaCSR[ 103 ][ 250 ],
   alphaCSR[ 103 ][ 251 ],
   alphaCSR[ 103 ][ 252 ],
   alphaCSR[ 103 ][ 253 ],
   alphaCSR[ 103 ][ 254 ],
   alphaCSR[ 103 ][ 255 ],
   alphaCSR[ 103 ][ 256 ],
   alphaCSR[ 103 ][ 257 ],
   alphaCSR[ 103 ][ 258 ],
   alphaCSR[ 103 ][ 259 ],
   alphaCSR[ 103 ][ 260 ],
   alphaCSR[ 103 ][ 261 ],
   alphaCSR[ 103 ][ 262 ],
   alphaCSR[ 103 ][ 263 ],
   alphaCSR[ 103 ][ 264 ],
   alphaCSR[ 103 ][ 265 ],
   alphaCSR[ 103 ][ 266 ],
   alphaCSR[ 103 ][ 267 ],
   alphaCSR[ 103 ][ 268 ],
   alphaCSR[ 103 ][ 269 ],
   alphaCSR[ 103 ][ 270 ],
   alphaCSR[ 103 ][ 271 ],
   alphaCSR[ 103 ][ 272 ],
   alphaCSR[ 103 ][ 273 ],
   alphaCSR[ 103 ][ 274 ],
   alphaCSR[ 103 ][ 275 ],
   alphaCSR[ 103 ][ 276 ],
   alphaCSR[ 103 ][ 277 ],
   alphaCSR[ 103 ][ 278 ],
   alphaCSR[ 103 ][ 279 ],
   alphaCSR[ 103 ][ 280 ],
   alphaCSR[ 103 ][ 281 ],
   alphaCSR[ 103 ][ 282 ],
   alphaCSR[ 103 ][ 283 ],
   alphaCSR[ 103 ][ 284 ],
   alphaCSR[ 103 ][ 285 ],
   alphaCSR[ 103 ][ 286 ],
   alphaCSR[ 103 ][ 287 ],
   alphaCSR[ 103 ][ 288 ],
   alphaCSR[ 103 ][ 289 ],
   alphaCSR[ 103 ][ 290 ],
   alphaCSR[ 103 ][ 291 ],
   alphaCSR[ 103 ][ 292 ],
   alphaCSR[ 103 ][ 293 ],
   alphaCSR[ 103 ][ 294 ],
   alphaCSR[ 103 ][ 295 ],
   alphaCSR[ 103 ][ 296 ],
   alphaCSR[ 103 ][ 297 ],
   alphaCSR[ 103 ][ 298 ],
   alphaCSR[ 103 ][ 299 ],
   alphaCSR[ 103 ][ 300 ],
   alphaCSR[ 103 ][ 301 ],
   alphaCSR[ 103 ][ 302 ],
   alphaCSR[ 103 ][ 303 ],
   alphaCSR[ 103 ][ 304 ],
   alphaCSR[ 103 ][ 305 ],
   alphaCSR[ 103 ][ 306 ],
   alphaCSR[ 103 ][ 307 ],
   alphaCSR[ 103 ][ 308 ],
   alphaCSR[ 103 ][ 309 ],
   alphaCSR[ 103 ][ 310 ],
   alphaCSR[ 103 ][ 311 ],
   alphaCSR[ 103 ][ 312 ],
   alphaCSR[ 103 ][ 313 ],
   alphaCSR[ 103 ][ 314 ],
   alphaCSR[ 103 ][ 315 ],
   alphaCSR[ 103 ][ 316 ],
   alphaCSR[ 103 ][ 317 ],
   alphaCSR[ 103 ][ 318 ],
   alphaCSR[ 103 ][ 319 ],
   alphaCSR[ 103 ][ 320 ],
   alphaCSR[ 103 ][ 321 ],
   alphaCSR[ 103 ][ 322 ],
   alphaCSR[ 103 ][ 323 ],
   alphaCSR[ 103 ][ 324 ],
   alphaCSR[ 103 ][ 325 ],
   alphaCSR[ 103 ][ 326 ],
   alphaCSR[ 103 ][ 327 ],
   alphaCSR[ 103 ][ 328 ],
   alphaCSR[ 103 ][ 329 ],
   alphaCSR[ 103 ][ 330 ],
   alphaCSR[ 103 ][ 331 ],
   alphaCSR[ 103 ][ 332 ],
   alphaCSR[ 103 ][ 333 ],
   alphaCSR[ 103 ][ 334 ],
   alphaCSR[ 103 ][ 335 ],
   alphaCSR[ 103 ][ 336 ],
   alphaCSR[ 103 ][ 337 ],
   alphaCSR[ 103 ][ 338 ],
   alphaCSR[ 103 ][ 339 ],
   alphaCSR[ 103 ][ 340 ],
   alphaCSR[ 103 ][ 341 ],
   alphaCSR[ 103 ][ 342 ],
   alphaCSR[ 103 ][ 343 ],
   alphaCSR[ 103 ][ 344 ],
   alphaCSR[ 103 ][ 345 ],
   alphaCSR[ 103 ][ 346 ],
   alphaCSR[ 103 ][ 347 ],
   alphaCSR[ 103 ][ 348 ],
   alphaCSR[ 103 ][ 349 ],
   alphaCSR[ 103 ][ 350 ],
   alphaCSR[ 103 ][ 351 ],
   alphaCSR[ 103 ][ 352 ],
   alphaCSR[ 103 ][ 353 ],
   alphaCSR[ 103 ][ 354 ],
   alphaCSR[ 103 ][ 355 ],
   alphaCSR[ 103 ][ 356 ],
   alphaCSR[ 103 ][ 357 ],
   alphaCSR[ 103 ][ 358 ],
   alphaCSR[ 103 ][ 359 ],
   alphaCSR[ 103 ][ 360 ],
   alphaCSR[ 103 ][ 361 ],
   alphaCSR[ 103 ][ 362 ],
   alphaCSR[ 103 ][ 363 ],
   alphaCSR[ 103 ][ 364 ],
   alphaCSR[ 103 ][ 365 ],
   alphaCSR[ 103 ][ 366 ],
   alphaCSR[ 103 ][ 367 ],
   alphaCSR[ 103 ][ 368 ],
   alphaCSR[ 103 ][ 369 ],
   alphaCSR[ 103 ][ 370 ],
   alphaCSR[ 103 ][ 371 ],
   alphaCSR[ 103 ][ 372 ],
   alphaCSR[ 103 ][ 373 ],
   alphaCSR[ 103 ][ 374 ],
   alphaCSR[ 103 ][ 375 ],
   alphaCSR[ 103 ][ 376 ],
   alphaCSR[ 103 ][ 377 ],
   alphaCSR[ 103 ][ 378 ],
   alphaCSR[ 103 ][ 379 ],
   alphaCSR[ 103 ][ 380 ],
   alphaCSR[ 103 ][ 381 ],
   alphaCSR[ 103 ][ 382 ],
   alphaCSR[ 103 ][ 383 ],
   alphaCSR[ 104 ][ 0 ],
   alphaCSR[ 104 ][ 1 ],
   alphaCSR[ 104 ][ 2 ],
   alphaCSR[ 104 ][ 3 ],
   alphaCSR[ 104 ][ 4 ],
   alphaCSR[ 104 ][ 5 ],
   alphaCSR[ 104 ][ 6 ],
   alphaCSR[ 104 ][ 7 ],
   alphaCSR[ 104 ][ 8 ],
   alphaCSR[ 104 ][ 9 ],
   alphaCSR[ 104 ][ 10 ],
   alphaCSR[ 104 ][ 11 ],
   alphaCSR[ 104 ][ 12 ],
   alphaCSR[ 104 ][ 13 ],
   alphaCSR[ 104 ][ 14 ],
   alphaCSR[ 104 ][ 15 ],
   alphaCSR[ 104 ][ 16 ],
   alphaCSR[ 104 ][ 17 ],
   alphaCSR[ 104 ][ 18 ],
   alphaCSR[ 104 ][ 19 ],
   alphaCSR[ 104 ][ 20 ],
   alphaCSR[ 104 ][ 21 ],
   alphaCSR[ 104 ][ 22 ],
   alphaCSR[ 104 ][ 23 ],
   alphaCSR[ 104 ][ 24 ],
   alphaCSR[ 104 ][ 25 ],
   alphaCSR[ 104 ][ 26 ],
   alphaCSR[ 104 ][ 27 ],
   alphaCSR[ 104 ][ 28 ],
   alphaCSR[ 104 ][ 29 ],
   alphaCSR[ 104 ][ 30 ],
   alphaCSR[ 104 ][ 31 ],
   alphaCSR[ 104 ][ 32 ],
   alphaCSR[ 104 ][ 33 ],
   alphaCSR[ 104 ][ 34 ],
   alphaCSR[ 104 ][ 35 ],
   alphaCSR[ 104 ][ 36 ],
   alphaCSR[ 104 ][ 37 ],
   alphaCSR[ 104 ][ 38 ],
   alphaCSR[ 104 ][ 39 ],
   alphaCSR[ 104 ][ 40 ],
   alphaCSR[ 104 ][ 41 ],
   alphaCSR[ 104 ][ 42 ],
   alphaCSR[ 104 ][ 43 ],
   alphaCSR[ 104 ][ 44 ],
   alphaCSR[ 104 ][ 45 ],
   alphaCSR[ 104 ][ 46 ],
   alphaCSR[ 104 ][ 47 ],
   alphaCSR[ 104 ][ 48 ],
   alphaCSR[ 104 ][ 49 ],
   alphaCSR[ 104 ][ 50 ],
   alphaCSR[ 104 ][ 51 ],
   alphaCSR[ 104 ][ 52 ],
   alphaCSR[ 104 ][ 53 ],
   alphaCSR[ 104 ][ 54 ],
   alphaCSR[ 104 ][ 55 ],
   alphaCSR[ 104 ][ 56 ],
   alphaCSR[ 104 ][ 57 ],
   alphaCSR[ 104 ][ 58 ],
   alphaCSR[ 104 ][ 59 ],
   alphaCSR[ 104 ][ 60 ],
   alphaCSR[ 104 ][ 61 ],
   alphaCSR[ 104 ][ 62 ],
   alphaCSR[ 104 ][ 63 ],
   alphaCSR[ 104 ][ 64 ],
   alphaCSR[ 104 ][ 65 ],
   alphaCSR[ 104 ][ 66 ],
   alphaCSR[ 104 ][ 67 ],
   alphaCSR[ 104 ][ 68 ],
   alphaCSR[ 104 ][ 69 ],
   alphaCSR[ 104 ][ 70 ],
   alphaCSR[ 104 ][ 71 ],
   alphaCSR[ 104 ][ 72 ],
   alphaCSR[ 104 ][ 73 ],
   alphaCSR[ 104 ][ 74 ],
   alphaCSR[ 104 ][ 75 ],
   alphaCSR[ 104 ][ 76 ],
   alphaCSR[ 104 ][ 77 ],
   alphaCSR[ 104 ][ 78 ],
   alphaCSR[ 104 ][ 79 ],
   alphaCSR[ 104 ][ 80 ],
   alphaCSR[ 104 ][ 81 ],
   alphaCSR[ 104 ][ 82 ],
   alphaCSR[ 104 ][ 83 ],
   alphaCSR[ 104 ][ 84 ],
   alphaCSR[ 104 ][ 85 ],
   alphaCSR[ 104 ][ 86 ],
   alphaCSR[ 104 ][ 87 ],
   alphaCSR[ 104 ][ 88 ],
   alphaCSR[ 104 ][ 89 ],
   alphaCSR[ 104 ][ 90 ],
   alphaCSR[ 104 ][ 91 ],
   alphaCSR[ 104 ][ 92 ],
   alphaCSR[ 104 ][ 93 ],
   alphaCSR[ 104 ][ 94 ],
   alphaCSR[ 104 ][ 95 ],
   alphaCSR[ 104 ][ 96 ],
   alphaCSR[ 104 ][ 97 ],
   alphaCSR[ 104 ][ 98 ],
   alphaCSR[ 104 ][ 99 ],
   alphaCSR[ 104 ][ 100 ],
   alphaCSR[ 104 ][ 101 ],
   alphaCSR[ 104 ][ 102 ],
   alphaCSR[ 104 ][ 103 ],
   alphaCSR[ 104 ][ 104 ],
   alphaCSR[ 104 ][ 105 ],
   alphaCSR[ 104 ][ 106 ],
   alphaCSR[ 104 ][ 107 ],
   alphaCSR[ 104 ][ 108 ],
   alphaCSR[ 104 ][ 109 ],
   alphaCSR[ 104 ][ 110 ],
   alphaCSR[ 104 ][ 111 ],
   alphaCSR[ 104 ][ 112 ],
   alphaCSR[ 104 ][ 113 ],
   alphaCSR[ 104 ][ 114 ],
   alphaCSR[ 104 ][ 115 ],
   alphaCSR[ 104 ][ 116 ],
   alphaCSR[ 104 ][ 117 ],
   alphaCSR[ 104 ][ 118 ],
   alphaCSR[ 104 ][ 119 ],
   alphaCSR[ 104 ][ 120 ],
   alphaCSR[ 104 ][ 121 ],
   alphaCSR[ 104 ][ 122 ],
   alphaCSR[ 104 ][ 123 ],
   alphaCSR[ 104 ][ 124 ],
   alphaCSR[ 104 ][ 125 ],
   alphaCSR[ 104 ][ 126 ],
   alphaCSR[ 104 ][ 127 ],
   alphaCSR[ 104 ][ 128 ],
   alphaCSR[ 104 ][ 129 ],
   alphaCSR[ 104 ][ 130 ],
   alphaCSR[ 104 ][ 131 ],
   alphaCSR[ 104 ][ 132 ],
   alphaCSR[ 104 ][ 133 ],
   alphaCSR[ 104 ][ 134 ],
   alphaCSR[ 104 ][ 135 ],
   alphaCSR[ 104 ][ 136 ],
   alphaCSR[ 104 ][ 137 ],
   alphaCSR[ 104 ][ 138 ],
   alphaCSR[ 104 ][ 139 ],
   alphaCSR[ 104 ][ 140 ],
   alphaCSR[ 104 ][ 141 ],
   alphaCSR[ 104 ][ 142 ],
   alphaCSR[ 104 ][ 143 ],
   alphaCSR[ 104 ][ 144 ],
   alphaCSR[ 104 ][ 145 ],
   alphaCSR[ 104 ][ 146 ],
   alphaCSR[ 104 ][ 147 ],
   alphaCSR[ 104 ][ 148 ],
   alphaCSR[ 104 ][ 149 ],
   alphaCSR[ 104 ][ 150 ],
   alphaCSR[ 104 ][ 151 ],
   alphaCSR[ 104 ][ 152 ],
   alphaCSR[ 104 ][ 153 ],
   alphaCSR[ 104 ][ 154 ],
   alphaCSR[ 104 ][ 155 ],
   alphaCSR[ 104 ][ 156 ],
   alphaCSR[ 104 ][ 157 ],
   alphaCSR[ 104 ][ 158 ],
   alphaCSR[ 104 ][ 159 ],
   alphaCSR[ 104 ][ 160 ],
   alphaCSR[ 104 ][ 161 ],
   alphaCSR[ 104 ][ 162 ],
   alphaCSR[ 104 ][ 163 ],
   alphaCSR[ 104 ][ 164 ],
   alphaCSR[ 104 ][ 165 ],
   alphaCSR[ 104 ][ 166 ],
   alphaCSR[ 104 ][ 167 ],
   alphaCSR[ 104 ][ 168 ],
   alphaCSR[ 104 ][ 169 ],
   alphaCSR[ 104 ][ 170 ],
   alphaCSR[ 104 ][ 171 ],
   alphaCSR[ 104 ][ 172 ],
   alphaCSR[ 104 ][ 173 ],
   alphaCSR[ 104 ][ 174 ],
   alphaCSR[ 104 ][ 175 ],
   alphaCSR[ 104 ][ 176 ],
   alphaCSR[ 104 ][ 177 ],
   alphaCSR[ 104 ][ 178 ],
   alphaCSR[ 104 ][ 179 ],
   alphaCSR[ 104 ][ 180 ],
   alphaCSR[ 104 ][ 181 ],
   alphaCSR[ 104 ][ 182 ],
   alphaCSR[ 104 ][ 183 ],
   alphaCSR[ 104 ][ 184 ],
   alphaCSR[ 104 ][ 185 ],
   alphaCSR[ 104 ][ 186 ],
   alphaCSR[ 104 ][ 187 ],
   alphaCSR[ 104 ][ 188 ],
   alphaCSR[ 104 ][ 189 ],
   alphaCSR[ 104 ][ 190 ],
   alphaCSR[ 104 ][ 191 ],
   alphaCSR[ 104 ][ 192 ],
   alphaCSR[ 104 ][ 193 ],
   alphaCSR[ 104 ][ 194 ],
   alphaCSR[ 104 ][ 195 ],
   alphaCSR[ 104 ][ 196 ],
   alphaCSR[ 104 ][ 197 ],
   alphaCSR[ 104 ][ 198 ],
   alphaCSR[ 104 ][ 199 ],
   alphaCSR[ 104 ][ 200 ],
   alphaCSR[ 104 ][ 201 ],
   alphaCSR[ 104 ][ 202 ],
   alphaCSR[ 104 ][ 203 ],
   alphaCSR[ 104 ][ 204 ],
   alphaCSR[ 104 ][ 205 ],
   alphaCSR[ 104 ][ 206 ],
   alphaCSR[ 104 ][ 207 ],
   alphaCSR[ 104 ][ 208 ],
   alphaCSR[ 104 ][ 209 ],
   alphaCSR[ 104 ][ 210 ],
   alphaCSR[ 104 ][ 211 ],
   alphaCSR[ 104 ][ 212 ],
   alphaCSR[ 104 ][ 213 ],
   alphaCSR[ 104 ][ 214 ],
   alphaCSR[ 104 ][ 215 ],
   alphaCSR[ 104 ][ 216 ],
   alphaCSR[ 104 ][ 217 ],
   alphaCSR[ 104 ][ 218 ],
   alphaCSR[ 104 ][ 219 ],
   alphaCSR[ 104 ][ 220 ],
   alphaCSR[ 104 ][ 221 ],
   alphaCSR[ 104 ][ 222 ],
   alphaCSR[ 104 ][ 223 ],
   alphaCSR[ 104 ][ 224 ],
   alphaCSR[ 104 ][ 225 ],
   alphaCSR[ 104 ][ 226 ],
   alphaCSR[ 104 ][ 227 ],
   alphaCSR[ 104 ][ 228 ],
   alphaCSR[ 104 ][ 229 ],
   alphaCSR[ 104 ][ 230 ],
   alphaCSR[ 104 ][ 231 ],
   alphaCSR[ 104 ][ 232 ],
   alphaCSR[ 104 ][ 233 ],
   alphaCSR[ 104 ][ 234 ],
   alphaCSR[ 104 ][ 235 ],
   alphaCSR[ 104 ][ 236 ],
   alphaCSR[ 104 ][ 237 ],
   alphaCSR[ 104 ][ 238 ],
   alphaCSR[ 104 ][ 239 ],
   alphaCSR[ 104 ][ 240 ],
   alphaCSR[ 104 ][ 241 ],
   alphaCSR[ 104 ][ 242 ],
   alphaCSR[ 104 ][ 243 ],
   alphaCSR[ 104 ][ 244 ],
   alphaCSR[ 104 ][ 245 ],
   alphaCSR[ 104 ][ 246 ],
   alphaCSR[ 104 ][ 247 ],
   alphaCSR[ 104 ][ 248 ],
   alphaCSR[ 104 ][ 249 ],
   alphaCSR[ 104 ][ 250 ],
   alphaCSR[ 104 ][ 251 ],
   alphaCSR[ 104 ][ 252 ],
   alphaCSR[ 104 ][ 253 ],
   alphaCSR[ 104 ][ 254 ],
   alphaCSR[ 104 ][ 255 ],
   alphaCSR[ 104 ][ 256 ],
   alphaCSR[ 104 ][ 257 ],
   alphaCSR[ 104 ][ 258 ],
   alphaCSR[ 104 ][ 259 ],
   alphaCSR[ 104 ][ 260 ],
   alphaCSR[ 104 ][ 261 ],
   alphaCSR[ 104 ][ 262 ],
   alphaCSR[ 104 ][ 263 ],
   alphaCSR[ 104 ][ 264 ],
   alphaCSR[ 104 ][ 265 ],
   alphaCSR[ 104 ][ 266 ],
   alphaCSR[ 104 ][ 267 ],
   alphaCSR[ 104 ][ 268 ],
   alphaCSR[ 104 ][ 269 ],
   alphaCSR[ 104 ][ 270 ],
   alphaCSR[ 104 ][ 271 ],
   alphaCSR[ 104 ][ 272 ],
   alphaCSR[ 104 ][ 273 ],
   alphaCSR[ 104 ][ 274 ],
   alphaCSR[ 104 ][ 275 ],
   alphaCSR[ 104 ][ 276 ],
   alphaCSR[ 104 ][ 277 ],
   alphaCSR[ 104 ][ 278 ],
   alphaCSR[ 104 ][ 279 ],
   alphaCSR[ 104 ][ 280 ],
   alphaCSR[ 104 ][ 281 ],
   alphaCSR[ 104 ][ 282 ],
   alphaCSR[ 104 ][ 283 ],
   alphaCSR[ 104 ][ 284 ],
   alphaCSR[ 104 ][ 285 ],
   alphaCSR[ 104 ][ 286 ],
   alphaCSR[ 104 ][ 287 ],
   alphaCSR[ 104 ][ 288 ],
   alphaCSR[ 104 ][ 289 ],
   alphaCSR[ 104 ][ 290 ],
   alphaCSR[ 104 ][ 291 ],
   alphaCSR[ 104 ][ 292 ],
   alphaCSR[ 104 ][ 293 ],
   alphaCSR[ 104 ][ 294 ],
   alphaCSR[ 104 ][ 295 ],
   alphaCSR[ 104 ][ 296 ],
   alphaCSR[ 104 ][ 297 ],
   alphaCSR[ 104 ][ 298 ],
   alphaCSR[ 104 ][ 299 ],
   alphaCSR[ 104 ][ 300 ],
   alphaCSR[ 104 ][ 301 ],
   alphaCSR[ 104 ][ 302 ],
   alphaCSR[ 104 ][ 303 ],
   alphaCSR[ 104 ][ 304 ],
   alphaCSR[ 104 ][ 305 ],
   alphaCSR[ 104 ][ 306 ],
   alphaCSR[ 104 ][ 307 ],
   alphaCSR[ 104 ][ 308 ],
   alphaCSR[ 104 ][ 309 ],
   alphaCSR[ 104 ][ 310 ],
   alphaCSR[ 104 ][ 311 ],
   alphaCSR[ 104 ][ 312 ],
   alphaCSR[ 104 ][ 313 ],
   alphaCSR[ 104 ][ 314 ],
   alphaCSR[ 104 ][ 315 ],
   alphaCSR[ 104 ][ 316 ],
   alphaCSR[ 104 ][ 317 ],
   alphaCSR[ 104 ][ 318 ],
   alphaCSR[ 104 ][ 319 ],
   alphaCSR[ 104 ][ 320 ],
   alphaCSR[ 104 ][ 321 ],
   alphaCSR[ 104 ][ 322 ],
   alphaCSR[ 104 ][ 323 ],
   alphaCSR[ 104 ][ 324 ],
   alphaCSR[ 104 ][ 325 ],
   alphaCSR[ 104 ][ 326 ],
   alphaCSR[ 104 ][ 327 ],
   alphaCSR[ 104 ][ 328 ],
   alphaCSR[ 104 ][ 329 ],
   alphaCSR[ 104 ][ 330 ],
   alphaCSR[ 104 ][ 331 ],
   alphaCSR[ 104 ][ 332 ],
   alphaCSR[ 104 ][ 333 ],
   alphaCSR[ 104 ][ 334 ],
   alphaCSR[ 104 ][ 335 ],
   alphaCSR[ 104 ][ 336 ],
   alphaCSR[ 104 ][ 337 ],
   alphaCSR[ 104 ][ 338 ],
   alphaCSR[ 104 ][ 339 ],
   alphaCSR[ 104 ][ 340 ],
   alphaCSR[ 104 ][ 341 ],
   alphaCSR[ 104 ][ 342 ],
   alphaCSR[ 104 ][ 343 ],
   alphaCSR[ 104 ][ 344 ],
   alphaCSR[ 104 ][ 345 ],
   alphaCSR[ 104 ][ 346 ],
   alphaCSR[ 104 ][ 347 ],
   alphaCSR[ 104 ][ 348 ],
   alphaCSR[ 104 ][ 349 ],
   alphaCSR[ 104 ][ 350 ],
   alphaCSR[ 104 ][ 351 ],
   alphaCSR[ 104 ][ 352 ],
   alphaCSR[ 104 ][ 353 ],
   alphaCSR[ 104 ][ 354 ],
   alphaCSR[ 104 ][ 355 ],
   alphaCSR[ 104 ][ 356 ],
   alphaCSR[ 104 ][ 357 ],
   alphaCSR[ 104 ][ 358 ],
   alphaCSR[ 104 ][ 359 ],
   alphaCSR[ 104 ][ 360 ],
   alphaCSR[ 104 ][ 361 ],
   alphaCSR[ 104 ][ 362 ],
   alphaCSR[ 104 ][ 363 ],
   alphaCSR[ 104 ][ 364 ],
   alphaCSR[ 104 ][ 365 ],
   alphaCSR[ 104 ][ 366 ],
   alphaCSR[ 104 ][ 367 ],
   alphaCSR[ 104 ][ 368 ],
   alphaCSR[ 104 ][ 369 ],
   alphaCSR[ 104 ][ 370 ],
   alphaCSR[ 104 ][ 371 ],
   alphaCSR[ 104 ][ 372 ],
   alphaCSR[ 104 ][ 373 ],
   alphaCSR[ 104 ][ 374 ],
   alphaCSR[ 104 ][ 375 ],
   alphaCSR[ 104 ][ 376 ],
   alphaCSR[ 104 ][ 377 ],
   alphaCSR[ 104 ][ 378 ],
   alphaCSR[ 104 ][ 379 ],
   alphaCSR[ 104 ][ 380 ],
   alphaCSR[ 104 ][ 381 ],
   alphaCSR[ 104 ][ 382 ],
   alphaCSR[ 104 ][ 383 ],
   alphaCSR[ 105 ][ 0 ],
   alphaCSR[ 105 ][ 1 ],
   alphaCSR[ 105 ][ 2 ],
   alphaCSR[ 105 ][ 3 ],
   alphaCSR[ 105 ][ 4 ],
   alphaCSR[ 105 ][ 5 ],
   alphaCSR[ 105 ][ 6 ],
   alphaCSR[ 105 ][ 7 ],
   alphaCSR[ 105 ][ 8 ],
   alphaCSR[ 105 ][ 9 ],
   alphaCSR[ 105 ][ 10 ],
   alphaCSR[ 105 ][ 11 ],
   alphaCSR[ 105 ][ 12 ],
   alphaCSR[ 105 ][ 13 ],
   alphaCSR[ 105 ][ 14 ],
   alphaCSR[ 105 ][ 15 ],
   alphaCSR[ 105 ][ 16 ],
   alphaCSR[ 105 ][ 17 ],
   alphaCSR[ 105 ][ 18 ],
   alphaCSR[ 105 ][ 19 ],
   alphaCSR[ 105 ][ 20 ],
   alphaCSR[ 105 ][ 21 ],
   alphaCSR[ 105 ][ 22 ],
   alphaCSR[ 105 ][ 23 ],
   alphaCSR[ 105 ][ 24 ],
   alphaCSR[ 105 ][ 25 ],
   alphaCSR[ 105 ][ 26 ],
   alphaCSR[ 105 ][ 27 ],
   alphaCSR[ 105 ][ 28 ],
   alphaCSR[ 105 ][ 29 ],
   alphaCSR[ 105 ][ 30 ],
   alphaCSR[ 105 ][ 31 ],
   alphaCSR[ 105 ][ 32 ],
   alphaCSR[ 105 ][ 33 ],
   alphaCSR[ 105 ][ 34 ],
   alphaCSR[ 105 ][ 35 ],
   alphaCSR[ 105 ][ 36 ],
   alphaCSR[ 105 ][ 37 ],
   alphaCSR[ 105 ][ 38 ],
   alphaCSR[ 105 ][ 39 ],
   alphaCSR[ 105 ][ 40 ],
   alphaCSR[ 105 ][ 41 ],
   alphaCSR[ 105 ][ 42 ],
   alphaCSR[ 105 ][ 43 ],
   alphaCSR[ 105 ][ 44 ],
   alphaCSR[ 105 ][ 45 ],
   alphaCSR[ 105 ][ 46 ],
   alphaCSR[ 105 ][ 47 ],
   alphaCSR[ 105 ][ 48 ],
   alphaCSR[ 105 ][ 49 ],
   alphaCSR[ 105 ][ 50 ],
   alphaCSR[ 105 ][ 51 ],
   alphaCSR[ 105 ][ 52 ],
   alphaCSR[ 105 ][ 53 ],
   alphaCSR[ 105 ][ 54 ],
   alphaCSR[ 105 ][ 55 ],
   alphaCSR[ 105 ][ 56 ],
   alphaCSR[ 105 ][ 57 ],
   alphaCSR[ 105 ][ 58 ],
   alphaCSR[ 105 ][ 59 ],
   alphaCSR[ 105 ][ 60 ],
   alphaCSR[ 105 ][ 61 ],
   alphaCSR[ 105 ][ 62 ],
   alphaCSR[ 105 ][ 63 ],
   alphaCSR[ 105 ][ 64 ],
   alphaCSR[ 105 ][ 65 ],
   alphaCSR[ 105 ][ 66 ],
   alphaCSR[ 105 ][ 67 ],
   alphaCSR[ 105 ][ 68 ],
   alphaCSR[ 105 ][ 69 ],
   alphaCSR[ 105 ][ 70 ],
   alphaCSR[ 105 ][ 71 ],
   alphaCSR[ 105 ][ 72 ],
   alphaCSR[ 105 ][ 73 ],
   alphaCSR[ 105 ][ 74 ],
   alphaCSR[ 105 ][ 75 ],
   alphaCSR[ 105 ][ 76 ],
   alphaCSR[ 105 ][ 77 ],
   alphaCSR[ 105 ][ 78 ],
   alphaCSR[ 105 ][ 79 ],
   alphaCSR[ 105 ][ 80 ],
   alphaCSR[ 105 ][ 81 ],
   alphaCSR[ 105 ][ 82 ],
   alphaCSR[ 105 ][ 83 ],
   alphaCSR[ 105 ][ 84 ],
   alphaCSR[ 105 ][ 85 ],
   alphaCSR[ 105 ][ 86 ],
   alphaCSR[ 105 ][ 87 ],
   alphaCSR[ 105 ][ 88 ],
   alphaCSR[ 105 ][ 89 ],
   alphaCSR[ 105 ][ 90 ],
   alphaCSR[ 105 ][ 91 ],
   alphaCSR[ 105 ][ 92 ],
   alphaCSR[ 105 ][ 93 ],
   alphaCSR[ 105 ][ 94 ],
   alphaCSR[ 105 ][ 95 ],
   alphaCSR[ 105 ][ 96 ],
   alphaCSR[ 105 ][ 97 ],
   alphaCSR[ 105 ][ 98 ],
   alphaCSR[ 105 ][ 99 ],
   alphaCSR[ 105 ][ 100 ],
   alphaCSR[ 105 ][ 101 ],
   alphaCSR[ 105 ][ 102 ],
   alphaCSR[ 105 ][ 103 ],
   alphaCSR[ 105 ][ 104 ],
   alphaCSR[ 105 ][ 105 ],
   alphaCSR[ 105 ][ 106 ],
   alphaCSR[ 105 ][ 107 ],
   alphaCSR[ 105 ][ 108 ],
   alphaCSR[ 105 ][ 109 ],
   alphaCSR[ 105 ][ 110 ],
   alphaCSR[ 105 ][ 111 ],
   alphaCSR[ 105 ][ 112 ],
   alphaCSR[ 105 ][ 113 ],
   alphaCSR[ 105 ][ 114 ],
   alphaCSR[ 105 ][ 115 ],
   alphaCSR[ 105 ][ 116 ],
   alphaCSR[ 105 ][ 117 ],
   alphaCSR[ 105 ][ 118 ],
   alphaCSR[ 105 ][ 119 ],
   alphaCSR[ 105 ][ 120 ],
   alphaCSR[ 105 ][ 121 ],
   alphaCSR[ 105 ][ 122 ],
   alphaCSR[ 105 ][ 123 ],
   alphaCSR[ 105 ][ 124 ],
   alphaCSR[ 105 ][ 125 ],
   alphaCSR[ 105 ][ 126 ],
   alphaCSR[ 105 ][ 127 ],
   alphaCSR[ 105 ][ 128 ],
   alphaCSR[ 105 ][ 129 ],
   alphaCSR[ 105 ][ 130 ],
   alphaCSR[ 105 ][ 131 ],
   alphaCSR[ 105 ][ 132 ],
   alphaCSR[ 105 ][ 133 ],
   alphaCSR[ 105 ][ 134 ],
   alphaCSR[ 105 ][ 135 ],
   alphaCSR[ 105 ][ 136 ],
   alphaCSR[ 105 ][ 137 ],
   alphaCSR[ 105 ][ 138 ],
   alphaCSR[ 105 ][ 139 ],
   alphaCSR[ 105 ][ 140 ],
   alphaCSR[ 105 ][ 141 ],
   alphaCSR[ 105 ][ 142 ],
   alphaCSR[ 105 ][ 143 ],
   alphaCSR[ 105 ][ 144 ],
   alphaCSR[ 105 ][ 145 ],
   alphaCSR[ 105 ][ 146 ],
   alphaCSR[ 105 ][ 147 ],
   alphaCSR[ 105 ][ 148 ],
   alphaCSR[ 105 ][ 149 ],
   alphaCSR[ 105 ][ 150 ],
   alphaCSR[ 105 ][ 151 ],
   alphaCSR[ 105 ][ 152 ],
   alphaCSR[ 105 ][ 153 ],
   alphaCSR[ 105 ][ 154 ],
   alphaCSR[ 105 ][ 155 ],
   alphaCSR[ 105 ][ 156 ],
   alphaCSR[ 105 ][ 157 ],
   alphaCSR[ 105 ][ 158 ],
   alphaCSR[ 105 ][ 159 ],
   alphaCSR[ 105 ][ 160 ],
   alphaCSR[ 105 ][ 161 ],
   alphaCSR[ 105 ][ 162 ],
   alphaCSR[ 105 ][ 163 ],
   alphaCSR[ 105 ][ 164 ],
   alphaCSR[ 105 ][ 165 ],
   alphaCSR[ 105 ][ 166 ],
   alphaCSR[ 105 ][ 167 ],
   alphaCSR[ 105 ][ 168 ],
   alphaCSR[ 105 ][ 169 ],
   alphaCSR[ 105 ][ 170 ],
   alphaCSR[ 105 ][ 171 ],
   alphaCSR[ 105 ][ 172 ],
   alphaCSR[ 105 ][ 173 ],
   alphaCSR[ 105 ][ 174 ],
   alphaCSR[ 105 ][ 175 ],
   alphaCSR[ 105 ][ 176 ],
   alphaCSR[ 105 ][ 177 ],
   alphaCSR[ 105 ][ 178 ],
   alphaCSR[ 105 ][ 179 ],
   alphaCSR[ 105 ][ 180 ],
   alphaCSR[ 105 ][ 181 ],
   alphaCSR[ 105 ][ 182 ],
   alphaCSR[ 105 ][ 183 ],
   alphaCSR[ 105 ][ 184 ],
   alphaCSR[ 105 ][ 185 ],
   alphaCSR[ 105 ][ 186 ],
   alphaCSR[ 105 ][ 187 ],
   alphaCSR[ 105 ][ 188 ],
   alphaCSR[ 105 ][ 189 ],
   alphaCSR[ 105 ][ 190 ],
   alphaCSR[ 105 ][ 191 ],
   alphaCSR[ 105 ][ 192 ],
   alphaCSR[ 105 ][ 193 ],
   alphaCSR[ 105 ][ 194 ],
   alphaCSR[ 105 ][ 195 ],
   alphaCSR[ 105 ][ 196 ],
   alphaCSR[ 105 ][ 197 ],
   alphaCSR[ 105 ][ 198 ],
   alphaCSR[ 105 ][ 199 ],
   alphaCSR[ 105 ][ 200 ],
   alphaCSR[ 105 ][ 201 ],
   alphaCSR[ 105 ][ 202 ],
   alphaCSR[ 105 ][ 203 ],
   alphaCSR[ 105 ][ 204 ],
   alphaCSR[ 105 ][ 205 ],
   alphaCSR[ 105 ][ 206 ],
   alphaCSR[ 105 ][ 207 ],
   alphaCSR[ 105 ][ 208 ],
   alphaCSR[ 105 ][ 209 ],
   alphaCSR[ 105 ][ 210 ],
   alphaCSR[ 105 ][ 211 ],
   alphaCSR[ 105 ][ 212 ],
   alphaCSR[ 105 ][ 213 ],
   alphaCSR[ 105 ][ 214 ],
   alphaCSR[ 105 ][ 215 ],
   alphaCSR[ 105 ][ 216 ],
   alphaCSR[ 105 ][ 217 ],
   alphaCSR[ 105 ][ 218 ],
   alphaCSR[ 105 ][ 219 ],
   alphaCSR[ 105 ][ 220 ],
   alphaCSR[ 105 ][ 221 ],
   alphaCSR[ 105 ][ 222 ],
   alphaCSR[ 105 ][ 223 ],
   alphaCSR[ 105 ][ 224 ],
   alphaCSR[ 105 ][ 225 ],
   alphaCSR[ 105 ][ 226 ],
   alphaCSR[ 105 ][ 227 ],
   alphaCSR[ 105 ][ 228 ],
   alphaCSR[ 105 ][ 229 ],
   alphaCSR[ 105 ][ 230 ],
   alphaCSR[ 105 ][ 231 ],
   alphaCSR[ 105 ][ 232 ],
   alphaCSR[ 105 ][ 233 ],
   alphaCSR[ 105 ][ 234 ],
   alphaCSR[ 105 ][ 235 ],
   alphaCSR[ 105 ][ 236 ],
   alphaCSR[ 105 ][ 237 ],
   alphaCSR[ 105 ][ 238 ],
   alphaCSR[ 105 ][ 239 ],
   alphaCSR[ 105 ][ 240 ],
   alphaCSR[ 105 ][ 241 ],
   alphaCSR[ 105 ][ 242 ],
   alphaCSR[ 105 ][ 243 ],
   alphaCSR[ 105 ][ 244 ],
   alphaCSR[ 105 ][ 245 ],
   alphaCSR[ 105 ][ 246 ],
   alphaCSR[ 105 ][ 247 ],
   alphaCSR[ 105 ][ 248 ],
   alphaCSR[ 105 ][ 249 ],
   alphaCSR[ 105 ][ 250 ],
   alphaCSR[ 105 ][ 251 ],
   alphaCSR[ 105 ][ 252 ],
   alphaCSR[ 105 ][ 253 ],
   alphaCSR[ 105 ][ 254 ],
   alphaCSR[ 105 ][ 255 ],
   alphaCSR[ 105 ][ 256 ],
   alphaCSR[ 105 ][ 257 ],
   alphaCSR[ 105 ][ 258 ],
   alphaCSR[ 105 ][ 259 ],
   alphaCSR[ 105 ][ 260 ],
   alphaCSR[ 105 ][ 261 ],
   alphaCSR[ 105 ][ 262 ],
   alphaCSR[ 105 ][ 263 ],
   alphaCSR[ 105 ][ 264 ],
   alphaCSR[ 105 ][ 265 ],
   alphaCSR[ 105 ][ 266 ],
   alphaCSR[ 105 ][ 267 ],
   alphaCSR[ 105 ][ 268 ],
   alphaCSR[ 105 ][ 269 ],
   alphaCSR[ 105 ][ 270 ],
   alphaCSR[ 105 ][ 271 ],
   alphaCSR[ 105 ][ 272 ],
   alphaCSR[ 105 ][ 273 ],
   alphaCSR[ 105 ][ 274 ],
   alphaCSR[ 105 ][ 275 ],
   alphaCSR[ 105 ][ 276 ],
   alphaCSR[ 105 ][ 277 ],
   alphaCSR[ 105 ][ 278 ],
   alphaCSR[ 105 ][ 279 ],
   alphaCSR[ 105 ][ 280 ],
   alphaCSR[ 105 ][ 281 ],
   alphaCSR[ 105 ][ 282 ],
   alphaCSR[ 105 ][ 283 ],
   alphaCSR[ 105 ][ 284 ],
   alphaCSR[ 105 ][ 285 ],
   alphaCSR[ 105 ][ 286 ],
   alphaCSR[ 105 ][ 287 ],
   alphaCSR[ 105 ][ 288 ],
   alphaCSR[ 105 ][ 289 ],
   alphaCSR[ 105 ][ 290 ],
   alphaCSR[ 105 ][ 291 ],
   alphaCSR[ 105 ][ 292 ],
   alphaCSR[ 105 ][ 293 ],
   alphaCSR[ 105 ][ 294 ],
   alphaCSR[ 105 ][ 295 ],
   alphaCSR[ 105 ][ 296 ],
   alphaCSR[ 105 ][ 297 ],
   alphaCSR[ 105 ][ 298 ],
   alphaCSR[ 105 ][ 299 ],
   alphaCSR[ 105 ][ 300 ],
   alphaCSR[ 105 ][ 301 ],
   alphaCSR[ 105 ][ 302 ],
   alphaCSR[ 105 ][ 303 ],
   alphaCSR[ 105 ][ 304 ],
   alphaCSR[ 105 ][ 305 ],
   alphaCSR[ 105 ][ 306 ],
   alphaCSR[ 105 ][ 307 ],
   alphaCSR[ 105 ][ 308 ],
   alphaCSR[ 105 ][ 309 ],
   alphaCSR[ 105 ][ 310 ],
   alphaCSR[ 105 ][ 311 ],
   alphaCSR[ 105 ][ 312 ],
   alphaCSR[ 105 ][ 313 ],
   alphaCSR[ 105 ][ 314 ],
   alphaCSR[ 105 ][ 315 ],
   alphaCSR[ 105 ][ 316 ],
   alphaCSR[ 105 ][ 317 ],
   alphaCSR[ 105 ][ 318 ],
   alphaCSR[ 105 ][ 319 ],
   alphaCSR[ 105 ][ 320 ],
   alphaCSR[ 105 ][ 321 ],
   alphaCSR[ 105 ][ 322 ],
   alphaCSR[ 105 ][ 323 ],
   alphaCSR[ 105 ][ 324 ],
   alphaCSR[ 105 ][ 325 ],
   alphaCSR[ 105 ][ 326 ],
   alphaCSR[ 105 ][ 327 ],
   alphaCSR[ 105 ][ 328 ],
   alphaCSR[ 105 ][ 329 ],
   alphaCSR[ 105 ][ 330 ],
   alphaCSR[ 105 ][ 331 ],
   alphaCSR[ 105 ][ 332 ],
   alphaCSR[ 105 ][ 333 ],
   alphaCSR[ 105 ][ 334 ],
   alphaCSR[ 105 ][ 335 ],
   alphaCSR[ 105 ][ 336 ],
   alphaCSR[ 105 ][ 337 ],
   alphaCSR[ 105 ][ 338 ],
   alphaCSR[ 105 ][ 339 ],
   alphaCSR[ 105 ][ 340 ],
   alphaCSR[ 105 ][ 341 ],
   alphaCSR[ 105 ][ 342 ],
   alphaCSR[ 105 ][ 343 ],
   alphaCSR[ 105 ][ 344 ],
   alphaCSR[ 105 ][ 345 ],
   alphaCSR[ 105 ][ 346 ],
   alphaCSR[ 105 ][ 347 ],
   alphaCSR[ 105 ][ 348 ],
   alphaCSR[ 105 ][ 349 ],
   alphaCSR[ 105 ][ 350 ],
   alphaCSR[ 105 ][ 351 ],
   alphaCSR[ 105 ][ 352 ],
   alphaCSR[ 105 ][ 353 ],
   alphaCSR[ 105 ][ 354 ],
   alphaCSR[ 105 ][ 355 ],
   alphaCSR[ 105 ][ 356 ],
   alphaCSR[ 105 ][ 357 ],
   alphaCSR[ 105 ][ 358 ],
   alphaCSR[ 105 ][ 359 ],
   alphaCSR[ 105 ][ 360 ],
   alphaCSR[ 105 ][ 361 ],
   alphaCSR[ 105 ][ 362 ],
   alphaCSR[ 105 ][ 363 ],
   alphaCSR[ 105 ][ 364 ],
   alphaCSR[ 105 ][ 365 ],
   alphaCSR[ 105 ][ 366 ],
   alphaCSR[ 105 ][ 367 ],
   alphaCSR[ 105 ][ 368 ],
   alphaCSR[ 105 ][ 369 ],
   alphaCSR[ 105 ][ 370 ],
   alphaCSR[ 105 ][ 371 ],
   alphaCSR[ 105 ][ 372 ],
   alphaCSR[ 105 ][ 373 ],
   alphaCSR[ 105 ][ 374 ],
   alphaCSR[ 105 ][ 375 ],
   alphaCSR[ 105 ][ 376 ],
   alphaCSR[ 105 ][ 377 ],
   alphaCSR[ 105 ][ 378 ],
   alphaCSR[ 105 ][ 379 ],
   alphaCSR[ 105 ][ 380 ],
   alphaCSR[ 105 ][ 381 ],
   alphaCSR[ 105 ][ 382 ],
   alphaCSR[ 105 ][ 383 ],
   alphaCSR[ 106 ][ 0 ],
   alphaCSR[ 106 ][ 1 ],
   alphaCSR[ 106 ][ 2 ],
   alphaCSR[ 106 ][ 3 ],
   alphaCSR[ 106 ][ 4 ],
   alphaCSR[ 106 ][ 5 ],
   alphaCSR[ 106 ][ 6 ],
   alphaCSR[ 106 ][ 7 ],
   alphaCSR[ 106 ][ 8 ],
   alphaCSR[ 106 ][ 9 ],
   alphaCSR[ 106 ][ 10 ],
   alphaCSR[ 106 ][ 11 ],
   alphaCSR[ 106 ][ 12 ],
   alphaCSR[ 106 ][ 13 ],
   alphaCSR[ 106 ][ 14 ],
   alphaCSR[ 106 ][ 15 ],
   alphaCSR[ 106 ][ 16 ],
   alphaCSR[ 106 ][ 17 ],
   alphaCSR[ 106 ][ 18 ],
   alphaCSR[ 106 ][ 19 ],
   alphaCSR[ 106 ][ 20 ],
   alphaCSR[ 106 ][ 21 ],
   alphaCSR[ 106 ][ 22 ],
   alphaCSR[ 106 ][ 23 ],
   alphaCSR[ 106 ][ 24 ],
   alphaCSR[ 106 ][ 25 ],
   alphaCSR[ 106 ][ 26 ],
   alphaCSR[ 106 ][ 27 ],
   alphaCSR[ 106 ][ 28 ],
   alphaCSR[ 106 ][ 29 ],
   alphaCSR[ 106 ][ 30 ],
   alphaCSR[ 106 ][ 31 ],
   alphaCSR[ 106 ][ 32 ],
   alphaCSR[ 106 ][ 33 ],
   alphaCSR[ 106 ][ 34 ],
   alphaCSR[ 106 ][ 35 ],
   alphaCSR[ 106 ][ 36 ],
   alphaCSR[ 106 ][ 37 ],
   alphaCSR[ 106 ][ 38 ],
   alphaCSR[ 106 ][ 39 ],
   alphaCSR[ 106 ][ 40 ],
   alphaCSR[ 106 ][ 41 ],
   alphaCSR[ 106 ][ 42 ],
   alphaCSR[ 106 ][ 43 ],
   alphaCSR[ 106 ][ 44 ],
   alphaCSR[ 106 ][ 45 ],
   alphaCSR[ 106 ][ 46 ],
   alphaCSR[ 106 ][ 47 ],
   alphaCSR[ 106 ][ 48 ],
   alphaCSR[ 106 ][ 49 ],
   alphaCSR[ 106 ][ 50 ],
   alphaCSR[ 106 ][ 51 ],
   alphaCSR[ 106 ][ 52 ],
   alphaCSR[ 106 ][ 53 ],
   alphaCSR[ 106 ][ 54 ],
   alphaCSR[ 106 ][ 55 ],
   alphaCSR[ 106 ][ 56 ],
   alphaCSR[ 106 ][ 57 ],
   alphaCSR[ 106 ][ 58 ],
   alphaCSR[ 106 ][ 59 ],
   alphaCSR[ 106 ][ 60 ],
   alphaCSR[ 106 ][ 61 ],
   alphaCSR[ 106 ][ 62 ],
   alphaCSR[ 106 ][ 63 ],
   alphaCSR[ 106 ][ 64 ],
   alphaCSR[ 106 ][ 65 ],
   alphaCSR[ 106 ][ 66 ],
   alphaCSR[ 106 ][ 67 ],
   alphaCSR[ 106 ][ 68 ],
   alphaCSR[ 106 ][ 69 ],
   alphaCSR[ 106 ][ 70 ],
   alphaCSR[ 106 ][ 71 ],
   alphaCSR[ 106 ][ 72 ],
   alphaCSR[ 106 ][ 73 ],
   alphaCSR[ 106 ][ 74 ],
   alphaCSR[ 106 ][ 75 ],
   alphaCSR[ 106 ][ 76 ],
   alphaCSR[ 106 ][ 77 ],
   alphaCSR[ 106 ][ 78 ],
   alphaCSR[ 106 ][ 79 ],
   alphaCSR[ 106 ][ 80 ],
   alphaCSR[ 106 ][ 81 ],
   alphaCSR[ 106 ][ 82 ],
   alphaCSR[ 106 ][ 83 ],
   alphaCSR[ 106 ][ 84 ],
   alphaCSR[ 106 ][ 85 ],
   alphaCSR[ 106 ][ 86 ],
   alphaCSR[ 106 ][ 87 ],
   alphaCSR[ 106 ][ 88 ],
   alphaCSR[ 106 ][ 89 ],
   alphaCSR[ 106 ][ 90 ],
   alphaCSR[ 106 ][ 91 ],
   alphaCSR[ 106 ][ 92 ],
   alphaCSR[ 106 ][ 93 ],
   alphaCSR[ 106 ][ 94 ],
   alphaCSR[ 106 ][ 95 ],
   alphaCSR[ 106 ][ 96 ],
   alphaCSR[ 106 ][ 97 ],
   alphaCSR[ 106 ][ 98 ],
   alphaCSR[ 106 ][ 99 ],
   alphaCSR[ 106 ][ 100 ],
   alphaCSR[ 106 ][ 101 ],
   alphaCSR[ 106 ][ 102 ],
   alphaCSR[ 106 ][ 103 ],
   alphaCSR[ 106 ][ 104 ],
   alphaCSR[ 106 ][ 105 ],
   alphaCSR[ 106 ][ 106 ],
   alphaCSR[ 106 ][ 107 ],
   alphaCSR[ 106 ][ 108 ],
   alphaCSR[ 106 ][ 109 ],
   alphaCSR[ 106 ][ 110 ],
   alphaCSR[ 106 ][ 111 ],
   alphaCSR[ 106 ][ 112 ],
   alphaCSR[ 106 ][ 113 ],
   alphaCSR[ 106 ][ 114 ],
   alphaCSR[ 106 ][ 115 ],
   alphaCSR[ 106 ][ 116 ],
   alphaCSR[ 106 ][ 117 ],
   alphaCSR[ 106 ][ 118 ],
   alphaCSR[ 106 ][ 119 ],
   alphaCSR[ 106 ][ 120 ],
   alphaCSR[ 106 ][ 121 ],
   alphaCSR[ 106 ][ 122 ],
   alphaCSR[ 106 ][ 123 ],
   alphaCSR[ 106 ][ 124 ],
   alphaCSR[ 106 ][ 125 ],
   alphaCSR[ 106 ][ 126 ],
   alphaCSR[ 106 ][ 127 ],
   alphaCSR[ 106 ][ 128 ],
   alphaCSR[ 106 ][ 129 ],
   alphaCSR[ 106 ][ 130 ],
   alphaCSR[ 106 ][ 131 ],
   alphaCSR[ 106 ][ 132 ],
   alphaCSR[ 106 ][ 133 ],
   alphaCSR[ 106 ][ 134 ],
   alphaCSR[ 106 ][ 135 ],
   alphaCSR[ 106 ][ 136 ],
   alphaCSR[ 106 ][ 137 ],
   alphaCSR[ 106 ][ 138 ],
   alphaCSR[ 106 ][ 139 ],
   alphaCSR[ 106 ][ 140 ],
   alphaCSR[ 106 ][ 141 ],
   alphaCSR[ 106 ][ 142 ],
   alphaCSR[ 106 ][ 143 ],
   alphaCSR[ 106 ][ 144 ],
   alphaCSR[ 106 ][ 145 ],
   alphaCSR[ 106 ][ 146 ],
   alphaCSR[ 106 ][ 147 ],
   alphaCSR[ 106 ][ 148 ],
   alphaCSR[ 106 ][ 149 ],
   alphaCSR[ 106 ][ 150 ],
   alphaCSR[ 106 ][ 151 ],
   alphaCSR[ 106 ][ 152 ],
   alphaCSR[ 106 ][ 153 ],
   alphaCSR[ 106 ][ 154 ],
   alphaCSR[ 106 ][ 155 ],
   alphaCSR[ 106 ][ 156 ],
   alphaCSR[ 106 ][ 157 ],
   alphaCSR[ 106 ][ 158 ],
   alphaCSR[ 106 ][ 159 ],
   alphaCSR[ 106 ][ 160 ],
   alphaCSR[ 106 ][ 161 ],
   alphaCSR[ 106 ][ 162 ],
   alphaCSR[ 106 ][ 163 ],
   alphaCSR[ 106 ][ 164 ],
   alphaCSR[ 106 ][ 165 ],
   alphaCSR[ 106 ][ 166 ],
   alphaCSR[ 106 ][ 167 ],
   alphaCSR[ 106 ][ 168 ],
   alphaCSR[ 106 ][ 169 ],
   alphaCSR[ 106 ][ 170 ],
   alphaCSR[ 106 ][ 171 ],
   alphaCSR[ 106 ][ 172 ],
   alphaCSR[ 106 ][ 173 ],
   alphaCSR[ 106 ][ 174 ],
   alphaCSR[ 106 ][ 175 ],
   alphaCSR[ 106 ][ 176 ],
   alphaCSR[ 106 ][ 177 ],
   alphaCSR[ 106 ][ 178 ],
   alphaCSR[ 106 ][ 179 ],
   alphaCSR[ 106 ][ 180 ],
   alphaCSR[ 106 ][ 181 ],
   alphaCSR[ 106 ][ 182 ],
   alphaCSR[ 106 ][ 183 ],
   alphaCSR[ 106 ][ 184 ],
   alphaCSR[ 106 ][ 185 ],
   alphaCSR[ 106 ][ 186 ],
   alphaCSR[ 106 ][ 187 ],
   alphaCSR[ 106 ][ 188 ],
   alphaCSR[ 106 ][ 189 ],
   alphaCSR[ 106 ][ 190 ],
   alphaCSR[ 106 ][ 191 ],
   alphaCSR[ 106 ][ 192 ],
   alphaCSR[ 106 ][ 193 ],
   alphaCSR[ 106 ][ 194 ],
   alphaCSR[ 106 ][ 195 ],
   alphaCSR[ 106 ][ 196 ],
   alphaCSR[ 106 ][ 197 ],
   alphaCSR[ 106 ][ 198 ],
   alphaCSR[ 106 ][ 199 ],
   alphaCSR[ 106 ][ 200 ],
   alphaCSR[ 106 ][ 201 ],
   alphaCSR[ 106 ][ 202 ],
   alphaCSR[ 106 ][ 203 ],
   alphaCSR[ 106 ][ 204 ],
   alphaCSR[ 106 ][ 205 ],
   alphaCSR[ 106 ][ 206 ],
   alphaCSR[ 106 ][ 207 ],
   alphaCSR[ 106 ][ 208 ],
   alphaCSR[ 106 ][ 209 ],
   alphaCSR[ 106 ][ 210 ],
   alphaCSR[ 106 ][ 211 ],
   alphaCSR[ 106 ][ 212 ],
   alphaCSR[ 106 ][ 213 ],
   alphaCSR[ 106 ][ 214 ],
   alphaCSR[ 106 ][ 215 ],
   alphaCSR[ 106 ][ 216 ],
   alphaCSR[ 106 ][ 217 ],
   alphaCSR[ 106 ][ 218 ],
   alphaCSR[ 106 ][ 219 ],
   alphaCSR[ 106 ][ 220 ],
   alphaCSR[ 106 ][ 221 ],
   alphaCSR[ 106 ][ 222 ],
   alphaCSR[ 106 ][ 223 ],
   alphaCSR[ 106 ][ 224 ],
   alphaCSR[ 106 ][ 225 ],
   alphaCSR[ 106 ][ 226 ],
   alphaCSR[ 106 ][ 227 ],
   alphaCSR[ 106 ][ 228 ],
   alphaCSR[ 106 ][ 229 ],
   alphaCSR[ 106 ][ 230 ],
   alphaCSR[ 106 ][ 231 ],
   alphaCSR[ 106 ][ 232 ],
   alphaCSR[ 106 ][ 233 ],
   alphaCSR[ 106 ][ 234 ],
   alphaCSR[ 106 ][ 235 ],
   alphaCSR[ 106 ][ 236 ],
   alphaCSR[ 106 ][ 237 ],
   alphaCSR[ 106 ][ 238 ],
   alphaCSR[ 106 ][ 239 ],
   alphaCSR[ 106 ][ 240 ],
   alphaCSR[ 106 ][ 241 ],
   alphaCSR[ 106 ][ 242 ],
   alphaCSR[ 106 ][ 243 ],
   alphaCSR[ 106 ][ 244 ],
   alphaCSR[ 106 ][ 245 ],
   alphaCSR[ 106 ][ 246 ],
   alphaCSR[ 106 ][ 247 ],
   alphaCSR[ 106 ][ 248 ],
   alphaCSR[ 106 ][ 249 ],
   alphaCSR[ 106 ][ 250 ],
   alphaCSR[ 106 ][ 251 ],
   alphaCSR[ 106 ][ 252 ],
   alphaCSR[ 106 ][ 253 ],
   alphaCSR[ 106 ][ 254 ],
   alphaCSR[ 106 ][ 255 ],
   alphaCSR[ 106 ][ 256 ],
   alphaCSR[ 106 ][ 257 ],
   alphaCSR[ 106 ][ 258 ],
   alphaCSR[ 106 ][ 259 ],
   alphaCSR[ 106 ][ 260 ],
   alphaCSR[ 106 ][ 261 ],
   alphaCSR[ 106 ][ 262 ],
   alphaCSR[ 106 ][ 263 ],
   alphaCSR[ 106 ][ 264 ],
   alphaCSR[ 106 ][ 265 ],
   alphaCSR[ 106 ][ 266 ],
   alphaCSR[ 106 ][ 267 ],
   alphaCSR[ 106 ][ 268 ],
   alphaCSR[ 106 ][ 269 ],
   alphaCSR[ 106 ][ 270 ],
   alphaCSR[ 106 ][ 271 ],
   alphaCSR[ 106 ][ 272 ],
   alphaCSR[ 106 ][ 273 ],
   alphaCSR[ 106 ][ 274 ],
   alphaCSR[ 106 ][ 275 ],
   alphaCSR[ 106 ][ 276 ],
   alphaCSR[ 106 ][ 277 ],
   alphaCSR[ 106 ][ 278 ],
   alphaCSR[ 106 ][ 279 ],
   alphaCSR[ 106 ][ 280 ],
   alphaCSR[ 106 ][ 281 ],
   alphaCSR[ 106 ][ 282 ],
   alphaCSR[ 106 ][ 283 ],
   alphaCSR[ 106 ][ 284 ],
   alphaCSR[ 106 ][ 285 ],
   alphaCSR[ 106 ][ 286 ],
   alphaCSR[ 106 ][ 287 ],
   alphaCSR[ 106 ][ 288 ],
   alphaCSR[ 106 ][ 289 ],
   alphaCSR[ 106 ][ 290 ],
   alphaCSR[ 106 ][ 291 ],
   alphaCSR[ 106 ][ 292 ],
   alphaCSR[ 106 ][ 293 ],
   alphaCSR[ 106 ][ 294 ],
   alphaCSR[ 106 ][ 295 ],
   alphaCSR[ 106 ][ 296 ],
   alphaCSR[ 106 ][ 297 ],
   alphaCSR[ 106 ][ 298 ],
   alphaCSR[ 106 ][ 299 ],
   alphaCSR[ 106 ][ 300 ],
   alphaCSR[ 106 ][ 301 ],
   alphaCSR[ 106 ][ 302 ],
   alphaCSR[ 106 ][ 303 ],
   alphaCSR[ 106 ][ 304 ],
   alphaCSR[ 106 ][ 305 ],
   alphaCSR[ 106 ][ 306 ],
   alphaCSR[ 106 ][ 307 ],
   alphaCSR[ 106 ][ 308 ],
   alphaCSR[ 106 ][ 309 ],
   alphaCSR[ 106 ][ 310 ],
   alphaCSR[ 106 ][ 311 ],
   alphaCSR[ 106 ][ 312 ],
   alphaCSR[ 106 ][ 313 ],
   alphaCSR[ 106 ][ 314 ],
   alphaCSR[ 106 ][ 315 ],
   alphaCSR[ 106 ][ 316 ],
   alphaCSR[ 106 ][ 317 ],
   alphaCSR[ 106 ][ 318 ],
   alphaCSR[ 106 ][ 319 ],
   alphaCSR[ 106 ][ 320 ],
   alphaCSR[ 106 ][ 321 ],
   alphaCSR[ 106 ][ 322 ],
   alphaCSR[ 106 ][ 323 ],
   alphaCSR[ 106 ][ 324 ],
   alphaCSR[ 106 ][ 325 ],
   alphaCSR[ 106 ][ 326 ],
   alphaCSR[ 106 ][ 327 ],
   alphaCSR[ 106 ][ 328 ],
   alphaCSR[ 106 ][ 329 ],
   alphaCSR[ 106 ][ 330 ],
   alphaCSR[ 106 ][ 331 ],
   alphaCSR[ 106 ][ 332 ],
   alphaCSR[ 106 ][ 333 ],
   alphaCSR[ 106 ][ 334 ],
   alphaCSR[ 106 ][ 335 ],
   alphaCSR[ 106 ][ 336 ],
   alphaCSR[ 106 ][ 337 ],
   alphaCSR[ 106 ][ 338 ],
   alphaCSR[ 106 ][ 339 ],
   alphaCSR[ 106 ][ 340 ],
   alphaCSR[ 106 ][ 341 ],
   alphaCSR[ 106 ][ 342 ],
   alphaCSR[ 106 ][ 343 ],
   alphaCSR[ 106 ][ 344 ],
   alphaCSR[ 106 ][ 345 ],
   alphaCSR[ 106 ][ 346 ],
   alphaCSR[ 106 ][ 347 ],
   alphaCSR[ 106 ][ 348 ],
   alphaCSR[ 106 ][ 349 ],
   alphaCSR[ 106 ][ 350 ],
   alphaCSR[ 106 ][ 351 ],
   alphaCSR[ 106 ][ 352 ],
   alphaCSR[ 106 ][ 353 ],
   alphaCSR[ 106 ][ 354 ],
   alphaCSR[ 106 ][ 355 ],
   alphaCSR[ 106 ][ 356 ],
   alphaCSR[ 106 ][ 357 ],
   alphaCSR[ 106 ][ 358 ],
   alphaCSR[ 106 ][ 359 ],
   alphaCSR[ 106 ][ 360 ],
   alphaCSR[ 106 ][ 361 ],
   alphaCSR[ 106 ][ 362 ],
   alphaCSR[ 106 ][ 363 ],
   alphaCSR[ 106 ][ 364 ],
   alphaCSR[ 106 ][ 365 ],
   alphaCSR[ 106 ][ 366 ],
   alphaCSR[ 106 ][ 367 ],
   alphaCSR[ 106 ][ 368 ],
   alphaCSR[ 106 ][ 369 ],
   alphaCSR[ 106 ][ 370 ],
   alphaCSR[ 106 ][ 371 ],
   alphaCSR[ 106 ][ 372 ],
   alphaCSR[ 106 ][ 373 ],
   alphaCSR[ 106 ][ 374 ],
   alphaCSR[ 106 ][ 375 ],
   alphaCSR[ 106 ][ 376 ],
   alphaCSR[ 106 ][ 377 ],
   alphaCSR[ 106 ][ 378 ],
   alphaCSR[ 106 ][ 379 ],
   alphaCSR[ 106 ][ 380 ],
   alphaCSR[ 106 ][ 381 ],
   alphaCSR[ 106 ][ 382 ],
   alphaCSR[ 106 ][ 383 ],
   alphaCSR[ 107 ][ 0 ],
   alphaCSR[ 107 ][ 1 ],
   alphaCSR[ 107 ][ 2 ],
   alphaCSR[ 107 ][ 3 ],
   alphaCSR[ 107 ][ 4 ],
   alphaCSR[ 107 ][ 5 ],
   alphaCSR[ 107 ][ 6 ],
   alphaCSR[ 107 ][ 7 ],
   alphaCSR[ 107 ][ 8 ],
   alphaCSR[ 107 ][ 9 ],
   alphaCSR[ 107 ][ 10 ],
   alphaCSR[ 107 ][ 11 ],
   alphaCSR[ 107 ][ 12 ],
   alphaCSR[ 107 ][ 13 ],
   alphaCSR[ 107 ][ 14 ],
   alphaCSR[ 107 ][ 15 ],
   alphaCSR[ 107 ][ 16 ],
   alphaCSR[ 107 ][ 17 ],
   alphaCSR[ 107 ][ 18 ],
   alphaCSR[ 107 ][ 19 ],
   alphaCSR[ 107 ][ 20 ],
   alphaCSR[ 107 ][ 21 ],
   alphaCSR[ 107 ][ 22 ],
   alphaCSR[ 107 ][ 23 ],
   alphaCSR[ 107 ][ 24 ],
   alphaCSR[ 107 ][ 25 ],
   alphaCSR[ 107 ][ 26 ],
   alphaCSR[ 107 ][ 27 ],
   alphaCSR[ 107 ][ 28 ],
   alphaCSR[ 107 ][ 29 ],
   alphaCSR[ 107 ][ 30 ],
   alphaCSR[ 107 ][ 31 ],
   alphaCSR[ 107 ][ 32 ],
   alphaCSR[ 107 ][ 33 ],
   alphaCSR[ 107 ][ 34 ],
   alphaCSR[ 107 ][ 35 ],
   alphaCSR[ 107 ][ 36 ],
   alphaCSR[ 107 ][ 37 ],
   alphaCSR[ 107 ][ 38 ],
   alphaCSR[ 107 ][ 39 ],
   alphaCSR[ 107 ][ 40 ],
   alphaCSR[ 107 ][ 41 ],
   alphaCSR[ 107 ][ 42 ],
   alphaCSR[ 107 ][ 43 ],
   alphaCSR[ 107 ][ 44 ],
   alphaCSR[ 107 ][ 45 ],
   alphaCSR[ 107 ][ 46 ],
   alphaCSR[ 107 ][ 47 ],
   alphaCSR[ 107 ][ 48 ],
   alphaCSR[ 107 ][ 49 ],
   alphaCSR[ 107 ][ 50 ],
   alphaCSR[ 107 ][ 51 ],
   alphaCSR[ 107 ][ 52 ],
   alphaCSR[ 107 ][ 53 ],
   alphaCSR[ 107 ][ 54 ],
   alphaCSR[ 107 ][ 55 ],
   alphaCSR[ 107 ][ 56 ],
   alphaCSR[ 107 ][ 57 ],
   alphaCSR[ 107 ][ 58 ],
   alphaCSR[ 107 ][ 59 ],
   alphaCSR[ 107 ][ 60 ],
   alphaCSR[ 107 ][ 61 ],
   alphaCSR[ 107 ][ 62 ],
   alphaCSR[ 107 ][ 63 ],
   alphaCSR[ 107 ][ 64 ],
   alphaCSR[ 107 ][ 65 ],
   alphaCSR[ 107 ][ 66 ],
   alphaCSR[ 107 ][ 67 ],
   alphaCSR[ 107 ][ 68 ],
   alphaCSR[ 107 ][ 69 ],
   alphaCSR[ 107 ][ 70 ],
   alphaCSR[ 107 ][ 71 ],
   alphaCSR[ 107 ][ 72 ],
   alphaCSR[ 107 ][ 73 ],
   alphaCSR[ 107 ][ 74 ],
   alphaCSR[ 107 ][ 75 ],
   alphaCSR[ 107 ][ 76 ],
   alphaCSR[ 107 ][ 77 ],
   alphaCSR[ 107 ][ 78 ],
   alphaCSR[ 107 ][ 79 ],
   alphaCSR[ 107 ][ 80 ],
   alphaCSR[ 107 ][ 81 ],
   alphaCSR[ 107 ][ 82 ],
   alphaCSR[ 107 ][ 83 ],
   alphaCSR[ 107 ][ 84 ],
   alphaCSR[ 107 ][ 85 ],
   alphaCSR[ 107 ][ 86 ],
   alphaCSR[ 107 ][ 87 ],
   alphaCSR[ 107 ][ 88 ],
   alphaCSR[ 107 ][ 89 ],
   alphaCSR[ 107 ][ 90 ],
   alphaCSR[ 107 ][ 91 ],
   alphaCSR[ 107 ][ 92 ],
   alphaCSR[ 107 ][ 93 ],
   alphaCSR[ 107 ][ 94 ],
   alphaCSR[ 107 ][ 95 ],
   alphaCSR[ 107 ][ 96 ],
   alphaCSR[ 107 ][ 97 ],
   alphaCSR[ 107 ][ 98 ],
   alphaCSR[ 107 ][ 99 ],
   alphaCSR[ 107 ][ 100 ],
   alphaCSR[ 107 ][ 101 ],
   alphaCSR[ 107 ][ 102 ],
   alphaCSR[ 107 ][ 103 ],
   alphaCSR[ 107 ][ 104 ],
   alphaCSR[ 107 ][ 105 ],
   alphaCSR[ 107 ][ 106 ],
   alphaCSR[ 107 ][ 107 ],
   alphaCSR[ 107 ][ 108 ],
   alphaCSR[ 107 ][ 109 ],
   alphaCSR[ 107 ][ 110 ],
   alphaCSR[ 107 ][ 111 ],
   alphaCSR[ 107 ][ 112 ],
   alphaCSR[ 107 ][ 113 ],
   alphaCSR[ 107 ][ 114 ],
   alphaCSR[ 107 ][ 115 ],
   alphaCSR[ 107 ][ 116 ],
   alphaCSR[ 107 ][ 117 ],
   alphaCSR[ 107 ][ 118 ],
   alphaCSR[ 107 ][ 119 ],
   alphaCSR[ 107 ][ 120 ],
   alphaCSR[ 107 ][ 121 ],
   alphaCSR[ 107 ][ 122 ],
   alphaCSR[ 107 ][ 123 ],
   alphaCSR[ 107 ][ 124 ],
   alphaCSR[ 107 ][ 125 ],
   alphaCSR[ 107 ][ 126 ],
   alphaCSR[ 107 ][ 127 ],
   alphaCSR[ 107 ][ 128 ],
   alphaCSR[ 107 ][ 129 ],
   alphaCSR[ 107 ][ 130 ],
   alphaCSR[ 107 ][ 131 ],
   alphaCSR[ 107 ][ 132 ],
   alphaCSR[ 107 ][ 133 ],
   alphaCSR[ 107 ][ 134 ],
   alphaCSR[ 107 ][ 135 ],
   alphaCSR[ 107 ][ 136 ],
   alphaCSR[ 107 ][ 137 ],
   alphaCSR[ 107 ][ 138 ],
   alphaCSR[ 107 ][ 139 ],
   alphaCSR[ 107 ][ 140 ],
   alphaCSR[ 107 ][ 141 ],
   alphaCSR[ 107 ][ 142 ],
   alphaCSR[ 107 ][ 143 ],
   alphaCSR[ 107 ][ 144 ],
   alphaCSR[ 107 ][ 145 ],
   alphaCSR[ 107 ][ 146 ],
   alphaCSR[ 107 ][ 147 ],
   alphaCSR[ 107 ][ 148 ],
   alphaCSR[ 107 ][ 149 ],
   alphaCSR[ 107 ][ 150 ],
   alphaCSR[ 107 ][ 151 ],
   alphaCSR[ 107 ][ 152 ],
   alphaCSR[ 107 ][ 153 ],
   alphaCSR[ 107 ][ 154 ],
   alphaCSR[ 107 ][ 155 ],
   alphaCSR[ 107 ][ 156 ],
   alphaCSR[ 107 ][ 157 ],
   alphaCSR[ 107 ][ 158 ],
   alphaCSR[ 107 ][ 159 ],
   alphaCSR[ 107 ][ 160 ],
   alphaCSR[ 107 ][ 161 ],
   alphaCSR[ 107 ][ 162 ],
   alphaCSR[ 107 ][ 163 ],
   alphaCSR[ 107 ][ 164 ],
   alphaCSR[ 107 ][ 165 ],
   alphaCSR[ 107 ][ 166 ],
   alphaCSR[ 107 ][ 167 ],
   alphaCSR[ 107 ][ 168 ],
   alphaCSR[ 107 ][ 169 ],
   alphaCSR[ 107 ][ 170 ],
   alphaCSR[ 107 ][ 171 ],
   alphaCSR[ 107 ][ 172 ],
   alphaCSR[ 107 ][ 173 ],
   alphaCSR[ 107 ][ 174 ],
   alphaCSR[ 107 ][ 175 ],
   alphaCSR[ 107 ][ 176 ],
   alphaCSR[ 107 ][ 177 ],
   alphaCSR[ 107 ][ 178 ],
   alphaCSR[ 107 ][ 179 ],
   alphaCSR[ 107 ][ 180 ],
   alphaCSR[ 107 ][ 181 ],
   alphaCSR[ 107 ][ 182 ],
   alphaCSR[ 107 ][ 183 ],
   alphaCSR[ 107 ][ 184 ],
   alphaCSR[ 107 ][ 185 ],
   alphaCSR[ 107 ][ 186 ],
   alphaCSR[ 107 ][ 187 ],
   alphaCSR[ 107 ][ 188 ],
   alphaCSR[ 107 ][ 189 ],
   alphaCSR[ 107 ][ 190 ],
   alphaCSR[ 107 ][ 191 ],
   alphaCSR[ 107 ][ 192 ],
   alphaCSR[ 107 ][ 193 ],
   alphaCSR[ 107 ][ 194 ],
   alphaCSR[ 107 ][ 195 ],
   alphaCSR[ 107 ][ 196 ],
   alphaCSR[ 107 ][ 197 ],
   alphaCSR[ 107 ][ 198 ],
   alphaCSR[ 107 ][ 199 ],
   alphaCSR[ 107 ][ 200 ],
   alphaCSR[ 107 ][ 201 ],
   alphaCSR[ 107 ][ 202 ],
   alphaCSR[ 107 ][ 203 ],
   alphaCSR[ 107 ][ 204 ],
   alphaCSR[ 107 ][ 205 ],
   alphaCSR[ 107 ][ 206 ],
   alphaCSR[ 107 ][ 207 ],
   alphaCSR[ 107 ][ 208 ],
   alphaCSR[ 107 ][ 209 ],
   alphaCSR[ 107 ][ 210 ],
   alphaCSR[ 107 ][ 211 ],
   alphaCSR[ 107 ][ 212 ],
   alphaCSR[ 107 ][ 213 ],
   alphaCSR[ 107 ][ 214 ],
   alphaCSR[ 107 ][ 215 ],
   alphaCSR[ 107 ][ 216 ],
   alphaCSR[ 107 ][ 217 ],
   alphaCSR[ 107 ][ 218 ],
   alphaCSR[ 107 ][ 219 ],
   alphaCSR[ 107 ][ 220 ],
   alphaCSR[ 107 ][ 221 ],
   alphaCSR[ 107 ][ 222 ],
   alphaCSR[ 107 ][ 223 ],
   alphaCSR[ 107 ][ 224 ],
   alphaCSR[ 107 ][ 225 ],
   alphaCSR[ 107 ][ 226 ],
   alphaCSR[ 107 ][ 227 ],
   alphaCSR[ 107 ][ 228 ],
   alphaCSR[ 107 ][ 229 ],
   alphaCSR[ 107 ][ 230 ],
   alphaCSR[ 107 ][ 231 ],
   alphaCSR[ 107 ][ 232 ],
   alphaCSR[ 107 ][ 233 ],
   alphaCSR[ 107 ][ 234 ],
   alphaCSR[ 107 ][ 235 ],
   alphaCSR[ 107 ][ 236 ],
   alphaCSR[ 107 ][ 237 ],
   alphaCSR[ 107 ][ 238 ],
   alphaCSR[ 107 ][ 239 ],
   alphaCSR[ 107 ][ 240 ],
   alphaCSR[ 107 ][ 241 ],
   alphaCSR[ 107 ][ 242 ],
   alphaCSR[ 107 ][ 243 ],
   alphaCSR[ 107 ][ 244 ],
   alphaCSR[ 107 ][ 245 ],
   alphaCSR[ 107 ][ 246 ],
   alphaCSR[ 107 ][ 247 ],
   alphaCSR[ 107 ][ 248 ],
   alphaCSR[ 107 ][ 249 ],
   alphaCSR[ 107 ][ 250 ],
   alphaCSR[ 107 ][ 251 ],
   alphaCSR[ 107 ][ 252 ],
   alphaCSR[ 107 ][ 253 ],
   alphaCSR[ 107 ][ 254 ],
   alphaCSR[ 107 ][ 255 ],
   alphaCSR[ 107 ][ 256 ],
   alphaCSR[ 107 ][ 257 ],
   alphaCSR[ 107 ][ 258 ],
   alphaCSR[ 107 ][ 259 ],
   alphaCSR[ 107 ][ 260 ],
   alphaCSR[ 107 ][ 261 ],
   alphaCSR[ 107 ][ 262 ],
   alphaCSR[ 107 ][ 263 ],
   alphaCSR[ 107 ][ 264 ],
   alphaCSR[ 107 ][ 265 ],
   alphaCSR[ 107 ][ 266 ],
   alphaCSR[ 107 ][ 267 ],
   alphaCSR[ 107 ][ 268 ],
   alphaCSR[ 107 ][ 269 ],
   alphaCSR[ 107 ][ 270 ],
   alphaCSR[ 107 ][ 271 ],
   alphaCSR[ 107 ][ 272 ],
   alphaCSR[ 107 ][ 273 ],
   alphaCSR[ 107 ][ 274 ],
   alphaCSR[ 107 ][ 275 ],
   alphaCSR[ 107 ][ 276 ],
   alphaCSR[ 107 ][ 277 ],
   alphaCSR[ 107 ][ 278 ],
   alphaCSR[ 107 ][ 279 ],
   alphaCSR[ 107 ][ 280 ],
   alphaCSR[ 107 ][ 281 ],
   alphaCSR[ 107 ][ 282 ],
   alphaCSR[ 107 ][ 283 ],
   alphaCSR[ 107 ][ 284 ],
   alphaCSR[ 107 ][ 285 ],
   alphaCSR[ 107 ][ 286 ],
   alphaCSR[ 107 ][ 287 ],
   alphaCSR[ 107 ][ 288 ],
   alphaCSR[ 107 ][ 289 ],
   alphaCSR[ 107 ][ 290 ],
   alphaCSR[ 107 ][ 291 ],
   alphaCSR[ 107 ][ 292 ],
   alphaCSR[ 107 ][ 293 ],
   alphaCSR[ 107 ][ 294 ],
   alphaCSR[ 107 ][ 295 ],
   alphaCSR[ 107 ][ 296 ],
   alphaCSR[ 107 ][ 297 ],
   alphaCSR[ 107 ][ 298 ],
   alphaCSR[ 107 ][ 299 ],
   alphaCSR[ 107 ][ 300 ],
   alphaCSR[ 107 ][ 301 ],
   alphaCSR[ 107 ][ 302 ],
   alphaCSR[ 107 ][ 303 ],
   alphaCSR[ 107 ][ 304 ],
   alphaCSR[ 107 ][ 305 ],
   alphaCSR[ 107 ][ 306 ],
   alphaCSR[ 107 ][ 307 ],
   alphaCSR[ 107 ][ 308 ],
   alphaCSR[ 107 ][ 309 ],
   alphaCSR[ 107 ][ 310 ],
   alphaCSR[ 107 ][ 311 ],
   alphaCSR[ 107 ][ 312 ],
   alphaCSR[ 107 ][ 313 ],
   alphaCSR[ 107 ][ 314 ],
   alphaCSR[ 107 ][ 315 ],
   alphaCSR[ 107 ][ 316 ],
   alphaCSR[ 107 ][ 317 ],
   alphaCSR[ 107 ][ 318 ],
   alphaCSR[ 107 ][ 319 ],
   alphaCSR[ 107 ][ 320 ],
   alphaCSR[ 107 ][ 321 ],
   alphaCSR[ 107 ][ 322 ],
   alphaCSR[ 107 ][ 323 ],
   alphaCSR[ 107 ][ 324 ],
   alphaCSR[ 107 ][ 325 ],
   alphaCSR[ 107 ][ 326 ],
   alphaCSR[ 107 ][ 327 ],
   alphaCSR[ 107 ][ 328 ],
   alphaCSR[ 107 ][ 329 ],
   alphaCSR[ 107 ][ 330 ],
   alphaCSR[ 107 ][ 331 ],
   alphaCSR[ 107 ][ 332 ],
   alphaCSR[ 107 ][ 333 ],
   alphaCSR[ 107 ][ 334 ],
   alphaCSR[ 107 ][ 335 ],
   alphaCSR[ 107 ][ 336 ],
   alphaCSR[ 107 ][ 337 ],
   alphaCSR[ 107 ][ 338 ],
   alphaCSR[ 107 ][ 339 ],
   alphaCSR[ 107 ][ 340 ],
   alphaCSR[ 107 ][ 341 ],
   alphaCSR[ 107 ][ 342 ],
   alphaCSR[ 107 ][ 343 ],
   alphaCSR[ 107 ][ 344 ],
   alphaCSR[ 107 ][ 345 ],
   alphaCSR[ 107 ][ 346 ],
   alphaCSR[ 107 ][ 347 ],
   alphaCSR[ 107 ][ 348 ],
   alphaCSR[ 107 ][ 349 ],
   alphaCSR[ 107 ][ 350 ],
   alphaCSR[ 107 ][ 351 ],
   alphaCSR[ 107 ][ 352 ],
   alphaCSR[ 107 ][ 353 ],
   alphaCSR[ 107 ][ 354 ],
   alphaCSR[ 107 ][ 355 ],
   alphaCSR[ 107 ][ 356 ],
   alphaCSR[ 107 ][ 357 ],
   alphaCSR[ 107 ][ 358 ],
   alphaCSR[ 107 ][ 359 ],
   alphaCSR[ 107 ][ 360 ],
   alphaCSR[ 107 ][ 361 ],
   alphaCSR[ 107 ][ 362 ],
   alphaCSR[ 107 ][ 363 ],
   alphaCSR[ 107 ][ 364 ],
   alphaCSR[ 107 ][ 365 ],
   alphaCSR[ 107 ][ 366 ],
   alphaCSR[ 107 ][ 367 ],
   alphaCSR[ 107 ][ 368 ],
   alphaCSR[ 107 ][ 369 ],
   alphaCSR[ 107 ][ 370 ],
   alphaCSR[ 107 ][ 371 ],
   alphaCSR[ 107 ][ 372 ],
   alphaCSR[ 107 ][ 373 ],
   alphaCSR[ 107 ][ 374 ],
   alphaCSR[ 107 ][ 375 ],
   alphaCSR[ 107 ][ 376 ],
   alphaCSR[ 107 ][ 377 ],
   alphaCSR[ 107 ][ 378 ],
   alphaCSR[ 107 ][ 379 ],
   alphaCSR[ 107 ][ 380 ],
   alphaCSR[ 107 ][ 381 ],
   alphaCSR[ 107 ][ 382 ],
   alphaCSR[ 107 ][ 383 ],
   alphaCSR[ 108 ][ 0 ],
   alphaCSR[ 108 ][ 1 ],
   alphaCSR[ 108 ][ 2 ],
   alphaCSR[ 108 ][ 3 ],
   alphaCSR[ 108 ][ 4 ],
   alphaCSR[ 108 ][ 5 ],
   alphaCSR[ 108 ][ 6 ],
   alphaCSR[ 108 ][ 7 ],
   alphaCSR[ 108 ][ 8 ],
   alphaCSR[ 108 ][ 9 ],
   alphaCSR[ 108 ][ 10 ],
   alphaCSR[ 108 ][ 11 ],
   alphaCSR[ 108 ][ 12 ],
   alphaCSR[ 108 ][ 13 ],
   alphaCSR[ 108 ][ 14 ],
   alphaCSR[ 108 ][ 15 ],
   alphaCSR[ 108 ][ 16 ],
   alphaCSR[ 108 ][ 17 ],
   alphaCSR[ 108 ][ 18 ],
   alphaCSR[ 108 ][ 19 ],
   alphaCSR[ 108 ][ 20 ],
   alphaCSR[ 108 ][ 21 ],
   alphaCSR[ 108 ][ 22 ],
   alphaCSR[ 108 ][ 23 ],
   alphaCSR[ 108 ][ 24 ],
   alphaCSR[ 108 ][ 25 ],
   alphaCSR[ 108 ][ 26 ],
   alphaCSR[ 108 ][ 27 ],
   alphaCSR[ 108 ][ 28 ],
   alphaCSR[ 108 ][ 29 ],
   alphaCSR[ 108 ][ 30 ],
   alphaCSR[ 108 ][ 31 ],
   alphaCSR[ 108 ][ 32 ],
   alphaCSR[ 108 ][ 33 ],
   alphaCSR[ 108 ][ 34 ],
   alphaCSR[ 108 ][ 35 ],
   alphaCSR[ 108 ][ 36 ],
   alphaCSR[ 108 ][ 37 ],
   alphaCSR[ 108 ][ 38 ],
   alphaCSR[ 108 ][ 39 ],
   alphaCSR[ 108 ][ 40 ],
   alphaCSR[ 108 ][ 41 ],
   alphaCSR[ 108 ][ 42 ],
   alphaCSR[ 108 ][ 43 ],
   alphaCSR[ 108 ][ 44 ],
   alphaCSR[ 108 ][ 45 ],
   alphaCSR[ 108 ][ 46 ],
   alphaCSR[ 108 ][ 47 ],
   alphaCSR[ 108 ][ 48 ],
   alphaCSR[ 108 ][ 49 ],
   alphaCSR[ 108 ][ 50 ],
   alphaCSR[ 108 ][ 51 ],
   alphaCSR[ 108 ][ 52 ],
   alphaCSR[ 108 ][ 53 ],
   alphaCSR[ 108 ][ 54 ],
   alphaCSR[ 108 ][ 55 ],
   alphaCSR[ 108 ][ 56 ],
   alphaCSR[ 108 ][ 57 ],
   alphaCSR[ 108 ][ 58 ],
   alphaCSR[ 108 ][ 59 ],
   alphaCSR[ 108 ][ 60 ],
   alphaCSR[ 108 ][ 61 ],
   alphaCSR[ 108 ][ 62 ],
   alphaCSR[ 108 ][ 63 ],
   alphaCSR[ 108 ][ 64 ],
   alphaCSR[ 108 ][ 65 ],
   alphaCSR[ 108 ][ 66 ],
   alphaCSR[ 108 ][ 67 ],
   alphaCSR[ 108 ][ 68 ],
   alphaCSR[ 108 ][ 69 ],
   alphaCSR[ 108 ][ 70 ],
   alphaCSR[ 108 ][ 71 ],
   alphaCSR[ 108 ][ 72 ],
   alphaCSR[ 108 ][ 73 ],
   alphaCSR[ 108 ][ 74 ],
   alphaCSR[ 108 ][ 75 ],
   alphaCSR[ 108 ][ 76 ],
   alphaCSR[ 108 ][ 77 ],
   alphaCSR[ 108 ][ 78 ],
   alphaCSR[ 108 ][ 79 ],
   alphaCSR[ 108 ][ 80 ],
   alphaCSR[ 108 ][ 81 ],
   alphaCSR[ 108 ][ 82 ],
   alphaCSR[ 108 ][ 83 ],
   alphaCSR[ 108 ][ 84 ],
   alphaCSR[ 108 ][ 85 ],
   alphaCSR[ 108 ][ 86 ],
   alphaCSR[ 108 ][ 87 ],
   alphaCSR[ 108 ][ 88 ],
   alphaCSR[ 108 ][ 89 ],
   alphaCSR[ 108 ][ 90 ],
   alphaCSR[ 108 ][ 91 ],
   alphaCSR[ 108 ][ 92 ],
   alphaCSR[ 108 ][ 93 ],
   alphaCSR[ 108 ][ 94 ],
   alphaCSR[ 108 ][ 95 ],
   alphaCSR[ 108 ][ 96 ],
   alphaCSR[ 108 ][ 97 ],
   alphaCSR[ 108 ][ 98 ],
   alphaCSR[ 108 ][ 99 ],
   alphaCSR[ 108 ][ 100 ],
   alphaCSR[ 108 ][ 101 ],
   alphaCSR[ 108 ][ 102 ],
   alphaCSR[ 108 ][ 103 ],
   alphaCSR[ 108 ][ 104 ],
   alphaCSR[ 108 ][ 105 ],
   alphaCSR[ 108 ][ 106 ],
   alphaCSR[ 108 ][ 107 ],
   alphaCSR[ 108 ][ 108 ],
   alphaCSR[ 108 ][ 109 ],
   alphaCSR[ 108 ][ 110 ],
   alphaCSR[ 108 ][ 111 ],
   alphaCSR[ 108 ][ 112 ],
   alphaCSR[ 108 ][ 113 ],
   alphaCSR[ 108 ][ 114 ],
   alphaCSR[ 108 ][ 115 ],
   alphaCSR[ 108 ][ 116 ],
   alphaCSR[ 108 ][ 117 ],
   alphaCSR[ 108 ][ 118 ],
   alphaCSR[ 108 ][ 119 ],
   alphaCSR[ 108 ][ 120 ],
   alphaCSR[ 108 ][ 121 ],
   alphaCSR[ 108 ][ 122 ],
   alphaCSR[ 108 ][ 123 ],
   alphaCSR[ 108 ][ 124 ],
   alphaCSR[ 108 ][ 125 ],
   alphaCSR[ 108 ][ 126 ],
   alphaCSR[ 108 ][ 127 ],
   alphaCSR[ 108 ][ 128 ],
   alphaCSR[ 108 ][ 129 ],
   alphaCSR[ 108 ][ 130 ],
   alphaCSR[ 108 ][ 131 ],
   alphaCSR[ 108 ][ 132 ],
   alphaCSR[ 108 ][ 133 ],
   alphaCSR[ 108 ][ 134 ],
   alphaCSR[ 108 ][ 135 ],
   alphaCSR[ 108 ][ 136 ],
   alphaCSR[ 108 ][ 137 ],
   alphaCSR[ 108 ][ 138 ],
   alphaCSR[ 108 ][ 139 ],
   alphaCSR[ 108 ][ 140 ],
   alphaCSR[ 108 ][ 141 ],
   alphaCSR[ 108 ][ 142 ],
   alphaCSR[ 108 ][ 143 ],
   alphaCSR[ 108 ][ 144 ],
   alphaCSR[ 108 ][ 145 ],
   alphaCSR[ 108 ][ 146 ],
   alphaCSR[ 108 ][ 147 ],
   alphaCSR[ 108 ][ 148 ],
   alphaCSR[ 108 ][ 149 ],
   alphaCSR[ 108 ][ 150 ],
   alphaCSR[ 108 ][ 151 ],
   alphaCSR[ 108 ][ 152 ],
   alphaCSR[ 108 ][ 153 ],
   alphaCSR[ 108 ][ 154 ],
   alphaCSR[ 108 ][ 155 ],
   alphaCSR[ 108 ][ 156 ],
   alphaCSR[ 108 ][ 157 ],
   alphaCSR[ 108 ][ 158 ],
   alphaCSR[ 108 ][ 159 ],
   alphaCSR[ 108 ][ 160 ],
   alphaCSR[ 108 ][ 161 ],
   alphaCSR[ 108 ][ 162 ],
   alphaCSR[ 108 ][ 163 ],
   alphaCSR[ 108 ][ 164 ],
   alphaCSR[ 108 ][ 165 ],
   alphaCSR[ 108 ][ 166 ],
   alphaCSR[ 108 ][ 167 ],
   alphaCSR[ 108 ][ 168 ],
   alphaCSR[ 108 ][ 169 ],
   alphaCSR[ 108 ][ 170 ],
   alphaCSR[ 108 ][ 171 ],
   alphaCSR[ 108 ][ 172 ],
   alphaCSR[ 108 ][ 173 ],
   alphaCSR[ 108 ][ 174 ],
   alphaCSR[ 108 ][ 175 ],
   alphaCSR[ 108 ][ 176 ],
   alphaCSR[ 108 ][ 177 ],
   alphaCSR[ 108 ][ 178 ],
   alphaCSR[ 108 ][ 179 ],
   alphaCSR[ 108 ][ 180 ],
   alphaCSR[ 108 ][ 181 ],
   alphaCSR[ 108 ][ 182 ],
   alphaCSR[ 108 ][ 183 ],
   alphaCSR[ 108 ][ 184 ],
   alphaCSR[ 108 ][ 185 ],
   alphaCSR[ 108 ][ 186 ],
   alphaCSR[ 108 ][ 187 ],
   alphaCSR[ 108 ][ 188 ],
   alphaCSR[ 108 ][ 189 ],
   alphaCSR[ 108 ][ 190 ],
   alphaCSR[ 108 ][ 191 ],
   alphaCSR[ 108 ][ 192 ],
   alphaCSR[ 108 ][ 193 ],
   alphaCSR[ 108 ][ 194 ],
   alphaCSR[ 108 ][ 195 ],
   alphaCSR[ 108 ][ 196 ],
   alphaCSR[ 108 ][ 197 ],
   alphaCSR[ 108 ][ 198 ],
   alphaCSR[ 108 ][ 199 ],
   alphaCSR[ 108 ][ 200 ],
   alphaCSR[ 108 ][ 201 ],
   alphaCSR[ 108 ][ 202 ],
   alphaCSR[ 108 ][ 203 ],
   alphaCSR[ 108 ][ 204 ],
   alphaCSR[ 108 ][ 205 ],
   alphaCSR[ 108 ][ 206 ],
   alphaCSR[ 108 ][ 207 ],
   alphaCSR[ 108 ][ 208 ],
   alphaCSR[ 108 ][ 209 ],
   alphaCSR[ 108 ][ 210 ],
   alphaCSR[ 108 ][ 211 ],
   alphaCSR[ 108 ][ 212 ],
   alphaCSR[ 108 ][ 213 ],
   alphaCSR[ 108 ][ 214 ],
   alphaCSR[ 108 ][ 215 ],
   alphaCSR[ 108 ][ 216 ],
   alphaCSR[ 108 ][ 217 ],
   alphaCSR[ 108 ][ 218 ],
   alphaCSR[ 108 ][ 219 ],
   alphaCSR[ 108 ][ 220 ],
   alphaCSR[ 108 ][ 221 ],
   alphaCSR[ 108 ][ 222 ],
   alphaCSR[ 108 ][ 223 ],
   alphaCSR[ 108 ][ 224 ],
   alphaCSR[ 108 ][ 225 ],
   alphaCSR[ 108 ][ 226 ],
   alphaCSR[ 108 ][ 227 ],
   alphaCSR[ 108 ][ 228 ],
   alphaCSR[ 108 ][ 229 ],
   alphaCSR[ 108 ][ 230 ],
   alphaCSR[ 108 ][ 231 ],
   alphaCSR[ 108 ][ 232 ],
   alphaCSR[ 108 ][ 233 ],
   alphaCSR[ 108 ][ 234 ],
   alphaCSR[ 108 ][ 235 ],
   alphaCSR[ 108 ][ 236 ],
   alphaCSR[ 108 ][ 237 ],
   alphaCSR[ 108 ][ 238 ],
   alphaCSR[ 108 ][ 239 ],
   alphaCSR[ 108 ][ 240 ],
   alphaCSR[ 108 ][ 241 ],
   alphaCSR[ 108 ][ 242 ],
   alphaCSR[ 108 ][ 243 ],
   alphaCSR[ 108 ][ 244 ],
   alphaCSR[ 108 ][ 245 ],
   alphaCSR[ 108 ][ 246 ],
   alphaCSR[ 108 ][ 247 ],
   alphaCSR[ 108 ][ 248 ],
   alphaCSR[ 108 ][ 249 ],
   alphaCSR[ 108 ][ 250 ],
   alphaCSR[ 108 ][ 251 ],
   alphaCSR[ 108 ][ 252 ],
   alphaCSR[ 108 ][ 253 ],
   alphaCSR[ 108 ][ 254 ],
   alphaCSR[ 108 ][ 255 ],
   alphaCSR[ 108 ][ 256 ],
   alphaCSR[ 108 ][ 257 ],
   alphaCSR[ 108 ][ 258 ],
   alphaCSR[ 108 ][ 259 ],
   alphaCSR[ 108 ][ 260 ],
   alphaCSR[ 108 ][ 261 ],
   alphaCSR[ 108 ][ 262 ],
   alphaCSR[ 108 ][ 263 ],
   alphaCSR[ 108 ][ 264 ],
   alphaCSR[ 108 ][ 265 ],
   alphaCSR[ 108 ][ 266 ],
   alphaCSR[ 108 ][ 267 ],
   alphaCSR[ 108 ][ 268 ],
   alphaCSR[ 108 ][ 269 ],
   alphaCSR[ 108 ][ 270 ],
   alphaCSR[ 108 ][ 271 ],
   alphaCSR[ 108 ][ 272 ],
   alphaCSR[ 108 ][ 273 ],
   alphaCSR[ 108 ][ 274 ],
   alphaCSR[ 108 ][ 275 ],
   alphaCSR[ 108 ][ 276 ],
   alphaCSR[ 108 ][ 277 ],
   alphaCSR[ 108 ][ 278 ],
   alphaCSR[ 108 ][ 279 ],
   alphaCSR[ 108 ][ 280 ],
   alphaCSR[ 108 ][ 281 ],
   alphaCSR[ 108 ][ 282 ],
   alphaCSR[ 108 ][ 283 ],
   alphaCSR[ 108 ][ 284 ],
   alphaCSR[ 108 ][ 285 ],
   alphaCSR[ 108 ][ 286 ],
   alphaCSR[ 108 ][ 287 ],
   alphaCSR[ 108 ][ 288 ],
   alphaCSR[ 108 ][ 289 ],
   alphaCSR[ 108 ][ 290 ],
   alphaCSR[ 108 ][ 291 ],
   alphaCSR[ 108 ][ 292 ],
   alphaCSR[ 108 ][ 293 ],
   alphaCSR[ 108 ][ 294 ],
   alphaCSR[ 108 ][ 295 ],
   alphaCSR[ 108 ][ 296 ],
   alphaCSR[ 108 ][ 297 ],
   alphaCSR[ 108 ][ 298 ],
   alphaCSR[ 108 ][ 299 ],
   alphaCSR[ 108 ][ 300 ],
   alphaCSR[ 108 ][ 301 ],
   alphaCSR[ 108 ][ 302 ],
   alphaCSR[ 108 ][ 303 ],
   alphaCSR[ 108 ][ 304 ],
   alphaCSR[ 108 ][ 305 ],
   alphaCSR[ 108 ][ 306 ],
   alphaCSR[ 108 ][ 307 ],
   alphaCSR[ 108 ][ 308 ],
   alphaCSR[ 108 ][ 309 ],
   alphaCSR[ 108 ][ 310 ],
   alphaCSR[ 108 ][ 311 ],
   alphaCSR[ 108 ][ 312 ],
   alphaCSR[ 108 ][ 313 ],
   alphaCSR[ 108 ][ 314 ],
   alphaCSR[ 108 ][ 315 ],
   alphaCSR[ 108 ][ 316 ],
   alphaCSR[ 108 ][ 317 ],
   alphaCSR[ 108 ][ 318 ],
   alphaCSR[ 108 ][ 319 ],
   alphaCSR[ 108 ][ 320 ],
   alphaCSR[ 108 ][ 321 ],
   alphaCSR[ 108 ][ 322 ],
   alphaCSR[ 108 ][ 323 ],
   alphaCSR[ 108 ][ 324 ],
   alphaCSR[ 108 ][ 325 ],
   alphaCSR[ 108 ][ 326 ],
   alphaCSR[ 108 ][ 327 ],
   alphaCSR[ 108 ][ 328 ],
   alphaCSR[ 108 ][ 329 ],
   alphaCSR[ 108 ][ 330 ],
   alphaCSR[ 108 ][ 331 ],
   alphaCSR[ 108 ][ 332 ],
   alphaCSR[ 108 ][ 333 ],
   alphaCSR[ 108 ][ 334 ],
   alphaCSR[ 108 ][ 335 ],
   alphaCSR[ 108 ][ 336 ],
   alphaCSR[ 108 ][ 337 ],
   alphaCSR[ 108 ][ 338 ],
   alphaCSR[ 108 ][ 339 ],
   alphaCSR[ 108 ][ 340 ],
   alphaCSR[ 108 ][ 341 ],
   alphaCSR[ 108 ][ 342 ],
   alphaCSR[ 108 ][ 343 ],
   alphaCSR[ 108 ][ 344 ],
   alphaCSR[ 108 ][ 345 ],
   alphaCSR[ 108 ][ 346 ],
   alphaCSR[ 108 ][ 347 ],
   alphaCSR[ 108 ][ 348 ],
   alphaCSR[ 108 ][ 349 ],
   alphaCSR[ 108 ][ 350 ],
   alphaCSR[ 108 ][ 351 ],
   alphaCSR[ 108 ][ 352 ],
   alphaCSR[ 108 ][ 353 ],
   alphaCSR[ 108 ][ 354 ],
   alphaCSR[ 108 ][ 355 ],
   alphaCSR[ 108 ][ 356 ],
   alphaCSR[ 108 ][ 357 ],
   alphaCSR[ 108 ][ 358 ],
   alphaCSR[ 108 ][ 359 ],
   alphaCSR[ 108 ][ 360 ],
   alphaCSR[ 108 ][ 361 ],
   alphaCSR[ 108 ][ 362 ],
   alphaCSR[ 108 ][ 363 ],
   alphaCSR[ 108 ][ 364 ],
   alphaCSR[ 108 ][ 365 ],
   alphaCSR[ 108 ][ 366 ],
   alphaCSR[ 108 ][ 367 ],
   alphaCSR[ 108 ][ 368 ],
   alphaCSR[ 108 ][ 369 ],
   alphaCSR[ 108 ][ 370 ],
   alphaCSR[ 108 ][ 371 ],
   alphaCSR[ 108 ][ 372 ],
   alphaCSR[ 108 ][ 373 ],
   alphaCSR[ 108 ][ 374 ],
   alphaCSR[ 108 ][ 375 ],
   alphaCSR[ 108 ][ 376 ],
   alphaCSR[ 108 ][ 377 ],
   alphaCSR[ 108 ][ 378 ],
   alphaCSR[ 108 ][ 379 ],
   alphaCSR[ 108 ][ 380 ],
   alphaCSR[ 108 ][ 381 ],
   alphaCSR[ 108 ][ 382 ],
   alphaCSR[ 108 ][ 383 ],
   alphaCSR[ 109 ][ 0 ],
   alphaCSR[ 109 ][ 1 ],
   alphaCSR[ 109 ][ 2 ],
   alphaCSR[ 109 ][ 3 ],
   alphaCSR[ 109 ][ 4 ],
   alphaCSR[ 109 ][ 5 ],
   alphaCSR[ 109 ][ 6 ],
   alphaCSR[ 109 ][ 7 ],
   alphaCSR[ 109 ][ 8 ],
   alphaCSR[ 109 ][ 9 ],
   alphaCSR[ 109 ][ 10 ],
   alphaCSR[ 109 ][ 11 ],
   alphaCSR[ 109 ][ 12 ],
   alphaCSR[ 109 ][ 13 ],
   alphaCSR[ 109 ][ 14 ],
   alphaCSR[ 109 ][ 15 ],
   alphaCSR[ 109 ][ 16 ],
   alphaCSR[ 109 ][ 17 ],
   alphaCSR[ 109 ][ 18 ],
   alphaCSR[ 109 ][ 19 ],
   alphaCSR[ 109 ][ 20 ],
   alphaCSR[ 109 ][ 21 ],
   alphaCSR[ 109 ][ 22 ],
   alphaCSR[ 109 ][ 23 ],
   alphaCSR[ 109 ][ 24 ],
   alphaCSR[ 109 ][ 25 ],
   alphaCSR[ 109 ][ 26 ],
   alphaCSR[ 109 ][ 27 ],
   alphaCSR[ 109 ][ 28 ],
   alphaCSR[ 109 ][ 29 ],
   alphaCSR[ 109 ][ 30 ],
   alphaCSR[ 109 ][ 31 ],
   alphaCSR[ 109 ][ 32 ],
   alphaCSR[ 109 ][ 33 ],
   alphaCSR[ 109 ][ 34 ],
   alphaCSR[ 109 ][ 35 ],
   alphaCSR[ 109 ][ 36 ],
   alphaCSR[ 109 ][ 37 ],
   alphaCSR[ 109 ][ 38 ],
   alphaCSR[ 109 ][ 39 ],
   alphaCSR[ 109 ][ 40 ],
   alphaCSR[ 109 ][ 41 ],
   alphaCSR[ 109 ][ 42 ],
   alphaCSR[ 109 ][ 43 ],
   alphaCSR[ 109 ][ 44 ],
   alphaCSR[ 109 ][ 45 ],
   alphaCSR[ 109 ][ 46 ],
   alphaCSR[ 109 ][ 47 ],
   alphaCSR[ 109 ][ 48 ],
   alphaCSR[ 109 ][ 49 ],
   alphaCSR[ 109 ][ 50 ],
   alphaCSR[ 109 ][ 51 ],
   alphaCSR[ 109 ][ 52 ],
   alphaCSR[ 109 ][ 53 ],
   alphaCSR[ 109 ][ 54 ],
   alphaCSR[ 109 ][ 55 ],
   alphaCSR[ 109 ][ 56 ],
   alphaCSR[ 109 ][ 57 ],
   alphaCSR[ 109 ][ 58 ],
   alphaCSR[ 109 ][ 59 ],
   alphaCSR[ 109 ][ 60 ],
   alphaCSR[ 109 ][ 61 ],
   alphaCSR[ 109 ][ 62 ],
   alphaCSR[ 109 ][ 63 ],
   alphaCSR[ 109 ][ 64 ],
   alphaCSR[ 109 ][ 65 ],
   alphaCSR[ 109 ][ 66 ],
   alphaCSR[ 109 ][ 67 ],
   alphaCSR[ 109 ][ 68 ],
   alphaCSR[ 109 ][ 69 ],
   alphaCSR[ 109 ][ 70 ],
   alphaCSR[ 109 ][ 71 ],
   alphaCSR[ 109 ][ 72 ],
   alphaCSR[ 109 ][ 73 ],
   alphaCSR[ 109 ][ 74 ],
   alphaCSR[ 109 ][ 75 ],
   alphaCSR[ 109 ][ 76 ],
   alphaCSR[ 109 ][ 77 ],
   alphaCSR[ 109 ][ 78 ],
   alphaCSR[ 109 ][ 79 ],
   alphaCSR[ 109 ][ 80 ],
   alphaCSR[ 109 ][ 81 ],
   alphaCSR[ 109 ][ 82 ],
   alphaCSR[ 109 ][ 83 ],
   alphaCSR[ 109 ][ 84 ],
   alphaCSR[ 109 ][ 85 ],
   alphaCSR[ 109 ][ 86 ],
   alphaCSR[ 109 ][ 87 ],
   alphaCSR[ 109 ][ 88 ],
   alphaCSR[ 109 ][ 89 ],
   alphaCSR[ 109 ][ 90 ],
   alphaCSR[ 109 ][ 91 ],
   alphaCSR[ 109 ][ 92 ],
   alphaCSR[ 109 ][ 93 ],
   alphaCSR[ 109 ][ 94 ],
   alphaCSR[ 109 ][ 95 ],
   alphaCSR[ 109 ][ 96 ],
   alphaCSR[ 109 ][ 97 ],
   alphaCSR[ 109 ][ 98 ],
   alphaCSR[ 109 ][ 99 ],
   alphaCSR[ 109 ][ 100 ],
   alphaCSR[ 109 ][ 101 ],
   alphaCSR[ 109 ][ 102 ],
   alphaCSR[ 109 ][ 103 ],
   alphaCSR[ 109 ][ 104 ],
   alphaCSR[ 109 ][ 105 ],
   alphaCSR[ 109 ][ 106 ],
   alphaCSR[ 109 ][ 107 ],
   alphaCSR[ 109 ][ 108 ],
   alphaCSR[ 109 ][ 109 ],
   alphaCSR[ 109 ][ 110 ],
   alphaCSR[ 109 ][ 111 ],
   alphaCSR[ 109 ][ 112 ],
   alphaCSR[ 109 ][ 113 ],
   alphaCSR[ 109 ][ 114 ],
   alphaCSR[ 109 ][ 115 ],
   alphaCSR[ 109 ][ 116 ],
   alphaCSR[ 109 ][ 117 ],
   alphaCSR[ 109 ][ 118 ],
   alphaCSR[ 109 ][ 119 ],
   alphaCSR[ 109 ][ 120 ],
   alphaCSR[ 109 ][ 121 ],
   alphaCSR[ 109 ][ 122 ],
   alphaCSR[ 109 ][ 123 ],
   alphaCSR[ 109 ][ 124 ],
   alphaCSR[ 109 ][ 125 ],
   alphaCSR[ 109 ][ 126 ],
   alphaCSR[ 109 ][ 127 ],
   alphaCSR[ 109 ][ 128 ],
   alphaCSR[ 109 ][ 129 ],
   alphaCSR[ 109 ][ 130 ],
   alphaCSR[ 109 ][ 131 ],
   alphaCSR[ 109 ][ 132 ],
   alphaCSR[ 109 ][ 133 ],
   alphaCSR[ 109 ][ 134 ],
   alphaCSR[ 109 ][ 135 ],
   alphaCSR[ 109 ][ 136 ],
   alphaCSR[ 109 ][ 137 ],
   alphaCSR[ 109 ][ 138 ],
   alphaCSR[ 109 ][ 139 ],
   alphaCSR[ 109 ][ 140 ],
   alphaCSR[ 109 ][ 141 ],
   alphaCSR[ 109 ][ 142 ],
   alphaCSR[ 109 ][ 143 ],
   alphaCSR[ 109 ][ 144 ],
   alphaCSR[ 109 ][ 145 ],
   alphaCSR[ 109 ][ 146 ],
   alphaCSR[ 109 ][ 147 ],
   alphaCSR[ 109 ][ 148 ],
   alphaCSR[ 109 ][ 149 ],
   alphaCSR[ 109 ][ 150 ],
   alphaCSR[ 109 ][ 151 ],
   alphaCSR[ 109 ][ 152 ],
   alphaCSR[ 109 ][ 153 ],
   alphaCSR[ 109 ][ 154 ],
   alphaCSR[ 109 ][ 155 ],
   alphaCSR[ 109 ][ 156 ],
   alphaCSR[ 109 ][ 157 ],
   alphaCSR[ 109 ][ 158 ],
   alphaCSR[ 109 ][ 159 ],
   alphaCSR[ 109 ][ 160 ],
   alphaCSR[ 109 ][ 161 ],
   alphaCSR[ 109 ][ 162 ],
   alphaCSR[ 109 ][ 163 ],
   alphaCSR[ 109 ][ 164 ],
   alphaCSR[ 109 ][ 165 ],
   alphaCSR[ 109 ][ 166 ],
   alphaCSR[ 109 ][ 167 ],
   alphaCSR[ 109 ][ 168 ],
   alphaCSR[ 109 ][ 169 ],
   alphaCSR[ 109 ][ 170 ],
   alphaCSR[ 109 ][ 171 ],
   alphaCSR[ 109 ][ 172 ],
   alphaCSR[ 109 ][ 173 ],
   alphaCSR[ 109 ][ 174 ],
   alphaCSR[ 109 ][ 175 ],
   alphaCSR[ 109 ][ 176 ],
   alphaCSR[ 109 ][ 177 ],
   alphaCSR[ 109 ][ 178 ],
   alphaCSR[ 109 ][ 179 ],
   alphaCSR[ 109 ][ 180 ],
   alphaCSR[ 109 ][ 181 ],
   alphaCSR[ 109 ][ 182 ],
   alphaCSR[ 109 ][ 183 ],
   alphaCSR[ 109 ][ 184 ],
   alphaCSR[ 109 ][ 185 ],
   alphaCSR[ 109 ][ 186 ],
   alphaCSR[ 109 ][ 187 ],
   alphaCSR[ 109 ][ 188 ],
   alphaCSR[ 109 ][ 189 ],
   alphaCSR[ 109 ][ 190 ],
   alphaCSR[ 109 ][ 191 ],
   alphaCSR[ 109 ][ 192 ],
   alphaCSR[ 109 ][ 193 ],
   alphaCSR[ 109 ][ 194 ],
   alphaCSR[ 109 ][ 195 ],
   alphaCSR[ 109 ][ 196 ],
   alphaCSR[ 109 ][ 197 ],
   alphaCSR[ 109 ][ 198 ],
   alphaCSR[ 109 ][ 199 ],
   alphaCSR[ 109 ][ 200 ],
   alphaCSR[ 109 ][ 201 ],
   alphaCSR[ 109 ][ 202 ],
   alphaCSR[ 109 ][ 203 ],
   alphaCSR[ 109 ][ 204 ],
   alphaCSR[ 109 ][ 205 ],
   alphaCSR[ 109 ][ 206 ],
   alphaCSR[ 109 ][ 207 ],
   alphaCSR[ 109 ][ 208 ],
   alphaCSR[ 109 ][ 209 ],
   alphaCSR[ 109 ][ 210 ],
   alphaCSR[ 109 ][ 211 ],
   alphaCSR[ 109 ][ 212 ],
   alphaCSR[ 109 ][ 213 ],
   alphaCSR[ 109 ][ 214 ],
   alphaCSR[ 109 ][ 215 ],
   alphaCSR[ 109 ][ 216 ],
   alphaCSR[ 109 ][ 217 ],
   alphaCSR[ 109 ][ 218 ],
   alphaCSR[ 109 ][ 219 ],
   alphaCSR[ 109 ][ 220 ],
   alphaCSR[ 109 ][ 221 ],
   alphaCSR[ 109 ][ 222 ],
   alphaCSR[ 109 ][ 223 ],
   alphaCSR[ 109 ][ 224 ],
   alphaCSR[ 109 ][ 225 ],
   alphaCSR[ 109 ][ 226 ],
   alphaCSR[ 109 ][ 227 ],
   alphaCSR[ 109 ][ 228 ],
   alphaCSR[ 109 ][ 229 ],
   alphaCSR[ 109 ][ 230 ],
   alphaCSR[ 109 ][ 231 ],
   alphaCSR[ 109 ][ 232 ],
   alphaCSR[ 109 ][ 233 ],
   alphaCSR[ 109 ][ 234 ],
   alphaCSR[ 109 ][ 235 ],
   alphaCSR[ 109 ][ 236 ],
   alphaCSR[ 109 ][ 237 ],
   alphaCSR[ 109 ][ 238 ],
   alphaCSR[ 109 ][ 239 ],
   alphaCSR[ 109 ][ 240 ],
   alphaCSR[ 109 ][ 241 ],
   alphaCSR[ 109 ][ 242 ],
   alphaCSR[ 109 ][ 243 ],
   alphaCSR[ 109 ][ 244 ],
   alphaCSR[ 109 ][ 245 ],
   alphaCSR[ 109 ][ 246 ],
   alphaCSR[ 109 ][ 247 ],
   alphaCSR[ 109 ][ 248 ],
   alphaCSR[ 109 ][ 249 ],
   alphaCSR[ 109 ][ 250 ],
   alphaCSR[ 109 ][ 251 ],
   alphaCSR[ 109 ][ 252 ],
   alphaCSR[ 109 ][ 253 ],
   alphaCSR[ 109 ][ 254 ],
   alphaCSR[ 109 ][ 255 ],
   alphaCSR[ 109 ][ 256 ],
   alphaCSR[ 109 ][ 257 ],
   alphaCSR[ 109 ][ 258 ],
   alphaCSR[ 109 ][ 259 ],
   alphaCSR[ 109 ][ 260 ],
   alphaCSR[ 109 ][ 261 ],
   alphaCSR[ 109 ][ 262 ],
   alphaCSR[ 109 ][ 263 ],
   alphaCSR[ 109 ][ 264 ],
   alphaCSR[ 109 ][ 265 ],
   alphaCSR[ 109 ][ 266 ],
   alphaCSR[ 109 ][ 267 ],
   alphaCSR[ 109 ][ 268 ],
   alphaCSR[ 109 ][ 269 ],
   alphaCSR[ 109 ][ 270 ],
   alphaCSR[ 109 ][ 271 ],
   alphaCSR[ 109 ][ 272 ],
   alphaCSR[ 109 ][ 273 ],
   alphaCSR[ 109 ][ 274 ],
   alphaCSR[ 109 ][ 275 ],
   alphaCSR[ 109 ][ 276 ],
   alphaCSR[ 109 ][ 277 ],
   alphaCSR[ 109 ][ 278 ],
   alphaCSR[ 109 ][ 279 ],
   alphaCSR[ 109 ][ 280 ],
   alphaCSR[ 109 ][ 281 ],
   alphaCSR[ 109 ][ 282 ],
   alphaCSR[ 109 ][ 283 ],
   alphaCSR[ 109 ][ 284 ],
   alphaCSR[ 109 ][ 285 ],
   alphaCSR[ 109 ][ 286 ],
   alphaCSR[ 109 ][ 287 ],
   alphaCSR[ 109 ][ 288 ],
   alphaCSR[ 109 ][ 289 ],
   alphaCSR[ 109 ][ 290 ],
   alphaCSR[ 109 ][ 291 ],
   alphaCSR[ 109 ][ 292 ],
   alphaCSR[ 109 ][ 293 ],
   alphaCSR[ 109 ][ 294 ],
   alphaCSR[ 109 ][ 295 ],
   alphaCSR[ 109 ][ 296 ],
   alphaCSR[ 109 ][ 297 ],
   alphaCSR[ 109 ][ 298 ],
   alphaCSR[ 109 ][ 299 ],
   alphaCSR[ 109 ][ 300 ],
   alphaCSR[ 109 ][ 301 ],
   alphaCSR[ 109 ][ 302 ],
   alphaCSR[ 109 ][ 303 ],
   alphaCSR[ 109 ][ 304 ],
   alphaCSR[ 109 ][ 305 ],
   alphaCSR[ 109 ][ 306 ],
   alphaCSR[ 109 ][ 307 ],
   alphaCSR[ 109 ][ 308 ],
   alphaCSR[ 109 ][ 309 ],
   alphaCSR[ 109 ][ 310 ],
   alphaCSR[ 109 ][ 311 ],
   alphaCSR[ 109 ][ 312 ],
   alphaCSR[ 109 ][ 313 ],
   alphaCSR[ 109 ][ 314 ],
   alphaCSR[ 109 ][ 315 ],
   alphaCSR[ 109 ][ 316 ],
   alphaCSR[ 109 ][ 317 ],
   alphaCSR[ 109 ][ 318 ],
   alphaCSR[ 109 ][ 319 ],
   alphaCSR[ 109 ][ 320 ],
   alphaCSR[ 109 ][ 321 ],
   alphaCSR[ 109 ][ 322 ],
   alphaCSR[ 109 ][ 323 ],
   alphaCSR[ 109 ][ 324 ],
   alphaCSR[ 109 ][ 325 ],
   alphaCSR[ 109 ][ 326 ],
   alphaCSR[ 109 ][ 327 ],
   alphaCSR[ 109 ][ 328 ],
   alphaCSR[ 109 ][ 329 ],
   alphaCSR[ 109 ][ 330 ],
   alphaCSR[ 109 ][ 331 ],
   alphaCSR[ 109 ][ 332 ],
   alphaCSR[ 109 ][ 333 ],
   alphaCSR[ 109 ][ 334 ],
   alphaCSR[ 109 ][ 335 ],
   alphaCSR[ 109 ][ 336 ],
   alphaCSR[ 109 ][ 337 ],
   alphaCSR[ 109 ][ 338 ],
   alphaCSR[ 109 ][ 339 ],
   alphaCSR[ 109 ][ 340 ],
   alphaCSR[ 109 ][ 341 ],
   alphaCSR[ 109 ][ 342 ],
   alphaCSR[ 109 ][ 343 ],
   alphaCSR[ 109 ][ 344 ],
   alphaCSR[ 109 ][ 345 ],
   alphaCSR[ 109 ][ 346 ],
   alphaCSR[ 109 ][ 347 ],
   alphaCSR[ 109 ][ 348 ],
   alphaCSR[ 109 ][ 349 ],
   alphaCSR[ 109 ][ 350 ],
   alphaCSR[ 109 ][ 351 ],
   alphaCSR[ 109 ][ 352 ],
   alphaCSR[ 109 ][ 353 ],
   alphaCSR[ 109 ][ 354 ],
   alphaCSR[ 109 ][ 355 ],
   alphaCSR[ 109 ][ 356 ],
   alphaCSR[ 109 ][ 357 ],
   alphaCSR[ 109 ][ 358 ],
   alphaCSR[ 109 ][ 359 ],
   alphaCSR[ 109 ][ 360 ],
   alphaCSR[ 109 ][ 361 ],
   alphaCSR[ 109 ][ 362 ],
   alphaCSR[ 109 ][ 363 ],
   alphaCSR[ 109 ][ 364 ],
   alphaCSR[ 109 ][ 365 ],
   alphaCSR[ 109 ][ 366 ],
   alphaCSR[ 109 ][ 367 ],
   alphaCSR[ 109 ][ 368 ],
   alphaCSR[ 109 ][ 369 ],
   alphaCSR[ 109 ][ 370 ],
   alphaCSR[ 109 ][ 371 ],
   alphaCSR[ 109 ][ 372 ],
   alphaCSR[ 109 ][ 373 ],
   alphaCSR[ 109 ][ 374 ],
   alphaCSR[ 109 ][ 375 ],
   alphaCSR[ 109 ][ 376 ],
   alphaCSR[ 109 ][ 377 ],
   alphaCSR[ 109 ][ 378 ],
   alphaCSR[ 109 ][ 379 ],
   alphaCSR[ 109 ][ 380 ],
   alphaCSR[ 109 ][ 381 ],
   alphaCSR[ 109 ][ 382 ],
   alphaCSR[ 109 ][ 383 ],
   alphaCSR[ 110 ][ 0 ],
   alphaCSR[ 110 ][ 1 ],
   alphaCSR[ 110 ][ 2 ],
   alphaCSR[ 110 ][ 3 ],
   alphaCSR[ 110 ][ 4 ],
   alphaCSR[ 110 ][ 5 ],
   alphaCSR[ 110 ][ 6 ],
   alphaCSR[ 110 ][ 7 ],
   alphaCSR[ 110 ][ 8 ],
   alphaCSR[ 110 ][ 9 ],
   alphaCSR[ 110 ][ 10 ],
   alphaCSR[ 110 ][ 11 ],
   alphaCSR[ 110 ][ 12 ],
   alphaCSR[ 110 ][ 13 ],
   alphaCSR[ 110 ][ 14 ],
   alphaCSR[ 110 ][ 15 ],
   alphaCSR[ 110 ][ 16 ],
   alphaCSR[ 110 ][ 17 ],
   alphaCSR[ 110 ][ 18 ],
   alphaCSR[ 110 ][ 19 ],
   alphaCSR[ 110 ][ 20 ],
   alphaCSR[ 110 ][ 21 ],
   alphaCSR[ 110 ][ 22 ],
   alphaCSR[ 110 ][ 23 ],
   alphaCSR[ 110 ][ 24 ],
   alphaCSR[ 110 ][ 25 ],
   alphaCSR[ 110 ][ 26 ],
   alphaCSR[ 110 ][ 27 ],
   alphaCSR[ 110 ][ 28 ],
   alphaCSR[ 110 ][ 29 ],
   alphaCSR[ 110 ][ 30 ],
   alphaCSR[ 110 ][ 31 ],
   alphaCSR[ 110 ][ 32 ],
   alphaCSR[ 110 ][ 33 ],
   alphaCSR[ 110 ][ 34 ],
   alphaCSR[ 110 ][ 35 ],
   alphaCSR[ 110 ][ 36 ],
   alphaCSR[ 110 ][ 37 ],
   alphaCSR[ 110 ][ 38 ],
   alphaCSR[ 110 ][ 39 ],
   alphaCSR[ 110 ][ 40 ],
   alphaCSR[ 110 ][ 41 ],
   alphaCSR[ 110 ][ 42 ],
   alphaCSR[ 110 ][ 43 ],
   alphaCSR[ 110 ][ 44 ],
   alphaCSR[ 110 ][ 45 ],
   alphaCSR[ 110 ][ 46 ],
   alphaCSR[ 110 ][ 47 ],
   alphaCSR[ 110 ][ 48 ],
   alphaCSR[ 110 ][ 49 ],
   alphaCSR[ 110 ][ 50 ],
   alphaCSR[ 110 ][ 51 ],
   alphaCSR[ 110 ][ 52 ],
   alphaCSR[ 110 ][ 53 ],
   alphaCSR[ 110 ][ 54 ],
   alphaCSR[ 110 ][ 55 ],
   alphaCSR[ 110 ][ 56 ],
   alphaCSR[ 110 ][ 57 ],
   alphaCSR[ 110 ][ 58 ],
   alphaCSR[ 110 ][ 59 ],
   alphaCSR[ 110 ][ 60 ],
   alphaCSR[ 110 ][ 61 ],
   alphaCSR[ 110 ][ 62 ],
   alphaCSR[ 110 ][ 63 ],
   alphaCSR[ 110 ][ 64 ],
   alphaCSR[ 110 ][ 65 ],
   alphaCSR[ 110 ][ 66 ],
   alphaCSR[ 110 ][ 67 ],
   alphaCSR[ 110 ][ 68 ],
   alphaCSR[ 110 ][ 69 ],
   alphaCSR[ 110 ][ 70 ],
   alphaCSR[ 110 ][ 71 ],
   alphaCSR[ 110 ][ 72 ],
   alphaCSR[ 110 ][ 73 ],
   alphaCSR[ 110 ][ 74 ],
   alphaCSR[ 110 ][ 75 ],
   alphaCSR[ 110 ][ 76 ],
   alphaCSR[ 110 ][ 77 ],
   alphaCSR[ 110 ][ 78 ],
   alphaCSR[ 110 ][ 79 ],
   alphaCSR[ 110 ][ 80 ],
   alphaCSR[ 110 ][ 81 ],
   alphaCSR[ 110 ][ 82 ],
   alphaCSR[ 110 ][ 83 ],
   alphaCSR[ 110 ][ 84 ],
   alphaCSR[ 110 ][ 85 ],
   alphaCSR[ 110 ][ 86 ],
   alphaCSR[ 110 ][ 87 ],
   alphaCSR[ 110 ][ 88 ],
   alphaCSR[ 110 ][ 89 ],
   alphaCSR[ 110 ][ 90 ],
   alphaCSR[ 110 ][ 91 ],
   alphaCSR[ 110 ][ 92 ],
   alphaCSR[ 110 ][ 93 ],
   alphaCSR[ 110 ][ 94 ],
   alphaCSR[ 110 ][ 95 ],
   alphaCSR[ 110 ][ 96 ],
   alphaCSR[ 110 ][ 97 ],
   alphaCSR[ 110 ][ 98 ],
   alphaCSR[ 110 ][ 99 ],
   alphaCSR[ 110 ][ 100 ],
   alphaCSR[ 110 ][ 101 ],
   alphaCSR[ 110 ][ 102 ],
   alphaCSR[ 110 ][ 103 ],
   alphaCSR[ 110 ][ 104 ],
   alphaCSR[ 110 ][ 105 ],
   alphaCSR[ 110 ][ 106 ],
   alphaCSR[ 110 ][ 107 ],
   alphaCSR[ 110 ][ 108 ],
   alphaCSR[ 110 ][ 109 ],
   alphaCSR[ 110 ][ 110 ],
   alphaCSR[ 110 ][ 111 ],
   alphaCSR[ 110 ][ 112 ],
   alphaCSR[ 110 ][ 113 ],
   alphaCSR[ 110 ][ 114 ],
   alphaCSR[ 110 ][ 115 ],
   alphaCSR[ 110 ][ 116 ],
   alphaCSR[ 110 ][ 117 ],
   alphaCSR[ 110 ][ 118 ],
   alphaCSR[ 110 ][ 119 ],
   alphaCSR[ 110 ][ 120 ],
   alphaCSR[ 110 ][ 121 ],
   alphaCSR[ 110 ][ 122 ],
   alphaCSR[ 110 ][ 123 ],
   alphaCSR[ 110 ][ 124 ],
   alphaCSR[ 110 ][ 125 ],
   alphaCSR[ 110 ][ 126 ],
   alphaCSR[ 110 ][ 127 ],
   alphaCSR[ 110 ][ 128 ],
   alphaCSR[ 110 ][ 129 ],
   alphaCSR[ 110 ][ 130 ],
   alphaCSR[ 110 ][ 131 ],
   alphaCSR[ 110 ][ 132 ],
   alphaCSR[ 110 ][ 133 ],
   alphaCSR[ 110 ][ 134 ],
   alphaCSR[ 110 ][ 135 ],
   alphaCSR[ 110 ][ 136 ],
   alphaCSR[ 110 ][ 137 ],
   alphaCSR[ 110 ][ 138 ],
   alphaCSR[ 110 ][ 139 ],
   alphaCSR[ 110 ][ 140 ],
   alphaCSR[ 110 ][ 141 ],
   alphaCSR[ 110 ][ 142 ],
   alphaCSR[ 110 ][ 143 ],
   alphaCSR[ 110 ][ 144 ],
   alphaCSR[ 110 ][ 145 ],
   alphaCSR[ 110 ][ 146 ],
   alphaCSR[ 110 ][ 147 ],
   alphaCSR[ 110 ][ 148 ],
   alphaCSR[ 110 ][ 149 ],
   alphaCSR[ 110 ][ 150 ],
   alphaCSR[ 110 ][ 151 ],
   alphaCSR[ 110 ][ 152 ],
   alphaCSR[ 110 ][ 153 ],
   alphaCSR[ 110 ][ 154 ],
   alphaCSR[ 110 ][ 155 ],
   alphaCSR[ 110 ][ 156 ],
   alphaCSR[ 110 ][ 157 ],
   alphaCSR[ 110 ][ 158 ],
   alphaCSR[ 110 ][ 159 ],
   alphaCSR[ 110 ][ 160 ],
   alphaCSR[ 110 ][ 161 ],
   alphaCSR[ 110 ][ 162 ],
   alphaCSR[ 110 ][ 163 ],
   alphaCSR[ 110 ][ 164 ],
   alphaCSR[ 110 ][ 165 ],
   alphaCSR[ 110 ][ 166 ],
   alphaCSR[ 110 ][ 167 ],
   alphaCSR[ 110 ][ 168 ],
   alphaCSR[ 110 ][ 169 ],
   alphaCSR[ 110 ][ 170 ],
   alphaCSR[ 110 ][ 171 ],
   alphaCSR[ 110 ][ 172 ],
   alphaCSR[ 110 ][ 173 ],
   alphaCSR[ 110 ][ 174 ],
   alphaCSR[ 110 ][ 175 ],
   alphaCSR[ 110 ][ 176 ],
   alphaCSR[ 110 ][ 177 ],
   alphaCSR[ 110 ][ 178 ],
   alphaCSR[ 110 ][ 179 ],
   alphaCSR[ 110 ][ 180 ],
   alphaCSR[ 110 ][ 181 ],
   alphaCSR[ 110 ][ 182 ],
   alphaCSR[ 110 ][ 183 ],
   alphaCSR[ 110 ][ 184 ],
   alphaCSR[ 110 ][ 185 ],
   alphaCSR[ 110 ][ 186 ],
   alphaCSR[ 110 ][ 187 ],
   alphaCSR[ 110 ][ 188 ],
   alphaCSR[ 110 ][ 189 ],
   alphaCSR[ 110 ][ 190 ],
   alphaCSR[ 110 ][ 191 ],
   alphaCSR[ 110 ][ 192 ],
   alphaCSR[ 110 ][ 193 ],
   alphaCSR[ 110 ][ 194 ],
   alphaCSR[ 110 ][ 195 ],
   alphaCSR[ 110 ][ 196 ],
   alphaCSR[ 110 ][ 197 ],
   alphaCSR[ 110 ][ 198 ],
   alphaCSR[ 110 ][ 199 ],
   alphaCSR[ 110 ][ 200 ],
   alphaCSR[ 110 ][ 201 ],
   alphaCSR[ 110 ][ 202 ],
   alphaCSR[ 110 ][ 203 ],
   alphaCSR[ 110 ][ 204 ],
   alphaCSR[ 110 ][ 205 ],
   alphaCSR[ 110 ][ 206 ],
   alphaCSR[ 110 ][ 207 ],
   alphaCSR[ 110 ][ 208 ],
   alphaCSR[ 110 ][ 209 ],
   alphaCSR[ 110 ][ 210 ],
   alphaCSR[ 110 ][ 211 ],
   alphaCSR[ 110 ][ 212 ],
   alphaCSR[ 110 ][ 213 ],
   alphaCSR[ 110 ][ 214 ],
   alphaCSR[ 110 ][ 215 ],
   alphaCSR[ 110 ][ 216 ],
   alphaCSR[ 110 ][ 217 ],
   alphaCSR[ 110 ][ 218 ],
   alphaCSR[ 110 ][ 219 ],
   alphaCSR[ 110 ][ 220 ],
   alphaCSR[ 110 ][ 221 ],
   alphaCSR[ 110 ][ 222 ],
   alphaCSR[ 110 ][ 223 ],
   alphaCSR[ 110 ][ 224 ],
   alphaCSR[ 110 ][ 225 ],
   alphaCSR[ 110 ][ 226 ],
   alphaCSR[ 110 ][ 227 ],
   alphaCSR[ 110 ][ 228 ],
   alphaCSR[ 110 ][ 229 ],
   alphaCSR[ 110 ][ 230 ],
   alphaCSR[ 110 ][ 231 ],
   alphaCSR[ 110 ][ 232 ],
   alphaCSR[ 110 ][ 233 ],
   alphaCSR[ 110 ][ 234 ],
   alphaCSR[ 110 ][ 235 ],
   alphaCSR[ 110 ][ 236 ],
   alphaCSR[ 110 ][ 237 ],
   alphaCSR[ 110 ][ 238 ],
   alphaCSR[ 110 ][ 239 ],
   alphaCSR[ 110 ][ 240 ],
   alphaCSR[ 110 ][ 241 ],
   alphaCSR[ 110 ][ 242 ],
   alphaCSR[ 110 ][ 243 ],
   alphaCSR[ 110 ][ 244 ],
   alphaCSR[ 110 ][ 245 ],
   alphaCSR[ 110 ][ 246 ],
   alphaCSR[ 110 ][ 247 ],
   alphaCSR[ 110 ][ 248 ],
   alphaCSR[ 110 ][ 249 ],
   alphaCSR[ 110 ][ 250 ],
   alphaCSR[ 110 ][ 251 ],
   alphaCSR[ 110 ][ 252 ],
   alphaCSR[ 110 ][ 253 ],
   alphaCSR[ 110 ][ 254 ],
   alphaCSR[ 110 ][ 255 ],
   alphaCSR[ 110 ][ 256 ],
   alphaCSR[ 110 ][ 257 ],
   alphaCSR[ 110 ][ 258 ],
   alphaCSR[ 110 ][ 259 ],
   alphaCSR[ 110 ][ 260 ],
   alphaCSR[ 110 ][ 261 ],
   alphaCSR[ 110 ][ 262 ],
   alphaCSR[ 110 ][ 263 ],
   alphaCSR[ 110 ][ 264 ],
   alphaCSR[ 110 ][ 265 ],
   alphaCSR[ 110 ][ 266 ],
   alphaCSR[ 110 ][ 267 ],
   alphaCSR[ 110 ][ 268 ],
   alphaCSR[ 110 ][ 269 ],
   alphaCSR[ 110 ][ 270 ],
   alphaCSR[ 110 ][ 271 ],
   alphaCSR[ 110 ][ 272 ],
   alphaCSR[ 110 ][ 273 ],
   alphaCSR[ 110 ][ 274 ],
   alphaCSR[ 110 ][ 275 ],
   alphaCSR[ 110 ][ 276 ],
   alphaCSR[ 110 ][ 277 ],
   alphaCSR[ 110 ][ 278 ],
   alphaCSR[ 110 ][ 279 ],
   alphaCSR[ 110 ][ 280 ],
   alphaCSR[ 110 ][ 281 ],
   alphaCSR[ 110 ][ 282 ],
   alphaCSR[ 110 ][ 283 ],
   alphaCSR[ 110 ][ 284 ],
   alphaCSR[ 110 ][ 285 ],
   alphaCSR[ 110 ][ 286 ],
   alphaCSR[ 110 ][ 287 ],
   alphaCSR[ 110 ][ 288 ],
   alphaCSR[ 110 ][ 289 ],
   alphaCSR[ 110 ][ 290 ],
   alphaCSR[ 110 ][ 291 ],
   alphaCSR[ 110 ][ 292 ],
   alphaCSR[ 110 ][ 293 ],
   alphaCSR[ 110 ][ 294 ],
   alphaCSR[ 110 ][ 295 ],
   alphaCSR[ 110 ][ 296 ],
   alphaCSR[ 110 ][ 297 ],
   alphaCSR[ 110 ][ 298 ],
   alphaCSR[ 110 ][ 299 ],
   alphaCSR[ 110 ][ 300 ],
   alphaCSR[ 110 ][ 301 ],
   alphaCSR[ 110 ][ 302 ],
   alphaCSR[ 110 ][ 303 ],
   alphaCSR[ 110 ][ 304 ],
   alphaCSR[ 110 ][ 305 ],
   alphaCSR[ 110 ][ 306 ],
   alphaCSR[ 110 ][ 307 ],
   alphaCSR[ 110 ][ 308 ],
   alphaCSR[ 110 ][ 309 ],
   alphaCSR[ 110 ][ 310 ],
   alphaCSR[ 110 ][ 311 ],
   alphaCSR[ 110 ][ 312 ],
   alphaCSR[ 110 ][ 313 ],
   alphaCSR[ 110 ][ 314 ],
   alphaCSR[ 110 ][ 315 ],
   alphaCSR[ 110 ][ 316 ],
   alphaCSR[ 110 ][ 317 ],
   alphaCSR[ 110 ][ 318 ],
   alphaCSR[ 110 ][ 319 ],
   alphaCSR[ 110 ][ 320 ],
   alphaCSR[ 110 ][ 321 ],
   alphaCSR[ 110 ][ 322 ],
   alphaCSR[ 110 ][ 323 ],
   alphaCSR[ 110 ][ 324 ],
   alphaCSR[ 110 ][ 325 ],
   alphaCSR[ 110 ][ 326 ],
   alphaCSR[ 110 ][ 327 ],
   alphaCSR[ 110 ][ 328 ],
   alphaCSR[ 110 ][ 329 ],
   alphaCSR[ 110 ][ 330 ],
   alphaCSR[ 110 ][ 331 ],
   alphaCSR[ 110 ][ 332 ],
   alphaCSR[ 110 ][ 333 ],
   alphaCSR[ 110 ][ 334 ],
   alphaCSR[ 110 ][ 335 ],
   alphaCSR[ 110 ][ 336 ],
   alphaCSR[ 110 ][ 337 ],
   alphaCSR[ 110 ][ 338 ],
   alphaCSR[ 110 ][ 339 ],
   alphaCSR[ 110 ][ 340 ],
   alphaCSR[ 110 ][ 341 ],
   alphaCSR[ 110 ][ 342 ],
   alphaCSR[ 110 ][ 343 ],
   alphaCSR[ 110 ][ 344 ],
   alphaCSR[ 110 ][ 345 ],
   alphaCSR[ 110 ][ 346 ],
   alphaCSR[ 110 ][ 347 ],
   alphaCSR[ 110 ][ 348 ],
   alphaCSR[ 110 ][ 349 ],
   alphaCSR[ 110 ][ 350 ],
   alphaCSR[ 110 ][ 351 ],
   alphaCSR[ 110 ][ 352 ],
   alphaCSR[ 110 ][ 353 ],
   alphaCSR[ 110 ][ 354 ],
   alphaCSR[ 110 ][ 355 ],
   alphaCSR[ 110 ][ 356 ],
   alphaCSR[ 110 ][ 357 ],
   alphaCSR[ 110 ][ 358 ],
   alphaCSR[ 110 ][ 359 ],
   alphaCSR[ 110 ][ 360 ],
   alphaCSR[ 110 ][ 361 ],
   alphaCSR[ 110 ][ 362 ],
   alphaCSR[ 110 ][ 363 ],
   alphaCSR[ 110 ][ 364 ],
   alphaCSR[ 110 ][ 365 ],
   alphaCSR[ 110 ][ 366 ],
   alphaCSR[ 110 ][ 367 ],
   alphaCSR[ 110 ][ 368 ],
   alphaCSR[ 110 ][ 369 ],
   alphaCSR[ 110 ][ 370 ],
   alphaCSR[ 110 ][ 371 ],
   alphaCSR[ 110 ][ 372 ],
   alphaCSR[ 110 ][ 373 ],
   alphaCSR[ 110 ][ 374 ],
   alphaCSR[ 110 ][ 375 ],
   alphaCSR[ 110 ][ 376 ],
   alphaCSR[ 110 ][ 377 ],
   alphaCSR[ 110 ][ 378 ],
   alphaCSR[ 110 ][ 379 ],
   alphaCSR[ 110 ][ 380 ],
   alphaCSR[ 110 ][ 381 ],
   alphaCSR[ 110 ][ 382 ],
   alphaCSR[ 110 ][ 383 ],
   alphaCSR[ 111 ][ 0 ],
   alphaCSR[ 111 ][ 1 ],
   alphaCSR[ 111 ][ 2 ],
   alphaCSR[ 111 ][ 3 ],
   alphaCSR[ 111 ][ 4 ],
   alphaCSR[ 111 ][ 5 ],
   alphaCSR[ 111 ][ 6 ],
   alphaCSR[ 111 ][ 7 ],
   alphaCSR[ 111 ][ 8 ],
   alphaCSR[ 111 ][ 9 ],
   alphaCSR[ 111 ][ 10 ],
   alphaCSR[ 111 ][ 11 ],
   alphaCSR[ 111 ][ 12 ],
   alphaCSR[ 111 ][ 13 ],
   alphaCSR[ 111 ][ 14 ],
   alphaCSR[ 111 ][ 15 ],
   alphaCSR[ 111 ][ 16 ],
   alphaCSR[ 111 ][ 17 ],
   alphaCSR[ 111 ][ 18 ],
   alphaCSR[ 111 ][ 19 ],
   alphaCSR[ 111 ][ 20 ],
   alphaCSR[ 111 ][ 21 ],
   alphaCSR[ 111 ][ 22 ],
   alphaCSR[ 111 ][ 23 ],
   alphaCSR[ 111 ][ 24 ],
   alphaCSR[ 111 ][ 25 ],
   alphaCSR[ 111 ][ 26 ],
   alphaCSR[ 111 ][ 27 ],
   alphaCSR[ 111 ][ 28 ],
   alphaCSR[ 111 ][ 29 ],
   alphaCSR[ 111 ][ 30 ],
   alphaCSR[ 111 ][ 31 ],
   alphaCSR[ 111 ][ 32 ],
   alphaCSR[ 111 ][ 33 ],
   alphaCSR[ 111 ][ 34 ],
   alphaCSR[ 111 ][ 35 ],
   alphaCSR[ 111 ][ 36 ],
   alphaCSR[ 111 ][ 37 ],
   alphaCSR[ 111 ][ 38 ],
   alphaCSR[ 111 ][ 39 ],
   alphaCSR[ 111 ][ 40 ],
   alphaCSR[ 111 ][ 41 ],
   alphaCSR[ 111 ][ 42 ],
   alphaCSR[ 111 ][ 43 ],
   alphaCSR[ 111 ][ 44 ],
   alphaCSR[ 111 ][ 45 ],
   alphaCSR[ 111 ][ 46 ],
   alphaCSR[ 111 ][ 47 ],
   alphaCSR[ 111 ][ 48 ],
   alphaCSR[ 111 ][ 49 ],
   alphaCSR[ 111 ][ 50 ],
   alphaCSR[ 111 ][ 51 ],
   alphaCSR[ 111 ][ 52 ],
   alphaCSR[ 111 ][ 53 ],
   alphaCSR[ 111 ][ 54 ],
   alphaCSR[ 111 ][ 55 ],
   alphaCSR[ 111 ][ 56 ],
   alphaCSR[ 111 ][ 57 ],
   alphaCSR[ 111 ][ 58 ],
   alphaCSR[ 111 ][ 59 ],
   alphaCSR[ 111 ][ 60 ],
   alphaCSR[ 111 ][ 61 ],
   alphaCSR[ 111 ][ 62 ],
   alphaCSR[ 111 ][ 63 ],
   alphaCSR[ 111 ][ 64 ],
   alphaCSR[ 111 ][ 65 ],
   alphaCSR[ 111 ][ 66 ],
   alphaCSR[ 111 ][ 67 ],
   alphaCSR[ 111 ][ 68 ],
   alphaCSR[ 111 ][ 69 ],
   alphaCSR[ 111 ][ 70 ],
   alphaCSR[ 111 ][ 71 ],
   alphaCSR[ 111 ][ 72 ],
   alphaCSR[ 111 ][ 73 ],
   alphaCSR[ 111 ][ 74 ],
   alphaCSR[ 111 ][ 75 ],
   alphaCSR[ 111 ][ 76 ],
   alphaCSR[ 111 ][ 77 ],
   alphaCSR[ 111 ][ 78 ],
   alphaCSR[ 111 ][ 79 ],
   alphaCSR[ 111 ][ 80 ],
   alphaCSR[ 111 ][ 81 ],
   alphaCSR[ 111 ][ 82 ],
   alphaCSR[ 111 ][ 83 ],
   alphaCSR[ 111 ][ 84 ],
   alphaCSR[ 111 ][ 85 ],
   alphaCSR[ 111 ][ 86 ],
   alphaCSR[ 111 ][ 87 ],
   alphaCSR[ 111 ][ 88 ],
   alphaCSR[ 111 ][ 89 ],
   alphaCSR[ 111 ][ 90 ],
   alphaCSR[ 111 ][ 91 ],
   alphaCSR[ 111 ][ 92 ],
   alphaCSR[ 111 ][ 93 ],
   alphaCSR[ 111 ][ 94 ],
   alphaCSR[ 111 ][ 95 ],
   alphaCSR[ 111 ][ 96 ],
   alphaCSR[ 111 ][ 97 ],
   alphaCSR[ 111 ][ 98 ],
   alphaCSR[ 111 ][ 99 ],
   alphaCSR[ 111 ][ 100 ],
   alphaCSR[ 111 ][ 101 ],
   alphaCSR[ 111 ][ 102 ],
   alphaCSR[ 111 ][ 103 ],
   alphaCSR[ 111 ][ 104 ],
   alphaCSR[ 111 ][ 105 ],
   alphaCSR[ 111 ][ 106 ],
   alphaCSR[ 111 ][ 107 ],
   alphaCSR[ 111 ][ 108 ],
   alphaCSR[ 111 ][ 109 ],
   alphaCSR[ 111 ][ 110 ],
   alphaCSR[ 111 ][ 111 ],
   alphaCSR[ 111 ][ 112 ],
   alphaCSR[ 111 ][ 113 ],
   alphaCSR[ 111 ][ 114 ],
   alphaCSR[ 111 ][ 115 ],
   alphaCSR[ 111 ][ 116 ],
   alphaCSR[ 111 ][ 117 ],
   alphaCSR[ 111 ][ 118 ],
   alphaCSR[ 111 ][ 119 ],
   alphaCSR[ 111 ][ 120 ],
   alphaCSR[ 111 ][ 121 ],
   alphaCSR[ 111 ][ 122 ],
   alphaCSR[ 111 ][ 123 ],
   alphaCSR[ 111 ][ 124 ],
   alphaCSR[ 111 ][ 125 ],
   alphaCSR[ 111 ][ 126 ],
   alphaCSR[ 111 ][ 127 ],
   alphaCSR[ 111 ][ 128 ],
   alphaCSR[ 111 ][ 129 ],
   alphaCSR[ 111 ][ 130 ],
   alphaCSR[ 111 ][ 131 ],
   alphaCSR[ 111 ][ 132 ],
   alphaCSR[ 111 ][ 133 ],
   alphaCSR[ 111 ][ 134 ],
   alphaCSR[ 111 ][ 135 ],
   alphaCSR[ 111 ][ 136 ],
   alphaCSR[ 111 ][ 137 ],
   alphaCSR[ 111 ][ 138 ],
   alphaCSR[ 111 ][ 139 ],
   alphaCSR[ 111 ][ 140 ],
   alphaCSR[ 111 ][ 141 ],
   alphaCSR[ 111 ][ 142 ],
   alphaCSR[ 111 ][ 143 ],
   alphaCSR[ 111 ][ 144 ],
   alphaCSR[ 111 ][ 145 ],
   alphaCSR[ 111 ][ 146 ],
   alphaCSR[ 111 ][ 147 ],
   alphaCSR[ 111 ][ 148 ],
   alphaCSR[ 111 ][ 149 ],
   alphaCSR[ 111 ][ 150 ],
   alphaCSR[ 111 ][ 151 ],
   alphaCSR[ 111 ][ 152 ],
   alphaCSR[ 111 ][ 153 ],
   alphaCSR[ 111 ][ 154 ],
   alphaCSR[ 111 ][ 155 ],
   alphaCSR[ 111 ][ 156 ],
   alphaCSR[ 111 ][ 157 ],
   alphaCSR[ 111 ][ 158 ],
   alphaCSR[ 111 ][ 159 ],
   alphaCSR[ 111 ][ 160 ],
   alphaCSR[ 111 ][ 161 ],
   alphaCSR[ 111 ][ 162 ],
   alphaCSR[ 111 ][ 163 ],
   alphaCSR[ 111 ][ 164 ],
   alphaCSR[ 111 ][ 165 ],
   alphaCSR[ 111 ][ 166 ],
   alphaCSR[ 111 ][ 167 ],
   alphaCSR[ 111 ][ 168 ],
   alphaCSR[ 111 ][ 169 ],
   alphaCSR[ 111 ][ 170 ],
   alphaCSR[ 111 ][ 171 ],
   alphaCSR[ 111 ][ 172 ],
   alphaCSR[ 111 ][ 173 ],
   alphaCSR[ 111 ][ 174 ],
   alphaCSR[ 111 ][ 175 ],
   alphaCSR[ 111 ][ 176 ],
   alphaCSR[ 111 ][ 177 ],
   alphaCSR[ 111 ][ 178 ],
   alphaCSR[ 111 ][ 179 ],
   alphaCSR[ 111 ][ 180 ],
   alphaCSR[ 111 ][ 181 ],
   alphaCSR[ 111 ][ 182 ],
   alphaCSR[ 111 ][ 183 ],
   alphaCSR[ 111 ][ 184 ],
   alphaCSR[ 111 ][ 185 ],
   alphaCSR[ 111 ][ 186 ],
   alphaCSR[ 111 ][ 187 ],
   alphaCSR[ 111 ][ 188 ],
   alphaCSR[ 111 ][ 189 ],
   alphaCSR[ 111 ][ 190 ],
   alphaCSR[ 111 ][ 191 ],
   alphaCSR[ 111 ][ 192 ],
   alphaCSR[ 111 ][ 193 ],
   alphaCSR[ 111 ][ 194 ],
   alphaCSR[ 111 ][ 195 ],
   alphaCSR[ 111 ][ 196 ],
   alphaCSR[ 111 ][ 197 ],
   alphaCSR[ 111 ][ 198 ],
   alphaCSR[ 111 ][ 199 ],
   alphaCSR[ 111 ][ 200 ],
   alphaCSR[ 111 ][ 201 ],
   alphaCSR[ 111 ][ 202 ],
   alphaCSR[ 111 ][ 203 ],
   alphaCSR[ 111 ][ 204 ],
   alphaCSR[ 111 ][ 205 ],
   alphaCSR[ 111 ][ 206 ],
   alphaCSR[ 111 ][ 207 ],
   alphaCSR[ 111 ][ 208 ],
   alphaCSR[ 111 ][ 209 ],
   alphaCSR[ 111 ][ 210 ],
   alphaCSR[ 111 ][ 211 ],
   alphaCSR[ 111 ][ 212 ],
   alphaCSR[ 111 ][ 213 ],
   alphaCSR[ 111 ][ 214 ],
   alphaCSR[ 111 ][ 215 ],
   alphaCSR[ 111 ][ 216 ],
   alphaCSR[ 111 ][ 217 ],
   alphaCSR[ 111 ][ 218 ],
   alphaCSR[ 111 ][ 219 ],
   alphaCSR[ 111 ][ 220 ],
   alphaCSR[ 111 ][ 221 ],
   alphaCSR[ 111 ][ 222 ],
   alphaCSR[ 111 ][ 223 ],
   alphaCSR[ 111 ][ 224 ],
   alphaCSR[ 111 ][ 225 ],
   alphaCSR[ 111 ][ 226 ],
   alphaCSR[ 111 ][ 227 ],
   alphaCSR[ 111 ][ 228 ],
   alphaCSR[ 111 ][ 229 ],
   alphaCSR[ 111 ][ 230 ],
   alphaCSR[ 111 ][ 231 ],
   alphaCSR[ 111 ][ 232 ],
   alphaCSR[ 111 ][ 233 ],
   alphaCSR[ 111 ][ 234 ],
   alphaCSR[ 111 ][ 235 ],
   alphaCSR[ 111 ][ 236 ],
   alphaCSR[ 111 ][ 237 ],
   alphaCSR[ 111 ][ 238 ],
   alphaCSR[ 111 ][ 239 ],
   alphaCSR[ 111 ][ 240 ],
   alphaCSR[ 111 ][ 241 ],
   alphaCSR[ 111 ][ 242 ],
   alphaCSR[ 111 ][ 243 ],
   alphaCSR[ 111 ][ 244 ],
   alphaCSR[ 111 ][ 245 ],
   alphaCSR[ 111 ][ 246 ],
   alphaCSR[ 111 ][ 247 ],
   alphaCSR[ 111 ][ 248 ],
   alphaCSR[ 111 ][ 249 ],
   alphaCSR[ 111 ][ 250 ],
   alphaCSR[ 111 ][ 251 ],
   alphaCSR[ 111 ][ 252 ],
   alphaCSR[ 111 ][ 253 ],
   alphaCSR[ 111 ][ 254 ],
   alphaCSR[ 111 ][ 255 ],
   alphaCSR[ 111 ][ 256 ],
   alphaCSR[ 111 ][ 257 ],
   alphaCSR[ 111 ][ 258 ],
   alphaCSR[ 111 ][ 259 ],
   alphaCSR[ 111 ][ 260 ],
   alphaCSR[ 111 ][ 261 ],
   alphaCSR[ 111 ][ 262 ],
   alphaCSR[ 111 ][ 263 ],
   alphaCSR[ 111 ][ 264 ],
   alphaCSR[ 111 ][ 265 ],
   alphaCSR[ 111 ][ 266 ],
   alphaCSR[ 111 ][ 267 ],
   alphaCSR[ 111 ][ 268 ],
   alphaCSR[ 111 ][ 269 ],
   alphaCSR[ 111 ][ 270 ],
   alphaCSR[ 111 ][ 271 ],
   alphaCSR[ 111 ][ 272 ],
   alphaCSR[ 111 ][ 273 ],
   alphaCSR[ 111 ][ 274 ],
   alphaCSR[ 111 ][ 275 ],
   alphaCSR[ 111 ][ 276 ],
   alphaCSR[ 111 ][ 277 ],
   alphaCSR[ 111 ][ 278 ],
   alphaCSR[ 111 ][ 279 ],
   alphaCSR[ 111 ][ 280 ],
   alphaCSR[ 111 ][ 281 ],
   alphaCSR[ 111 ][ 282 ],
   alphaCSR[ 111 ][ 283 ],
   alphaCSR[ 111 ][ 284 ],
   alphaCSR[ 111 ][ 285 ],
   alphaCSR[ 111 ][ 286 ],
   alphaCSR[ 111 ][ 287 ],
   alphaCSR[ 111 ][ 288 ],
   alphaCSR[ 111 ][ 289 ],
   alphaCSR[ 111 ][ 290 ],
   alphaCSR[ 111 ][ 291 ],
   alphaCSR[ 111 ][ 292 ],
   alphaCSR[ 111 ][ 293 ],
   alphaCSR[ 111 ][ 294 ],
   alphaCSR[ 111 ][ 295 ],
   alphaCSR[ 111 ][ 296 ],
   alphaCSR[ 111 ][ 297 ],
   alphaCSR[ 111 ][ 298 ],
   alphaCSR[ 111 ][ 299 ],
   alphaCSR[ 111 ][ 300 ],
   alphaCSR[ 111 ][ 301 ],
   alphaCSR[ 111 ][ 302 ],
   alphaCSR[ 111 ][ 303 ],
   alphaCSR[ 111 ][ 304 ],
   alphaCSR[ 111 ][ 305 ],
   alphaCSR[ 111 ][ 306 ],
   alphaCSR[ 111 ][ 307 ],
   alphaCSR[ 111 ][ 308 ],
   alphaCSR[ 111 ][ 309 ],
   alphaCSR[ 111 ][ 310 ],
   alphaCSR[ 111 ][ 311 ],
   alphaCSR[ 111 ][ 312 ],
   alphaCSR[ 111 ][ 313 ],
   alphaCSR[ 111 ][ 314 ],
   alphaCSR[ 111 ][ 315 ],
   alphaCSR[ 111 ][ 316 ],
   alphaCSR[ 111 ][ 317 ],
   alphaCSR[ 111 ][ 318 ],
   alphaCSR[ 111 ][ 319 ],
   alphaCSR[ 111 ][ 320 ],
   alphaCSR[ 111 ][ 321 ],
   alphaCSR[ 111 ][ 322 ],
   alphaCSR[ 111 ][ 323 ],
   alphaCSR[ 111 ][ 324 ],
   alphaCSR[ 111 ][ 325 ],
   alphaCSR[ 111 ][ 326 ],
   alphaCSR[ 111 ][ 327 ],
   alphaCSR[ 111 ][ 328 ],
   alphaCSR[ 111 ][ 329 ],
   alphaCSR[ 111 ][ 330 ],
   alphaCSR[ 111 ][ 331 ],
   alphaCSR[ 111 ][ 332 ],
   alphaCSR[ 111 ][ 333 ],
   alphaCSR[ 111 ][ 334 ],
   alphaCSR[ 111 ][ 335 ],
   alphaCSR[ 111 ][ 336 ],
   alphaCSR[ 111 ][ 337 ],
   alphaCSR[ 111 ][ 338 ],
   alphaCSR[ 111 ][ 339 ],
   alphaCSR[ 111 ][ 340 ],
   alphaCSR[ 111 ][ 341 ],
   alphaCSR[ 111 ][ 342 ],
   alphaCSR[ 111 ][ 343 ],
   alphaCSR[ 111 ][ 344 ],
   alphaCSR[ 111 ][ 345 ],
   alphaCSR[ 111 ][ 346 ],
   alphaCSR[ 111 ][ 347 ],
   alphaCSR[ 111 ][ 348 ],
   alphaCSR[ 111 ][ 349 ],
   alphaCSR[ 111 ][ 350 ],
   alphaCSR[ 111 ][ 351 ],
   alphaCSR[ 111 ][ 352 ],
   alphaCSR[ 111 ][ 353 ],
   alphaCSR[ 111 ][ 354 ],
   alphaCSR[ 111 ][ 355 ],
   alphaCSR[ 111 ][ 356 ],
   alphaCSR[ 111 ][ 357 ],
   alphaCSR[ 111 ][ 358 ],
   alphaCSR[ 111 ][ 359 ],
   alphaCSR[ 111 ][ 360 ],
   alphaCSR[ 111 ][ 361 ],
   alphaCSR[ 111 ][ 362 ],
   alphaCSR[ 111 ][ 363 ],
   alphaCSR[ 111 ][ 364 ],
   alphaCSR[ 111 ][ 365 ],
   alphaCSR[ 111 ][ 366 ],
   alphaCSR[ 111 ][ 367 ],
   alphaCSR[ 111 ][ 368 ],
   alphaCSR[ 111 ][ 369 ],
   alphaCSR[ 111 ][ 370 ],
   alphaCSR[ 111 ][ 371 ],
   alphaCSR[ 111 ][ 372 ],
   alphaCSR[ 111 ][ 373 ],
   alphaCSR[ 111 ][ 374 ],
   alphaCSR[ 111 ][ 375 ],
   alphaCSR[ 111 ][ 376 ],
   alphaCSR[ 111 ][ 377 ],
   alphaCSR[ 111 ][ 378 ],
   alphaCSR[ 111 ][ 379 ],
   alphaCSR[ 111 ][ 380 ],
   alphaCSR[ 111 ][ 381 ],
   alphaCSR[ 111 ][ 382 ],
   alphaCSR[ 111 ][ 383 ],
   alphaCSR[ 112 ][ 0 ],
   alphaCSR[ 112 ][ 1 ],
   alphaCSR[ 112 ][ 2 ],
   alphaCSR[ 112 ][ 3 ],
   alphaCSR[ 112 ][ 4 ],
   alphaCSR[ 112 ][ 5 ],
   alphaCSR[ 112 ][ 6 ],
   alphaCSR[ 112 ][ 7 ],
   alphaCSR[ 112 ][ 8 ],
   alphaCSR[ 112 ][ 9 ],
   alphaCSR[ 112 ][ 10 ],
   alphaCSR[ 112 ][ 11 ],
   alphaCSR[ 112 ][ 12 ],
   alphaCSR[ 112 ][ 13 ],
   alphaCSR[ 112 ][ 14 ],
   alphaCSR[ 112 ][ 15 ],
   alphaCSR[ 112 ][ 16 ],
   alphaCSR[ 112 ][ 17 ],
   alphaCSR[ 112 ][ 18 ],
   alphaCSR[ 112 ][ 19 ],
   alphaCSR[ 112 ][ 20 ],
   alphaCSR[ 112 ][ 21 ],
   alphaCSR[ 112 ][ 22 ],
   alphaCSR[ 112 ][ 23 ],
   alphaCSR[ 112 ][ 24 ],
   alphaCSR[ 112 ][ 25 ],
   alphaCSR[ 112 ][ 26 ],
   alphaCSR[ 112 ][ 27 ],
   alphaCSR[ 112 ][ 28 ],
   alphaCSR[ 112 ][ 29 ],
   alphaCSR[ 112 ][ 30 ],
   alphaCSR[ 112 ][ 31 ],
   alphaCSR[ 112 ][ 32 ],
   alphaCSR[ 112 ][ 33 ],
   alphaCSR[ 112 ][ 34 ],
   alphaCSR[ 112 ][ 35 ],
   alphaCSR[ 112 ][ 36 ],
   alphaCSR[ 112 ][ 37 ],
   alphaCSR[ 112 ][ 38 ],
   alphaCSR[ 112 ][ 39 ],
   alphaCSR[ 112 ][ 40 ],
   alphaCSR[ 112 ][ 41 ],
   alphaCSR[ 112 ][ 42 ],
   alphaCSR[ 112 ][ 43 ],
   alphaCSR[ 112 ][ 44 ],
   alphaCSR[ 112 ][ 45 ],
   alphaCSR[ 112 ][ 46 ],
   alphaCSR[ 112 ][ 47 ],
   alphaCSR[ 112 ][ 48 ],
   alphaCSR[ 112 ][ 49 ],
   alphaCSR[ 112 ][ 50 ],
   alphaCSR[ 112 ][ 51 ],
   alphaCSR[ 112 ][ 52 ],
   alphaCSR[ 112 ][ 53 ],
   alphaCSR[ 112 ][ 54 ],
   alphaCSR[ 112 ][ 55 ],
   alphaCSR[ 112 ][ 56 ],
   alphaCSR[ 112 ][ 57 ],
   alphaCSR[ 112 ][ 58 ],
   alphaCSR[ 112 ][ 59 ],
   alphaCSR[ 112 ][ 60 ],
   alphaCSR[ 112 ][ 61 ],
   alphaCSR[ 112 ][ 62 ],
   alphaCSR[ 112 ][ 63 ],
   alphaCSR[ 112 ][ 64 ],
   alphaCSR[ 112 ][ 65 ],
   alphaCSR[ 112 ][ 66 ],
   alphaCSR[ 112 ][ 67 ],
   alphaCSR[ 112 ][ 68 ],
   alphaCSR[ 112 ][ 69 ],
   alphaCSR[ 112 ][ 70 ],
   alphaCSR[ 112 ][ 71 ],
   alphaCSR[ 112 ][ 72 ],
   alphaCSR[ 112 ][ 73 ],
   alphaCSR[ 112 ][ 74 ],
   alphaCSR[ 112 ][ 75 ],
   alphaCSR[ 112 ][ 76 ],
   alphaCSR[ 112 ][ 77 ],
   alphaCSR[ 112 ][ 78 ],
   alphaCSR[ 112 ][ 79 ],
   alphaCSR[ 112 ][ 80 ],
   alphaCSR[ 112 ][ 81 ],
   alphaCSR[ 112 ][ 82 ],
   alphaCSR[ 112 ][ 83 ],
   alphaCSR[ 112 ][ 84 ],
   alphaCSR[ 112 ][ 85 ],
   alphaCSR[ 112 ][ 86 ],
   alphaCSR[ 112 ][ 87 ],
   alphaCSR[ 112 ][ 88 ],
   alphaCSR[ 112 ][ 89 ],
   alphaCSR[ 112 ][ 90 ],
   alphaCSR[ 112 ][ 91 ],
   alphaCSR[ 112 ][ 92 ],
   alphaCSR[ 112 ][ 93 ],
   alphaCSR[ 112 ][ 94 ],
   alphaCSR[ 112 ][ 95 ],
   alphaCSR[ 112 ][ 96 ],
   alphaCSR[ 112 ][ 97 ],
   alphaCSR[ 112 ][ 98 ],
   alphaCSR[ 112 ][ 99 ],
   alphaCSR[ 112 ][ 100 ],
   alphaCSR[ 112 ][ 101 ],
   alphaCSR[ 112 ][ 102 ],
   alphaCSR[ 112 ][ 103 ],
   alphaCSR[ 112 ][ 104 ],
   alphaCSR[ 112 ][ 105 ],
   alphaCSR[ 112 ][ 106 ],
   alphaCSR[ 112 ][ 107 ],
   alphaCSR[ 112 ][ 108 ],
   alphaCSR[ 112 ][ 109 ],
   alphaCSR[ 112 ][ 110 ],
   alphaCSR[ 112 ][ 111 ],
   alphaCSR[ 112 ][ 112 ],
   alphaCSR[ 112 ][ 113 ],
   alphaCSR[ 112 ][ 114 ],
   alphaCSR[ 112 ][ 115 ],
   alphaCSR[ 112 ][ 116 ],
   alphaCSR[ 112 ][ 117 ],
   alphaCSR[ 112 ][ 118 ],
   alphaCSR[ 112 ][ 119 ],
   alphaCSR[ 112 ][ 120 ],
   alphaCSR[ 112 ][ 121 ],
   alphaCSR[ 112 ][ 122 ],
   alphaCSR[ 112 ][ 123 ],
   alphaCSR[ 112 ][ 124 ],
   alphaCSR[ 112 ][ 125 ],
   alphaCSR[ 112 ][ 126 ],
   alphaCSR[ 112 ][ 127 ],
   alphaCSR[ 112 ][ 128 ],
   alphaCSR[ 112 ][ 129 ],
   alphaCSR[ 112 ][ 130 ],
   alphaCSR[ 112 ][ 131 ],
   alphaCSR[ 112 ][ 132 ],
   alphaCSR[ 112 ][ 133 ],
   alphaCSR[ 112 ][ 134 ],
   alphaCSR[ 112 ][ 135 ],
   alphaCSR[ 112 ][ 136 ],
   alphaCSR[ 112 ][ 137 ],
   alphaCSR[ 112 ][ 138 ],
   alphaCSR[ 112 ][ 139 ],
   alphaCSR[ 112 ][ 140 ],
   alphaCSR[ 112 ][ 141 ],
   alphaCSR[ 112 ][ 142 ],
   alphaCSR[ 112 ][ 143 ],
   alphaCSR[ 112 ][ 144 ],
   alphaCSR[ 112 ][ 145 ],
   alphaCSR[ 112 ][ 146 ],
   alphaCSR[ 112 ][ 147 ],
   alphaCSR[ 112 ][ 148 ],
   alphaCSR[ 112 ][ 149 ],
   alphaCSR[ 112 ][ 150 ],
   alphaCSR[ 112 ][ 151 ],
   alphaCSR[ 112 ][ 152 ],
   alphaCSR[ 112 ][ 153 ],
   alphaCSR[ 112 ][ 154 ],
   alphaCSR[ 112 ][ 155 ],
   alphaCSR[ 112 ][ 156 ],
   alphaCSR[ 112 ][ 157 ],
   alphaCSR[ 112 ][ 158 ],
   alphaCSR[ 112 ][ 159 ],
   alphaCSR[ 112 ][ 160 ],
   alphaCSR[ 112 ][ 161 ],
   alphaCSR[ 112 ][ 162 ],
   alphaCSR[ 112 ][ 163 ],
   alphaCSR[ 112 ][ 164 ],
   alphaCSR[ 112 ][ 165 ],
   alphaCSR[ 112 ][ 166 ],
   alphaCSR[ 112 ][ 167 ],
   alphaCSR[ 112 ][ 168 ],
   alphaCSR[ 112 ][ 169 ],
   alphaCSR[ 112 ][ 170 ],
   alphaCSR[ 112 ][ 171 ],
   alphaCSR[ 112 ][ 172 ],
   alphaCSR[ 112 ][ 173 ],
   alphaCSR[ 112 ][ 174 ],
   alphaCSR[ 112 ][ 175 ],
   alphaCSR[ 112 ][ 176 ],
   alphaCSR[ 112 ][ 177 ],
   alphaCSR[ 112 ][ 178 ],
   alphaCSR[ 112 ][ 179 ],
   alphaCSR[ 112 ][ 180 ],
   alphaCSR[ 112 ][ 181 ],
   alphaCSR[ 112 ][ 182 ],
   alphaCSR[ 112 ][ 183 ],
   alphaCSR[ 112 ][ 184 ],
   alphaCSR[ 112 ][ 185 ],
   alphaCSR[ 112 ][ 186 ],
   alphaCSR[ 112 ][ 187 ],
   alphaCSR[ 112 ][ 188 ],
   alphaCSR[ 112 ][ 189 ],
   alphaCSR[ 112 ][ 190 ],
   alphaCSR[ 112 ][ 191 ],
   alphaCSR[ 112 ][ 192 ],
   alphaCSR[ 112 ][ 193 ],
   alphaCSR[ 112 ][ 194 ],
   alphaCSR[ 112 ][ 195 ],
   alphaCSR[ 112 ][ 196 ],
   alphaCSR[ 112 ][ 197 ],
   alphaCSR[ 112 ][ 198 ],
   alphaCSR[ 112 ][ 199 ],
   alphaCSR[ 112 ][ 200 ],
   alphaCSR[ 112 ][ 201 ],
   alphaCSR[ 112 ][ 202 ],
   alphaCSR[ 112 ][ 203 ],
   alphaCSR[ 112 ][ 204 ],
   alphaCSR[ 112 ][ 205 ],
   alphaCSR[ 112 ][ 206 ],
   alphaCSR[ 112 ][ 207 ],
   alphaCSR[ 112 ][ 208 ],
   alphaCSR[ 112 ][ 209 ],
   alphaCSR[ 112 ][ 210 ],
   alphaCSR[ 112 ][ 211 ],
   alphaCSR[ 112 ][ 212 ],
   alphaCSR[ 112 ][ 213 ],
   alphaCSR[ 112 ][ 214 ],
   alphaCSR[ 112 ][ 215 ],
   alphaCSR[ 112 ][ 216 ],
   alphaCSR[ 112 ][ 217 ],
   alphaCSR[ 112 ][ 218 ],
   alphaCSR[ 112 ][ 219 ],
   alphaCSR[ 112 ][ 220 ],
   alphaCSR[ 112 ][ 221 ],
   alphaCSR[ 112 ][ 222 ],
   alphaCSR[ 112 ][ 223 ],
   alphaCSR[ 112 ][ 224 ],
   alphaCSR[ 112 ][ 225 ],
   alphaCSR[ 112 ][ 226 ],
   alphaCSR[ 112 ][ 227 ],
   alphaCSR[ 112 ][ 228 ],
   alphaCSR[ 112 ][ 229 ],
   alphaCSR[ 112 ][ 230 ],
   alphaCSR[ 112 ][ 231 ],
   alphaCSR[ 112 ][ 232 ],
   alphaCSR[ 112 ][ 233 ],
   alphaCSR[ 112 ][ 234 ],
   alphaCSR[ 112 ][ 235 ],
   alphaCSR[ 112 ][ 236 ],
   alphaCSR[ 112 ][ 237 ],
   alphaCSR[ 112 ][ 238 ],
   alphaCSR[ 112 ][ 239 ],
   alphaCSR[ 112 ][ 240 ],
   alphaCSR[ 112 ][ 241 ],
   alphaCSR[ 112 ][ 242 ],
   alphaCSR[ 112 ][ 243 ],
   alphaCSR[ 112 ][ 244 ],
   alphaCSR[ 112 ][ 245 ],
   alphaCSR[ 112 ][ 246 ],
   alphaCSR[ 112 ][ 247 ],
   alphaCSR[ 112 ][ 248 ],
   alphaCSR[ 112 ][ 249 ],
   alphaCSR[ 112 ][ 250 ],
   alphaCSR[ 112 ][ 251 ],
   alphaCSR[ 112 ][ 252 ],
   alphaCSR[ 112 ][ 253 ],
   alphaCSR[ 112 ][ 254 ],
   alphaCSR[ 112 ][ 255 ],
   alphaCSR[ 112 ][ 256 ],
   alphaCSR[ 112 ][ 257 ],
   alphaCSR[ 112 ][ 258 ],
   alphaCSR[ 112 ][ 259 ],
   alphaCSR[ 112 ][ 260 ],
   alphaCSR[ 112 ][ 261 ],
   alphaCSR[ 112 ][ 262 ],
   alphaCSR[ 112 ][ 263 ],
   alphaCSR[ 112 ][ 264 ],
   alphaCSR[ 112 ][ 265 ],
   alphaCSR[ 112 ][ 266 ],
   alphaCSR[ 112 ][ 267 ],
   alphaCSR[ 112 ][ 268 ],
   alphaCSR[ 112 ][ 269 ],
   alphaCSR[ 112 ][ 270 ],
   alphaCSR[ 112 ][ 271 ],
   alphaCSR[ 112 ][ 272 ],
   alphaCSR[ 112 ][ 273 ],
   alphaCSR[ 112 ][ 274 ],
   alphaCSR[ 112 ][ 275 ],
   alphaCSR[ 112 ][ 276 ],
   alphaCSR[ 112 ][ 277 ],
   alphaCSR[ 112 ][ 278 ],
   alphaCSR[ 112 ][ 279 ],
   alphaCSR[ 112 ][ 280 ],
   alphaCSR[ 112 ][ 281 ],
   alphaCSR[ 112 ][ 282 ],
   alphaCSR[ 112 ][ 283 ],
   alphaCSR[ 112 ][ 284 ],
   alphaCSR[ 112 ][ 285 ],
   alphaCSR[ 112 ][ 286 ],
   alphaCSR[ 112 ][ 287 ],
   alphaCSR[ 112 ][ 288 ],
   alphaCSR[ 112 ][ 289 ],
   alphaCSR[ 112 ][ 290 ],
   alphaCSR[ 112 ][ 291 ],
   alphaCSR[ 112 ][ 292 ],
   alphaCSR[ 112 ][ 293 ],
   alphaCSR[ 112 ][ 294 ],
   alphaCSR[ 112 ][ 295 ],
   alphaCSR[ 112 ][ 296 ],
   alphaCSR[ 112 ][ 297 ],
   alphaCSR[ 112 ][ 298 ],
   alphaCSR[ 112 ][ 299 ],
   alphaCSR[ 112 ][ 300 ],
   alphaCSR[ 112 ][ 301 ],
   alphaCSR[ 112 ][ 302 ],
   alphaCSR[ 112 ][ 303 ],
   alphaCSR[ 112 ][ 304 ],
   alphaCSR[ 112 ][ 305 ],
   alphaCSR[ 112 ][ 306 ],
   alphaCSR[ 112 ][ 307 ],
   alphaCSR[ 112 ][ 308 ],
   alphaCSR[ 112 ][ 309 ],
   alphaCSR[ 112 ][ 310 ],
   alphaCSR[ 112 ][ 311 ],
   alphaCSR[ 112 ][ 312 ],
   alphaCSR[ 112 ][ 313 ],
   alphaCSR[ 112 ][ 314 ],
   alphaCSR[ 112 ][ 315 ],
   alphaCSR[ 112 ][ 316 ],
   alphaCSR[ 112 ][ 317 ],
   alphaCSR[ 112 ][ 318 ],
   alphaCSR[ 112 ][ 319 ],
   alphaCSR[ 112 ][ 320 ],
   alphaCSR[ 112 ][ 321 ],
   alphaCSR[ 112 ][ 322 ],
   alphaCSR[ 112 ][ 323 ],
   alphaCSR[ 112 ][ 324 ],
   alphaCSR[ 112 ][ 325 ],
   alphaCSR[ 112 ][ 326 ],
   alphaCSR[ 112 ][ 327 ],
   alphaCSR[ 112 ][ 328 ],
   alphaCSR[ 112 ][ 329 ],
   alphaCSR[ 112 ][ 330 ],
   alphaCSR[ 112 ][ 331 ],
   alphaCSR[ 112 ][ 332 ],
   alphaCSR[ 112 ][ 333 ],
   alphaCSR[ 112 ][ 334 ],
   alphaCSR[ 112 ][ 335 ],
   alphaCSR[ 112 ][ 336 ],
   alphaCSR[ 112 ][ 337 ],
   alphaCSR[ 112 ][ 338 ],
   alphaCSR[ 112 ][ 339 ],
   alphaCSR[ 112 ][ 340 ],
   alphaCSR[ 112 ][ 341 ],
   alphaCSR[ 112 ][ 342 ],
   alphaCSR[ 112 ][ 343 ],
   alphaCSR[ 112 ][ 344 ],
   alphaCSR[ 112 ][ 345 ],
   alphaCSR[ 112 ][ 346 ],
   alphaCSR[ 112 ][ 347 ],
   alphaCSR[ 112 ][ 348 ],
   alphaCSR[ 112 ][ 349 ],
   alphaCSR[ 112 ][ 350 ],
   alphaCSR[ 112 ][ 351 ],
   alphaCSR[ 112 ][ 352 ],
   alphaCSR[ 112 ][ 353 ],
   alphaCSR[ 112 ][ 354 ],
   alphaCSR[ 112 ][ 355 ],
   alphaCSR[ 112 ][ 356 ],
   alphaCSR[ 112 ][ 357 ],
   alphaCSR[ 112 ][ 358 ],
   alphaCSR[ 112 ][ 359 ],
   alphaCSR[ 112 ][ 360 ],
   alphaCSR[ 112 ][ 361 ],
   alphaCSR[ 112 ][ 362 ],
   alphaCSR[ 112 ][ 363 ],
   alphaCSR[ 112 ][ 364 ],
   alphaCSR[ 112 ][ 365 ],
   alphaCSR[ 112 ][ 366 ],
   alphaCSR[ 112 ][ 367 ],
   alphaCSR[ 112 ][ 368 ],
   alphaCSR[ 112 ][ 369 ],
   alphaCSR[ 112 ][ 370 ],
   alphaCSR[ 112 ][ 371 ],
   alphaCSR[ 112 ][ 372 ],
   alphaCSR[ 112 ][ 373 ],
   alphaCSR[ 112 ][ 374 ],
   alphaCSR[ 112 ][ 375 ],
   alphaCSR[ 112 ][ 376 ],
   alphaCSR[ 112 ][ 377 ],
   alphaCSR[ 112 ][ 378 ],
   alphaCSR[ 112 ][ 379 ],
   alphaCSR[ 112 ][ 380 ],
   alphaCSR[ 112 ][ 381 ],
   alphaCSR[ 112 ][ 382 ],
   alphaCSR[ 112 ][ 383 ],
   alphaCSR[ 113 ][ 0 ],
   alphaCSR[ 113 ][ 1 ],
   alphaCSR[ 113 ][ 2 ],
   alphaCSR[ 113 ][ 3 ],
   alphaCSR[ 113 ][ 4 ],
   alphaCSR[ 113 ][ 5 ],
   alphaCSR[ 113 ][ 6 ],
   alphaCSR[ 113 ][ 7 ],
   alphaCSR[ 113 ][ 8 ],
   alphaCSR[ 113 ][ 9 ],
   alphaCSR[ 113 ][ 10 ],
   alphaCSR[ 113 ][ 11 ],
   alphaCSR[ 113 ][ 12 ],
   alphaCSR[ 113 ][ 13 ],
   alphaCSR[ 113 ][ 14 ],
   alphaCSR[ 113 ][ 15 ],
   alphaCSR[ 113 ][ 16 ],
   alphaCSR[ 113 ][ 17 ],
   alphaCSR[ 113 ][ 18 ],
   alphaCSR[ 113 ][ 19 ],
   alphaCSR[ 113 ][ 20 ],
   alphaCSR[ 113 ][ 21 ],
   alphaCSR[ 113 ][ 22 ],
   alphaCSR[ 113 ][ 23 ],
   alphaCSR[ 113 ][ 24 ],
   alphaCSR[ 113 ][ 25 ],
   alphaCSR[ 113 ][ 26 ],
   alphaCSR[ 113 ][ 27 ],
   alphaCSR[ 113 ][ 28 ],
   alphaCSR[ 113 ][ 29 ],
   alphaCSR[ 113 ][ 30 ],
   alphaCSR[ 113 ][ 31 ],
   alphaCSR[ 113 ][ 32 ],
   alphaCSR[ 113 ][ 33 ],
   alphaCSR[ 113 ][ 34 ],
   alphaCSR[ 113 ][ 35 ],
   alphaCSR[ 113 ][ 36 ],
   alphaCSR[ 113 ][ 37 ],
   alphaCSR[ 113 ][ 38 ],
   alphaCSR[ 113 ][ 39 ],
   alphaCSR[ 113 ][ 40 ],
   alphaCSR[ 113 ][ 41 ],
   alphaCSR[ 113 ][ 42 ],
   alphaCSR[ 113 ][ 43 ],
   alphaCSR[ 113 ][ 44 ],
   alphaCSR[ 113 ][ 45 ],
   alphaCSR[ 113 ][ 46 ],
   alphaCSR[ 113 ][ 47 ],
   alphaCSR[ 113 ][ 48 ],
   alphaCSR[ 113 ][ 49 ],
   alphaCSR[ 113 ][ 50 ],
   alphaCSR[ 113 ][ 51 ],
   alphaCSR[ 113 ][ 52 ],
   alphaCSR[ 113 ][ 53 ],
   alphaCSR[ 113 ][ 54 ],
   alphaCSR[ 113 ][ 55 ],
   alphaCSR[ 113 ][ 56 ],
   alphaCSR[ 113 ][ 57 ],
   alphaCSR[ 113 ][ 58 ],
   alphaCSR[ 113 ][ 59 ],
   alphaCSR[ 113 ][ 60 ],
   alphaCSR[ 113 ][ 61 ],
   alphaCSR[ 113 ][ 62 ],
   alphaCSR[ 113 ][ 63 ],
   alphaCSR[ 113 ][ 64 ],
   alphaCSR[ 113 ][ 65 ],
   alphaCSR[ 113 ][ 66 ],
   alphaCSR[ 113 ][ 67 ],
   alphaCSR[ 113 ][ 68 ],
   alphaCSR[ 113 ][ 69 ],
   alphaCSR[ 113 ][ 70 ],
   alphaCSR[ 113 ][ 71 ],
   alphaCSR[ 113 ][ 72 ],
   alphaCSR[ 113 ][ 73 ],
   alphaCSR[ 113 ][ 74 ],
   alphaCSR[ 113 ][ 75 ],
   alphaCSR[ 113 ][ 76 ],
   alphaCSR[ 113 ][ 77 ],
   alphaCSR[ 113 ][ 78 ],
   alphaCSR[ 113 ][ 79 ],
   alphaCSR[ 113 ][ 80 ],
   alphaCSR[ 113 ][ 81 ],
   alphaCSR[ 113 ][ 82 ],
   alphaCSR[ 113 ][ 83 ],
   alphaCSR[ 113 ][ 84 ],
   alphaCSR[ 113 ][ 85 ],
   alphaCSR[ 113 ][ 86 ],
   alphaCSR[ 113 ][ 87 ],
   alphaCSR[ 113 ][ 88 ],
   alphaCSR[ 113 ][ 89 ],
   alphaCSR[ 113 ][ 90 ],
   alphaCSR[ 113 ][ 91 ],
   alphaCSR[ 113 ][ 92 ],
   alphaCSR[ 113 ][ 93 ],
   alphaCSR[ 113 ][ 94 ],
   alphaCSR[ 113 ][ 95 ],
   alphaCSR[ 113 ][ 96 ],
   alphaCSR[ 113 ][ 97 ],
   alphaCSR[ 113 ][ 98 ],
   alphaCSR[ 113 ][ 99 ],
   alphaCSR[ 113 ][ 100 ],
   alphaCSR[ 113 ][ 101 ],
   alphaCSR[ 113 ][ 102 ],
   alphaCSR[ 113 ][ 103 ],
   alphaCSR[ 113 ][ 104 ],
   alphaCSR[ 113 ][ 105 ],
   alphaCSR[ 113 ][ 106 ],
   alphaCSR[ 113 ][ 107 ],
   alphaCSR[ 113 ][ 108 ],
   alphaCSR[ 113 ][ 109 ],
   alphaCSR[ 113 ][ 110 ],
   alphaCSR[ 113 ][ 111 ],
   alphaCSR[ 113 ][ 112 ],
   alphaCSR[ 113 ][ 113 ],
   alphaCSR[ 113 ][ 114 ],
   alphaCSR[ 113 ][ 115 ],
   alphaCSR[ 113 ][ 116 ],
   alphaCSR[ 113 ][ 117 ],
   alphaCSR[ 113 ][ 118 ],
   alphaCSR[ 113 ][ 119 ],
   alphaCSR[ 113 ][ 120 ],
   alphaCSR[ 113 ][ 121 ],
   alphaCSR[ 113 ][ 122 ],
   alphaCSR[ 113 ][ 123 ],
   alphaCSR[ 113 ][ 124 ],
   alphaCSR[ 113 ][ 125 ],
   alphaCSR[ 113 ][ 126 ],
   alphaCSR[ 113 ][ 127 ],
   alphaCSR[ 113 ][ 128 ],
   alphaCSR[ 113 ][ 129 ],
   alphaCSR[ 113 ][ 130 ],
   alphaCSR[ 113 ][ 131 ],
   alphaCSR[ 113 ][ 132 ],
   alphaCSR[ 113 ][ 133 ],
   alphaCSR[ 113 ][ 134 ],
   alphaCSR[ 113 ][ 135 ],
   alphaCSR[ 113 ][ 136 ],
   alphaCSR[ 113 ][ 137 ],
   alphaCSR[ 113 ][ 138 ],
   alphaCSR[ 113 ][ 139 ],
   alphaCSR[ 113 ][ 140 ],
   alphaCSR[ 113 ][ 141 ],
   alphaCSR[ 113 ][ 142 ],
   alphaCSR[ 113 ][ 143 ],
   alphaCSR[ 113 ][ 144 ],
   alphaCSR[ 113 ][ 145 ],
   alphaCSR[ 113 ][ 146 ],
   alphaCSR[ 113 ][ 147 ],
   alphaCSR[ 113 ][ 148 ],
   alphaCSR[ 113 ][ 149 ],
   alphaCSR[ 113 ][ 150 ],
   alphaCSR[ 113 ][ 151 ],
   alphaCSR[ 113 ][ 152 ],
   alphaCSR[ 113 ][ 153 ],
   alphaCSR[ 113 ][ 154 ],
   alphaCSR[ 113 ][ 155 ],
   alphaCSR[ 113 ][ 156 ],
   alphaCSR[ 113 ][ 157 ],
   alphaCSR[ 113 ][ 158 ],
   alphaCSR[ 113 ][ 159 ],
   alphaCSR[ 113 ][ 160 ],
   alphaCSR[ 113 ][ 161 ],
   alphaCSR[ 113 ][ 162 ],
   alphaCSR[ 113 ][ 163 ],
   alphaCSR[ 113 ][ 164 ],
   alphaCSR[ 113 ][ 165 ],
   alphaCSR[ 113 ][ 166 ],
   alphaCSR[ 113 ][ 167 ],
   alphaCSR[ 113 ][ 168 ],
   alphaCSR[ 113 ][ 169 ],
   alphaCSR[ 113 ][ 170 ],
   alphaCSR[ 113 ][ 171 ],
   alphaCSR[ 113 ][ 172 ],
   alphaCSR[ 113 ][ 173 ],
   alphaCSR[ 113 ][ 174 ],
   alphaCSR[ 113 ][ 175 ],
   alphaCSR[ 113 ][ 176 ],
   alphaCSR[ 113 ][ 177 ],
   alphaCSR[ 113 ][ 178 ],
   alphaCSR[ 113 ][ 179 ],
   alphaCSR[ 113 ][ 180 ],
   alphaCSR[ 113 ][ 181 ],
   alphaCSR[ 113 ][ 182 ],
   alphaCSR[ 113 ][ 183 ],
   alphaCSR[ 113 ][ 184 ],
   alphaCSR[ 113 ][ 185 ],
   alphaCSR[ 113 ][ 186 ],
   alphaCSR[ 113 ][ 187 ],
   alphaCSR[ 113 ][ 188 ],
   alphaCSR[ 113 ][ 189 ],
   alphaCSR[ 113 ][ 190 ],
   alphaCSR[ 113 ][ 191 ],
   alphaCSR[ 113 ][ 192 ],
   alphaCSR[ 113 ][ 193 ],
   alphaCSR[ 113 ][ 194 ],
   alphaCSR[ 113 ][ 195 ],
   alphaCSR[ 113 ][ 196 ],
   alphaCSR[ 113 ][ 197 ],
   alphaCSR[ 113 ][ 198 ],
   alphaCSR[ 113 ][ 199 ],
   alphaCSR[ 113 ][ 200 ],
   alphaCSR[ 113 ][ 201 ],
   alphaCSR[ 113 ][ 202 ],
   alphaCSR[ 113 ][ 203 ],
   alphaCSR[ 113 ][ 204 ],
   alphaCSR[ 113 ][ 205 ],
   alphaCSR[ 113 ][ 206 ],
   alphaCSR[ 113 ][ 207 ],
   alphaCSR[ 113 ][ 208 ],
   alphaCSR[ 113 ][ 209 ],
   alphaCSR[ 113 ][ 210 ],
   alphaCSR[ 113 ][ 211 ],
   alphaCSR[ 113 ][ 212 ],
   alphaCSR[ 113 ][ 213 ],
   alphaCSR[ 113 ][ 214 ],
   alphaCSR[ 113 ][ 215 ],
   alphaCSR[ 113 ][ 216 ],
   alphaCSR[ 113 ][ 217 ],
   alphaCSR[ 113 ][ 218 ],
   alphaCSR[ 113 ][ 219 ],
   alphaCSR[ 113 ][ 220 ],
   alphaCSR[ 113 ][ 221 ],
   alphaCSR[ 113 ][ 222 ],
   alphaCSR[ 113 ][ 223 ],
   alphaCSR[ 113 ][ 224 ],
   alphaCSR[ 113 ][ 225 ],
   alphaCSR[ 113 ][ 226 ],
   alphaCSR[ 113 ][ 227 ],
   alphaCSR[ 113 ][ 228 ],
   alphaCSR[ 113 ][ 229 ],
   alphaCSR[ 113 ][ 230 ],
   alphaCSR[ 113 ][ 231 ],
   alphaCSR[ 113 ][ 232 ],
   alphaCSR[ 113 ][ 233 ],
   alphaCSR[ 113 ][ 234 ],
   alphaCSR[ 113 ][ 235 ],
   alphaCSR[ 113 ][ 236 ],
   alphaCSR[ 113 ][ 237 ],
   alphaCSR[ 113 ][ 238 ],
   alphaCSR[ 113 ][ 239 ],
   alphaCSR[ 113 ][ 240 ],
   alphaCSR[ 113 ][ 241 ],
   alphaCSR[ 113 ][ 242 ],
   alphaCSR[ 113 ][ 243 ],
   alphaCSR[ 113 ][ 244 ],
   alphaCSR[ 113 ][ 245 ],
   alphaCSR[ 113 ][ 246 ],
   alphaCSR[ 113 ][ 247 ],
   alphaCSR[ 113 ][ 248 ],
   alphaCSR[ 113 ][ 249 ],
   alphaCSR[ 113 ][ 250 ],
   alphaCSR[ 113 ][ 251 ],
   alphaCSR[ 113 ][ 252 ],
   alphaCSR[ 113 ][ 253 ],
   alphaCSR[ 113 ][ 254 ],
   alphaCSR[ 113 ][ 255 ],
   alphaCSR[ 113 ][ 256 ],
   alphaCSR[ 113 ][ 257 ],
   alphaCSR[ 113 ][ 258 ],
   alphaCSR[ 113 ][ 259 ],
   alphaCSR[ 113 ][ 260 ],
   alphaCSR[ 113 ][ 261 ],
   alphaCSR[ 113 ][ 262 ],
   alphaCSR[ 113 ][ 263 ],
   alphaCSR[ 113 ][ 264 ],
   alphaCSR[ 113 ][ 265 ],
   alphaCSR[ 113 ][ 266 ],
   alphaCSR[ 113 ][ 267 ],
   alphaCSR[ 113 ][ 268 ],
   alphaCSR[ 113 ][ 269 ],
   alphaCSR[ 113 ][ 270 ],
   alphaCSR[ 113 ][ 271 ],
   alphaCSR[ 113 ][ 272 ],
   alphaCSR[ 113 ][ 273 ],
   alphaCSR[ 113 ][ 274 ],
   alphaCSR[ 113 ][ 275 ],
   alphaCSR[ 113 ][ 276 ],
   alphaCSR[ 113 ][ 277 ],
   alphaCSR[ 113 ][ 278 ],
   alphaCSR[ 113 ][ 279 ],
   alphaCSR[ 113 ][ 280 ],
   alphaCSR[ 113 ][ 281 ],
   alphaCSR[ 113 ][ 282 ],
   alphaCSR[ 113 ][ 283 ],
   alphaCSR[ 113 ][ 284 ],
   alphaCSR[ 113 ][ 285 ],
   alphaCSR[ 113 ][ 286 ],
   alphaCSR[ 113 ][ 287 ],
   alphaCSR[ 113 ][ 288 ],
   alphaCSR[ 113 ][ 289 ],
   alphaCSR[ 113 ][ 290 ],
   alphaCSR[ 113 ][ 291 ],
   alphaCSR[ 113 ][ 292 ],
   alphaCSR[ 113 ][ 293 ],
   alphaCSR[ 113 ][ 294 ],
   alphaCSR[ 113 ][ 295 ],
   alphaCSR[ 113 ][ 296 ],
   alphaCSR[ 113 ][ 297 ],
   alphaCSR[ 113 ][ 298 ],
   alphaCSR[ 113 ][ 299 ],
   alphaCSR[ 113 ][ 300 ],
   alphaCSR[ 113 ][ 301 ],
   alphaCSR[ 113 ][ 302 ],
   alphaCSR[ 113 ][ 303 ],
   alphaCSR[ 113 ][ 304 ],
   alphaCSR[ 113 ][ 305 ],
   alphaCSR[ 113 ][ 306 ],
   alphaCSR[ 113 ][ 307 ],
   alphaCSR[ 113 ][ 308 ],
   alphaCSR[ 113 ][ 309 ],
   alphaCSR[ 113 ][ 310 ],
   alphaCSR[ 113 ][ 311 ],
   alphaCSR[ 113 ][ 312 ],
   alphaCSR[ 113 ][ 313 ],
   alphaCSR[ 113 ][ 314 ],
   alphaCSR[ 113 ][ 315 ],
   alphaCSR[ 113 ][ 316 ],
   alphaCSR[ 113 ][ 317 ],
   alphaCSR[ 113 ][ 318 ],
   alphaCSR[ 113 ][ 319 ],
   alphaCSR[ 113 ][ 320 ],
   alphaCSR[ 113 ][ 321 ],
   alphaCSR[ 113 ][ 322 ],
   alphaCSR[ 113 ][ 323 ],
   alphaCSR[ 113 ][ 324 ],
   alphaCSR[ 113 ][ 325 ],
   alphaCSR[ 113 ][ 326 ],
   alphaCSR[ 113 ][ 327 ],
   alphaCSR[ 113 ][ 328 ],
   alphaCSR[ 113 ][ 329 ],
   alphaCSR[ 113 ][ 330 ],
   alphaCSR[ 113 ][ 331 ],
   alphaCSR[ 113 ][ 332 ],
   alphaCSR[ 113 ][ 333 ],
   alphaCSR[ 113 ][ 334 ],
   alphaCSR[ 113 ][ 335 ],
   alphaCSR[ 113 ][ 336 ],
   alphaCSR[ 113 ][ 337 ],
   alphaCSR[ 113 ][ 338 ],
   alphaCSR[ 113 ][ 339 ],
   alphaCSR[ 113 ][ 340 ],
   alphaCSR[ 113 ][ 341 ],
   alphaCSR[ 113 ][ 342 ],
   alphaCSR[ 113 ][ 343 ],
   alphaCSR[ 113 ][ 344 ],
   alphaCSR[ 113 ][ 345 ],
   alphaCSR[ 113 ][ 346 ],
   alphaCSR[ 113 ][ 347 ],
   alphaCSR[ 113 ][ 348 ],
   alphaCSR[ 113 ][ 349 ],
   alphaCSR[ 113 ][ 350 ],
   alphaCSR[ 113 ][ 351 ],
   alphaCSR[ 113 ][ 352 ],
   alphaCSR[ 113 ][ 353 ],
   alphaCSR[ 113 ][ 354 ],
   alphaCSR[ 113 ][ 355 ],
   alphaCSR[ 113 ][ 356 ],
   alphaCSR[ 113 ][ 357 ],
   alphaCSR[ 113 ][ 358 ],
   alphaCSR[ 113 ][ 359 ],
   alphaCSR[ 113 ][ 360 ],
   alphaCSR[ 113 ][ 361 ],
   alphaCSR[ 113 ][ 362 ],
   alphaCSR[ 113 ][ 363 ],
   alphaCSR[ 113 ][ 364 ],
   alphaCSR[ 113 ][ 365 ],
   alphaCSR[ 113 ][ 366 ],
   alphaCSR[ 113 ][ 367 ],
   alphaCSR[ 113 ][ 368 ],
   alphaCSR[ 113 ][ 369 ],
   alphaCSR[ 113 ][ 370 ],
   alphaCSR[ 113 ][ 371 ],
   alphaCSR[ 113 ][ 372 ],
   alphaCSR[ 113 ][ 373 ],
   alphaCSR[ 113 ][ 374 ],
   alphaCSR[ 113 ][ 375 ],
   alphaCSR[ 113 ][ 376 ],
   alphaCSR[ 113 ][ 377 ],
   alphaCSR[ 113 ][ 378 ],
   alphaCSR[ 113 ][ 379 ],
   alphaCSR[ 113 ][ 380 ],
   alphaCSR[ 113 ][ 381 ],
   alphaCSR[ 113 ][ 382 ],
   alphaCSR[ 113 ][ 383 ],
   alphaCSR[ 114 ][ 0 ],
   alphaCSR[ 114 ][ 1 ],
   alphaCSR[ 114 ][ 2 ],
   alphaCSR[ 114 ][ 3 ],
   alphaCSR[ 114 ][ 4 ],
   alphaCSR[ 114 ][ 5 ],
   alphaCSR[ 114 ][ 6 ],
   alphaCSR[ 114 ][ 7 ],
   alphaCSR[ 114 ][ 8 ],
   alphaCSR[ 114 ][ 9 ],
   alphaCSR[ 114 ][ 10 ],
   alphaCSR[ 114 ][ 11 ],
   alphaCSR[ 114 ][ 12 ],
   alphaCSR[ 114 ][ 13 ],
   alphaCSR[ 114 ][ 14 ],
   alphaCSR[ 114 ][ 15 ],
   alphaCSR[ 114 ][ 16 ],
   alphaCSR[ 114 ][ 17 ],
   alphaCSR[ 114 ][ 18 ],
   alphaCSR[ 114 ][ 19 ],
   alphaCSR[ 114 ][ 20 ],
   alphaCSR[ 114 ][ 21 ],
   alphaCSR[ 114 ][ 22 ],
   alphaCSR[ 114 ][ 23 ],
   alphaCSR[ 114 ][ 24 ],
   alphaCSR[ 114 ][ 25 ],
   alphaCSR[ 114 ][ 26 ],
   alphaCSR[ 114 ][ 27 ],
   alphaCSR[ 114 ][ 28 ],
   alphaCSR[ 114 ][ 29 ],
   alphaCSR[ 114 ][ 30 ],
   alphaCSR[ 114 ][ 31 ],
   alphaCSR[ 114 ][ 32 ],
   alphaCSR[ 114 ][ 33 ],
   alphaCSR[ 114 ][ 34 ],
   alphaCSR[ 114 ][ 35 ],
   alphaCSR[ 114 ][ 36 ],
   alphaCSR[ 114 ][ 37 ],
   alphaCSR[ 114 ][ 38 ],
   alphaCSR[ 114 ][ 39 ],
   alphaCSR[ 114 ][ 40 ],
   alphaCSR[ 114 ][ 41 ],
   alphaCSR[ 114 ][ 42 ],
   alphaCSR[ 114 ][ 43 ],
   alphaCSR[ 114 ][ 44 ],
   alphaCSR[ 114 ][ 45 ],
   alphaCSR[ 114 ][ 46 ],
   alphaCSR[ 114 ][ 47 ],
   alphaCSR[ 114 ][ 48 ],
   alphaCSR[ 114 ][ 49 ],
   alphaCSR[ 114 ][ 50 ],
   alphaCSR[ 114 ][ 51 ],
   alphaCSR[ 114 ][ 52 ],
   alphaCSR[ 114 ][ 53 ],
   alphaCSR[ 114 ][ 54 ],
   alphaCSR[ 114 ][ 55 ],
   alphaCSR[ 114 ][ 56 ],
   alphaCSR[ 114 ][ 57 ],
   alphaCSR[ 114 ][ 58 ],
   alphaCSR[ 114 ][ 59 ],
   alphaCSR[ 114 ][ 60 ],
   alphaCSR[ 114 ][ 61 ],
   alphaCSR[ 114 ][ 62 ],
   alphaCSR[ 114 ][ 63 ],
   alphaCSR[ 114 ][ 64 ],
   alphaCSR[ 114 ][ 65 ],
   alphaCSR[ 114 ][ 66 ],
   alphaCSR[ 114 ][ 67 ],
   alphaCSR[ 114 ][ 68 ],
   alphaCSR[ 114 ][ 69 ],
   alphaCSR[ 114 ][ 70 ],
   alphaCSR[ 114 ][ 71 ],
   alphaCSR[ 114 ][ 72 ],
   alphaCSR[ 114 ][ 73 ],
   alphaCSR[ 114 ][ 74 ],
   alphaCSR[ 114 ][ 75 ],
   alphaCSR[ 114 ][ 76 ],
   alphaCSR[ 114 ][ 77 ],
   alphaCSR[ 114 ][ 78 ],
   alphaCSR[ 114 ][ 79 ],
   alphaCSR[ 114 ][ 80 ],
   alphaCSR[ 114 ][ 81 ],
   alphaCSR[ 114 ][ 82 ],
   alphaCSR[ 114 ][ 83 ],
   alphaCSR[ 114 ][ 84 ],
   alphaCSR[ 114 ][ 85 ],
   alphaCSR[ 114 ][ 86 ],
   alphaCSR[ 114 ][ 87 ],
   alphaCSR[ 114 ][ 88 ],
   alphaCSR[ 114 ][ 89 ],
   alphaCSR[ 114 ][ 90 ],
   alphaCSR[ 114 ][ 91 ],
   alphaCSR[ 114 ][ 92 ],
   alphaCSR[ 114 ][ 93 ],
   alphaCSR[ 114 ][ 94 ],
   alphaCSR[ 114 ][ 95 ],
   alphaCSR[ 114 ][ 96 ],
   alphaCSR[ 114 ][ 97 ],
   alphaCSR[ 114 ][ 98 ],
   alphaCSR[ 114 ][ 99 ],
   alphaCSR[ 114 ][ 100 ],
   alphaCSR[ 114 ][ 101 ],
   alphaCSR[ 114 ][ 102 ],
   alphaCSR[ 114 ][ 103 ],
   alphaCSR[ 114 ][ 104 ],
   alphaCSR[ 114 ][ 105 ],
   alphaCSR[ 114 ][ 106 ],
   alphaCSR[ 114 ][ 107 ],
   alphaCSR[ 114 ][ 108 ],
   alphaCSR[ 114 ][ 109 ],
   alphaCSR[ 114 ][ 110 ],
   alphaCSR[ 114 ][ 111 ],
   alphaCSR[ 114 ][ 112 ],
   alphaCSR[ 114 ][ 113 ],
   alphaCSR[ 114 ][ 114 ],
   alphaCSR[ 114 ][ 115 ],
   alphaCSR[ 114 ][ 116 ],
   alphaCSR[ 114 ][ 117 ],
   alphaCSR[ 114 ][ 118 ],
   alphaCSR[ 114 ][ 119 ],
   alphaCSR[ 114 ][ 120 ],
   alphaCSR[ 114 ][ 121 ],
   alphaCSR[ 114 ][ 122 ],
   alphaCSR[ 114 ][ 123 ],
   alphaCSR[ 114 ][ 124 ],
   alphaCSR[ 114 ][ 125 ],
   alphaCSR[ 114 ][ 126 ],
   alphaCSR[ 114 ][ 127 ],
   alphaCSR[ 114 ][ 128 ],
   alphaCSR[ 114 ][ 129 ],
   alphaCSR[ 114 ][ 130 ],
   alphaCSR[ 114 ][ 131 ],
   alphaCSR[ 114 ][ 132 ],
   alphaCSR[ 114 ][ 133 ],
   alphaCSR[ 114 ][ 134 ],
   alphaCSR[ 114 ][ 135 ],
   alphaCSR[ 114 ][ 136 ],
   alphaCSR[ 114 ][ 137 ],
   alphaCSR[ 114 ][ 138 ],
   alphaCSR[ 114 ][ 139 ],
   alphaCSR[ 114 ][ 140 ],
   alphaCSR[ 114 ][ 141 ],
   alphaCSR[ 114 ][ 142 ],
   alphaCSR[ 114 ][ 143 ],
   alphaCSR[ 114 ][ 144 ],
   alphaCSR[ 114 ][ 145 ],
   alphaCSR[ 114 ][ 146 ],
   alphaCSR[ 114 ][ 147 ],
   alphaCSR[ 114 ][ 148 ],
   alphaCSR[ 114 ][ 149 ],
   alphaCSR[ 114 ][ 150 ],
   alphaCSR[ 114 ][ 151 ],
   alphaCSR[ 114 ][ 152 ],
   alphaCSR[ 114 ][ 153 ],
   alphaCSR[ 114 ][ 154 ],
   alphaCSR[ 114 ][ 155 ],
   alphaCSR[ 114 ][ 156 ],
   alphaCSR[ 114 ][ 157 ],
   alphaCSR[ 114 ][ 158 ],
   alphaCSR[ 114 ][ 159 ],
   alphaCSR[ 114 ][ 160 ],
   alphaCSR[ 114 ][ 161 ],
   alphaCSR[ 114 ][ 162 ],
   alphaCSR[ 114 ][ 163 ],
   alphaCSR[ 114 ][ 164 ],
   alphaCSR[ 114 ][ 165 ],
   alphaCSR[ 114 ][ 166 ],
   alphaCSR[ 114 ][ 167 ],
   alphaCSR[ 114 ][ 168 ],
   alphaCSR[ 114 ][ 169 ],
   alphaCSR[ 114 ][ 170 ],
   alphaCSR[ 114 ][ 171 ],
   alphaCSR[ 114 ][ 172 ],
   alphaCSR[ 114 ][ 173 ],
   alphaCSR[ 114 ][ 174 ],
   alphaCSR[ 114 ][ 175 ],
   alphaCSR[ 114 ][ 176 ],
   alphaCSR[ 114 ][ 177 ],
   alphaCSR[ 114 ][ 178 ],
   alphaCSR[ 114 ][ 179 ],
   alphaCSR[ 114 ][ 180 ],
   alphaCSR[ 114 ][ 181 ],
   alphaCSR[ 114 ][ 182 ],
   alphaCSR[ 114 ][ 183 ],
   alphaCSR[ 114 ][ 184 ],
   alphaCSR[ 114 ][ 185 ],
   alphaCSR[ 114 ][ 186 ],
   alphaCSR[ 114 ][ 187 ],
   alphaCSR[ 114 ][ 188 ],
   alphaCSR[ 114 ][ 189 ],
   alphaCSR[ 114 ][ 190 ],
   alphaCSR[ 114 ][ 191 ],
   alphaCSR[ 114 ][ 192 ],
   alphaCSR[ 114 ][ 193 ],
   alphaCSR[ 114 ][ 194 ],
   alphaCSR[ 114 ][ 195 ],
   alphaCSR[ 114 ][ 196 ],
   alphaCSR[ 114 ][ 197 ],
   alphaCSR[ 114 ][ 198 ],
   alphaCSR[ 114 ][ 199 ],
   alphaCSR[ 114 ][ 200 ],
   alphaCSR[ 114 ][ 201 ],
   alphaCSR[ 114 ][ 202 ],
   alphaCSR[ 114 ][ 203 ],
   alphaCSR[ 114 ][ 204 ],
   alphaCSR[ 114 ][ 205 ],
   alphaCSR[ 114 ][ 206 ],
   alphaCSR[ 114 ][ 207 ],
   alphaCSR[ 114 ][ 208 ],
   alphaCSR[ 114 ][ 209 ],
   alphaCSR[ 114 ][ 210 ],
   alphaCSR[ 114 ][ 211 ],
   alphaCSR[ 114 ][ 212 ],
   alphaCSR[ 114 ][ 213 ],
   alphaCSR[ 114 ][ 214 ],
   alphaCSR[ 114 ][ 215 ],
   alphaCSR[ 114 ][ 216 ],
   alphaCSR[ 114 ][ 217 ],
   alphaCSR[ 114 ][ 218 ],
   alphaCSR[ 114 ][ 219 ],
   alphaCSR[ 114 ][ 220 ],
   alphaCSR[ 114 ][ 221 ],
   alphaCSR[ 114 ][ 222 ],
   alphaCSR[ 114 ][ 223 ],
   alphaCSR[ 114 ][ 224 ],
   alphaCSR[ 114 ][ 225 ],
   alphaCSR[ 114 ][ 226 ],
   alphaCSR[ 114 ][ 227 ],
   alphaCSR[ 114 ][ 228 ],
   alphaCSR[ 114 ][ 229 ],
   alphaCSR[ 114 ][ 230 ],
   alphaCSR[ 114 ][ 231 ],
   alphaCSR[ 114 ][ 232 ],
   alphaCSR[ 114 ][ 233 ],
   alphaCSR[ 114 ][ 234 ],
   alphaCSR[ 114 ][ 235 ],
   alphaCSR[ 114 ][ 236 ],
   alphaCSR[ 114 ][ 237 ],
   alphaCSR[ 114 ][ 238 ],
   alphaCSR[ 114 ][ 239 ],
   alphaCSR[ 114 ][ 240 ],
   alphaCSR[ 114 ][ 241 ],
   alphaCSR[ 114 ][ 242 ],
   alphaCSR[ 114 ][ 243 ],
   alphaCSR[ 114 ][ 244 ],
   alphaCSR[ 114 ][ 245 ],
   alphaCSR[ 114 ][ 246 ],
   alphaCSR[ 114 ][ 247 ],
   alphaCSR[ 114 ][ 248 ],
   alphaCSR[ 114 ][ 249 ],
   alphaCSR[ 114 ][ 250 ],
   alphaCSR[ 114 ][ 251 ],
   alphaCSR[ 114 ][ 252 ],
   alphaCSR[ 114 ][ 253 ],
   alphaCSR[ 114 ][ 254 ],
   alphaCSR[ 114 ][ 255 ],
   alphaCSR[ 114 ][ 256 ],
   alphaCSR[ 114 ][ 257 ],
   alphaCSR[ 114 ][ 258 ],
   alphaCSR[ 114 ][ 259 ],
   alphaCSR[ 114 ][ 260 ],
   alphaCSR[ 114 ][ 261 ],
   alphaCSR[ 114 ][ 262 ],
   alphaCSR[ 114 ][ 263 ],
   alphaCSR[ 114 ][ 264 ],
   alphaCSR[ 114 ][ 265 ],
   alphaCSR[ 114 ][ 266 ],
   alphaCSR[ 114 ][ 267 ],
   alphaCSR[ 114 ][ 268 ],
   alphaCSR[ 114 ][ 269 ],
   alphaCSR[ 114 ][ 270 ],
   alphaCSR[ 114 ][ 271 ],
   alphaCSR[ 114 ][ 272 ],
   alphaCSR[ 114 ][ 273 ],
   alphaCSR[ 114 ][ 274 ],
   alphaCSR[ 114 ][ 275 ],
   alphaCSR[ 114 ][ 276 ],
   alphaCSR[ 114 ][ 277 ],
   alphaCSR[ 114 ][ 278 ],
   alphaCSR[ 114 ][ 279 ],
   alphaCSR[ 114 ][ 280 ],
   alphaCSR[ 114 ][ 281 ],
   alphaCSR[ 114 ][ 282 ],
   alphaCSR[ 114 ][ 283 ],
   alphaCSR[ 114 ][ 284 ],
   alphaCSR[ 114 ][ 285 ],
   alphaCSR[ 114 ][ 286 ],
   alphaCSR[ 114 ][ 287 ],
   alphaCSR[ 114 ][ 288 ],
   alphaCSR[ 114 ][ 289 ],
   alphaCSR[ 114 ][ 290 ],
   alphaCSR[ 114 ][ 291 ],
   alphaCSR[ 114 ][ 292 ],
   alphaCSR[ 114 ][ 293 ],
   alphaCSR[ 114 ][ 294 ],
   alphaCSR[ 114 ][ 295 ],
   alphaCSR[ 114 ][ 296 ],
   alphaCSR[ 114 ][ 297 ],
   alphaCSR[ 114 ][ 298 ],
   alphaCSR[ 114 ][ 299 ],
   alphaCSR[ 114 ][ 300 ],
   alphaCSR[ 114 ][ 301 ],
   alphaCSR[ 114 ][ 302 ],
   alphaCSR[ 114 ][ 303 ],
   alphaCSR[ 114 ][ 304 ],
   alphaCSR[ 114 ][ 305 ],
   alphaCSR[ 114 ][ 306 ],
   alphaCSR[ 114 ][ 307 ],
   alphaCSR[ 114 ][ 308 ],
   alphaCSR[ 114 ][ 309 ],
   alphaCSR[ 114 ][ 310 ],
   alphaCSR[ 114 ][ 311 ],
   alphaCSR[ 114 ][ 312 ],
   alphaCSR[ 114 ][ 313 ],
   alphaCSR[ 114 ][ 314 ],
   alphaCSR[ 114 ][ 315 ],
   alphaCSR[ 114 ][ 316 ],
   alphaCSR[ 114 ][ 317 ],
   alphaCSR[ 114 ][ 318 ],
   alphaCSR[ 114 ][ 319 ],
   alphaCSR[ 114 ][ 320 ],
   alphaCSR[ 114 ][ 321 ],
   alphaCSR[ 114 ][ 322 ],
   alphaCSR[ 114 ][ 323 ],
   alphaCSR[ 114 ][ 324 ],
   alphaCSR[ 114 ][ 325 ],
   alphaCSR[ 114 ][ 326 ],
   alphaCSR[ 114 ][ 327 ],
   alphaCSR[ 114 ][ 328 ],
   alphaCSR[ 114 ][ 329 ],
   alphaCSR[ 114 ][ 330 ],
   alphaCSR[ 114 ][ 331 ],
   alphaCSR[ 114 ][ 332 ],
   alphaCSR[ 114 ][ 333 ],
   alphaCSR[ 114 ][ 334 ],
   alphaCSR[ 114 ][ 335 ],
   alphaCSR[ 114 ][ 336 ],
   alphaCSR[ 114 ][ 337 ],
   alphaCSR[ 114 ][ 338 ],
   alphaCSR[ 114 ][ 339 ],
   alphaCSR[ 114 ][ 340 ],
   alphaCSR[ 114 ][ 341 ],
   alphaCSR[ 114 ][ 342 ],
   alphaCSR[ 114 ][ 343 ],
   alphaCSR[ 114 ][ 344 ],
   alphaCSR[ 114 ][ 345 ],
   alphaCSR[ 114 ][ 346 ],
   alphaCSR[ 114 ][ 347 ],
   alphaCSR[ 114 ][ 348 ],
   alphaCSR[ 114 ][ 349 ],
   alphaCSR[ 114 ][ 350 ],
   alphaCSR[ 114 ][ 351 ],
   alphaCSR[ 114 ][ 352 ],
   alphaCSR[ 114 ][ 353 ],
   alphaCSR[ 114 ][ 354 ],
   alphaCSR[ 114 ][ 355 ],
   alphaCSR[ 114 ][ 356 ],
   alphaCSR[ 114 ][ 357 ],
   alphaCSR[ 114 ][ 358 ],
   alphaCSR[ 114 ][ 359 ],
   alphaCSR[ 114 ][ 360 ],
   alphaCSR[ 114 ][ 361 ],
   alphaCSR[ 114 ][ 362 ],
   alphaCSR[ 114 ][ 363 ],
   alphaCSR[ 114 ][ 364 ],
   alphaCSR[ 114 ][ 365 ],
   alphaCSR[ 114 ][ 366 ],
   alphaCSR[ 114 ][ 367 ],
   alphaCSR[ 114 ][ 368 ],
   alphaCSR[ 114 ][ 369 ],
   alphaCSR[ 114 ][ 370 ],
   alphaCSR[ 114 ][ 371 ],
   alphaCSR[ 114 ][ 372 ],
   alphaCSR[ 114 ][ 373 ],
   alphaCSR[ 114 ][ 374 ],
   alphaCSR[ 114 ][ 375 ],
   alphaCSR[ 114 ][ 376 ],
   alphaCSR[ 114 ][ 377 ],
   alphaCSR[ 114 ][ 378 ],
   alphaCSR[ 114 ][ 379 ],
   alphaCSR[ 114 ][ 380 ],
   alphaCSR[ 114 ][ 381 ],
   alphaCSR[ 114 ][ 382 ],
   alphaCSR[ 114 ][ 383 ],
   alphaCSR[ 115 ][ 0 ],
   alphaCSR[ 115 ][ 1 ],
   alphaCSR[ 115 ][ 2 ],
   alphaCSR[ 115 ][ 3 ],
   alphaCSR[ 115 ][ 4 ],
   alphaCSR[ 115 ][ 5 ],
   alphaCSR[ 115 ][ 6 ],
   alphaCSR[ 115 ][ 7 ],
   alphaCSR[ 115 ][ 8 ],
   alphaCSR[ 115 ][ 9 ],
   alphaCSR[ 115 ][ 10 ],
   alphaCSR[ 115 ][ 11 ],
   alphaCSR[ 115 ][ 12 ],
   alphaCSR[ 115 ][ 13 ],
   alphaCSR[ 115 ][ 14 ],
   alphaCSR[ 115 ][ 15 ],
   alphaCSR[ 115 ][ 16 ],
   alphaCSR[ 115 ][ 17 ],
   alphaCSR[ 115 ][ 18 ],
   alphaCSR[ 115 ][ 19 ],
   alphaCSR[ 115 ][ 20 ],
   alphaCSR[ 115 ][ 21 ],
   alphaCSR[ 115 ][ 22 ],
   alphaCSR[ 115 ][ 23 ],
   alphaCSR[ 115 ][ 24 ],
   alphaCSR[ 115 ][ 25 ],
   alphaCSR[ 115 ][ 26 ],
   alphaCSR[ 115 ][ 27 ],
   alphaCSR[ 115 ][ 28 ],
   alphaCSR[ 115 ][ 29 ],
   alphaCSR[ 115 ][ 30 ],
   alphaCSR[ 115 ][ 31 ],
   alphaCSR[ 115 ][ 32 ],
   alphaCSR[ 115 ][ 33 ],
   alphaCSR[ 115 ][ 34 ],
   alphaCSR[ 115 ][ 35 ],
   alphaCSR[ 115 ][ 36 ],
   alphaCSR[ 115 ][ 37 ],
   alphaCSR[ 115 ][ 38 ],
   alphaCSR[ 115 ][ 39 ],
   alphaCSR[ 115 ][ 40 ],
   alphaCSR[ 115 ][ 41 ],
   alphaCSR[ 115 ][ 42 ],
   alphaCSR[ 115 ][ 43 ],
   alphaCSR[ 115 ][ 44 ],
   alphaCSR[ 115 ][ 45 ],
   alphaCSR[ 115 ][ 46 ],
   alphaCSR[ 115 ][ 47 ],
   alphaCSR[ 115 ][ 48 ],
   alphaCSR[ 115 ][ 49 ],
   alphaCSR[ 115 ][ 50 ],
   alphaCSR[ 115 ][ 51 ],
   alphaCSR[ 115 ][ 52 ],
   alphaCSR[ 115 ][ 53 ],
   alphaCSR[ 115 ][ 54 ],
   alphaCSR[ 115 ][ 55 ],
   alphaCSR[ 115 ][ 56 ],
   alphaCSR[ 115 ][ 57 ],
   alphaCSR[ 115 ][ 58 ],
   alphaCSR[ 115 ][ 59 ],
   alphaCSR[ 115 ][ 60 ],
   alphaCSR[ 115 ][ 61 ],
   alphaCSR[ 115 ][ 62 ],
   alphaCSR[ 115 ][ 63 ],
   alphaCSR[ 115 ][ 64 ],
   alphaCSR[ 115 ][ 65 ],
   alphaCSR[ 115 ][ 66 ],
   alphaCSR[ 115 ][ 67 ],
   alphaCSR[ 115 ][ 68 ],
   alphaCSR[ 115 ][ 69 ],
   alphaCSR[ 115 ][ 70 ],
   alphaCSR[ 115 ][ 71 ],
   alphaCSR[ 115 ][ 72 ],
   alphaCSR[ 115 ][ 73 ],
   alphaCSR[ 115 ][ 74 ],
   alphaCSR[ 115 ][ 75 ],
   alphaCSR[ 115 ][ 76 ],
   alphaCSR[ 115 ][ 77 ],
   alphaCSR[ 115 ][ 78 ],
   alphaCSR[ 115 ][ 79 ],
   alphaCSR[ 115 ][ 80 ],
   alphaCSR[ 115 ][ 81 ],
   alphaCSR[ 115 ][ 82 ],
   alphaCSR[ 115 ][ 83 ],
   alphaCSR[ 115 ][ 84 ],
   alphaCSR[ 115 ][ 85 ],
   alphaCSR[ 115 ][ 86 ],
   alphaCSR[ 115 ][ 87 ],
   alphaCSR[ 115 ][ 88 ],
   alphaCSR[ 115 ][ 89 ],
   alphaCSR[ 115 ][ 90 ],
   alphaCSR[ 115 ][ 91 ],
   alphaCSR[ 115 ][ 92 ],
   alphaCSR[ 115 ][ 93 ],
   alphaCSR[ 115 ][ 94 ],
   alphaCSR[ 115 ][ 95 ],
   alphaCSR[ 115 ][ 96 ],
   alphaCSR[ 115 ][ 97 ],
   alphaCSR[ 115 ][ 98 ],
   alphaCSR[ 115 ][ 99 ],
   alphaCSR[ 115 ][ 100 ],
   alphaCSR[ 115 ][ 101 ],
   alphaCSR[ 115 ][ 102 ],
   alphaCSR[ 115 ][ 103 ],
   alphaCSR[ 115 ][ 104 ],
   alphaCSR[ 115 ][ 105 ],
   alphaCSR[ 115 ][ 106 ],
   alphaCSR[ 115 ][ 107 ],
   alphaCSR[ 115 ][ 108 ],
   alphaCSR[ 115 ][ 109 ],
   alphaCSR[ 115 ][ 110 ],
   alphaCSR[ 115 ][ 111 ],
   alphaCSR[ 115 ][ 112 ],
   alphaCSR[ 115 ][ 113 ],
   alphaCSR[ 115 ][ 114 ],
   alphaCSR[ 115 ][ 115 ],
   alphaCSR[ 115 ][ 116 ],
   alphaCSR[ 115 ][ 117 ],
   alphaCSR[ 115 ][ 118 ],
   alphaCSR[ 115 ][ 119 ],
   alphaCSR[ 115 ][ 120 ],
   alphaCSR[ 115 ][ 121 ],
   alphaCSR[ 115 ][ 122 ],
   alphaCSR[ 115 ][ 123 ],
   alphaCSR[ 115 ][ 124 ],
   alphaCSR[ 115 ][ 125 ],
   alphaCSR[ 115 ][ 126 ],
   alphaCSR[ 115 ][ 127 ],
   alphaCSR[ 115 ][ 128 ],
   alphaCSR[ 115 ][ 129 ],
   alphaCSR[ 115 ][ 130 ],
   alphaCSR[ 115 ][ 131 ],
   alphaCSR[ 115 ][ 132 ],
   alphaCSR[ 115 ][ 133 ],
   alphaCSR[ 115 ][ 134 ],
   alphaCSR[ 115 ][ 135 ],
   alphaCSR[ 115 ][ 136 ],
   alphaCSR[ 115 ][ 137 ],
   alphaCSR[ 115 ][ 138 ],
   alphaCSR[ 115 ][ 139 ],
   alphaCSR[ 115 ][ 140 ],
   alphaCSR[ 115 ][ 141 ],
   alphaCSR[ 115 ][ 142 ],
   alphaCSR[ 115 ][ 143 ],
   alphaCSR[ 115 ][ 144 ],
   alphaCSR[ 115 ][ 145 ],
   alphaCSR[ 115 ][ 146 ],
   alphaCSR[ 115 ][ 147 ],
   alphaCSR[ 115 ][ 148 ],
   alphaCSR[ 115 ][ 149 ],
   alphaCSR[ 115 ][ 150 ],
   alphaCSR[ 115 ][ 151 ],
   alphaCSR[ 115 ][ 152 ],
   alphaCSR[ 115 ][ 153 ],
   alphaCSR[ 115 ][ 154 ],
   alphaCSR[ 115 ][ 155 ],
   alphaCSR[ 115 ][ 156 ],
   alphaCSR[ 115 ][ 157 ],
   alphaCSR[ 115 ][ 158 ],
   alphaCSR[ 115 ][ 159 ],
   alphaCSR[ 115 ][ 160 ],
   alphaCSR[ 115 ][ 161 ],
   alphaCSR[ 115 ][ 162 ],
   alphaCSR[ 115 ][ 163 ],
   alphaCSR[ 115 ][ 164 ],
   alphaCSR[ 115 ][ 165 ],
   alphaCSR[ 115 ][ 166 ],
   alphaCSR[ 115 ][ 167 ],
   alphaCSR[ 115 ][ 168 ],
   alphaCSR[ 115 ][ 169 ],
   alphaCSR[ 115 ][ 170 ],
   alphaCSR[ 115 ][ 171 ],
   alphaCSR[ 115 ][ 172 ],
   alphaCSR[ 115 ][ 173 ],
   alphaCSR[ 115 ][ 174 ],
   alphaCSR[ 115 ][ 175 ],
   alphaCSR[ 115 ][ 176 ],
   alphaCSR[ 115 ][ 177 ],
   alphaCSR[ 115 ][ 178 ],
   alphaCSR[ 115 ][ 179 ],
   alphaCSR[ 115 ][ 180 ],
   alphaCSR[ 115 ][ 181 ],
   alphaCSR[ 115 ][ 182 ],
   alphaCSR[ 115 ][ 183 ],
   alphaCSR[ 115 ][ 184 ],
   alphaCSR[ 115 ][ 185 ],
   alphaCSR[ 115 ][ 186 ],
   alphaCSR[ 115 ][ 187 ],
   alphaCSR[ 115 ][ 188 ],
   alphaCSR[ 115 ][ 189 ],
   alphaCSR[ 115 ][ 190 ],
   alphaCSR[ 115 ][ 191 ],
   alphaCSR[ 115 ][ 192 ],
   alphaCSR[ 115 ][ 193 ],
   alphaCSR[ 115 ][ 194 ],
   alphaCSR[ 115 ][ 195 ],
   alphaCSR[ 115 ][ 196 ],
   alphaCSR[ 115 ][ 197 ],
   alphaCSR[ 115 ][ 198 ],
   alphaCSR[ 115 ][ 199 ],
   alphaCSR[ 115 ][ 200 ],
   alphaCSR[ 115 ][ 201 ],
   alphaCSR[ 115 ][ 202 ],
   alphaCSR[ 115 ][ 203 ],
   alphaCSR[ 115 ][ 204 ],
   alphaCSR[ 115 ][ 205 ],
   alphaCSR[ 115 ][ 206 ],
   alphaCSR[ 115 ][ 207 ],
   alphaCSR[ 115 ][ 208 ],
   alphaCSR[ 115 ][ 209 ],
   alphaCSR[ 115 ][ 210 ],
   alphaCSR[ 115 ][ 211 ],
   alphaCSR[ 115 ][ 212 ],
   alphaCSR[ 115 ][ 213 ],
   alphaCSR[ 115 ][ 214 ],
   alphaCSR[ 115 ][ 215 ],
   alphaCSR[ 115 ][ 216 ],
   alphaCSR[ 115 ][ 217 ],
   alphaCSR[ 115 ][ 218 ],
   alphaCSR[ 115 ][ 219 ],
   alphaCSR[ 115 ][ 220 ],
   alphaCSR[ 115 ][ 221 ],
   alphaCSR[ 115 ][ 222 ],
   alphaCSR[ 115 ][ 223 ],
   alphaCSR[ 115 ][ 224 ],
   alphaCSR[ 115 ][ 225 ],
   alphaCSR[ 115 ][ 226 ],
   alphaCSR[ 115 ][ 227 ],
   alphaCSR[ 115 ][ 228 ],
   alphaCSR[ 115 ][ 229 ],
   alphaCSR[ 115 ][ 230 ],
   alphaCSR[ 115 ][ 231 ],
   alphaCSR[ 115 ][ 232 ],
   alphaCSR[ 115 ][ 233 ],
   alphaCSR[ 115 ][ 234 ],
   alphaCSR[ 115 ][ 235 ],
   alphaCSR[ 115 ][ 236 ],
   alphaCSR[ 115 ][ 237 ],
   alphaCSR[ 115 ][ 238 ],
   alphaCSR[ 115 ][ 239 ],
   alphaCSR[ 115 ][ 240 ],
   alphaCSR[ 115 ][ 241 ],
   alphaCSR[ 115 ][ 242 ],
   alphaCSR[ 115 ][ 243 ],
   alphaCSR[ 115 ][ 244 ],
   alphaCSR[ 115 ][ 245 ],
   alphaCSR[ 115 ][ 246 ],
   alphaCSR[ 115 ][ 247 ],
   alphaCSR[ 115 ][ 248 ],
   alphaCSR[ 115 ][ 249 ],
   alphaCSR[ 115 ][ 250 ],
   alphaCSR[ 115 ][ 251 ],
   alphaCSR[ 115 ][ 252 ],
   alphaCSR[ 115 ][ 253 ],
   alphaCSR[ 115 ][ 254 ],
   alphaCSR[ 115 ][ 255 ],
   alphaCSR[ 115 ][ 256 ],
   alphaCSR[ 115 ][ 257 ],
   alphaCSR[ 115 ][ 258 ],
   alphaCSR[ 115 ][ 259 ],
   alphaCSR[ 115 ][ 260 ],
   alphaCSR[ 115 ][ 261 ],
   alphaCSR[ 115 ][ 262 ],
   alphaCSR[ 115 ][ 263 ],
   alphaCSR[ 115 ][ 264 ],
   alphaCSR[ 115 ][ 265 ],
   alphaCSR[ 115 ][ 266 ],
   alphaCSR[ 115 ][ 267 ],
   alphaCSR[ 115 ][ 268 ],
   alphaCSR[ 115 ][ 269 ],
   alphaCSR[ 115 ][ 270 ],
   alphaCSR[ 115 ][ 271 ],
   alphaCSR[ 115 ][ 272 ],
   alphaCSR[ 115 ][ 273 ],
   alphaCSR[ 115 ][ 274 ],
   alphaCSR[ 115 ][ 275 ],
   alphaCSR[ 115 ][ 276 ],
   alphaCSR[ 115 ][ 277 ],
   alphaCSR[ 115 ][ 278 ],
   alphaCSR[ 115 ][ 279 ],
   alphaCSR[ 115 ][ 280 ],
   alphaCSR[ 115 ][ 281 ],
   alphaCSR[ 115 ][ 282 ],
   alphaCSR[ 115 ][ 283 ],
   alphaCSR[ 115 ][ 284 ],
   alphaCSR[ 115 ][ 285 ],
   alphaCSR[ 115 ][ 286 ],
   alphaCSR[ 115 ][ 287 ],
   alphaCSR[ 115 ][ 288 ],
   alphaCSR[ 115 ][ 289 ],
   alphaCSR[ 115 ][ 290 ],
   alphaCSR[ 115 ][ 291 ],
   alphaCSR[ 115 ][ 292 ],
   alphaCSR[ 115 ][ 293 ],
   alphaCSR[ 115 ][ 294 ],
   alphaCSR[ 115 ][ 295 ],
   alphaCSR[ 115 ][ 296 ],
   alphaCSR[ 115 ][ 297 ],
   alphaCSR[ 115 ][ 298 ],
   alphaCSR[ 115 ][ 299 ],
   alphaCSR[ 115 ][ 300 ],
   alphaCSR[ 115 ][ 301 ],
   alphaCSR[ 115 ][ 302 ],
   alphaCSR[ 115 ][ 303 ],
   alphaCSR[ 115 ][ 304 ],
   alphaCSR[ 115 ][ 305 ],
   alphaCSR[ 115 ][ 306 ],
   alphaCSR[ 115 ][ 307 ],
   alphaCSR[ 115 ][ 308 ],
   alphaCSR[ 115 ][ 309 ],
   alphaCSR[ 115 ][ 310 ],
   alphaCSR[ 115 ][ 311 ],
   alphaCSR[ 115 ][ 312 ],
   alphaCSR[ 115 ][ 313 ],
   alphaCSR[ 115 ][ 314 ],
   alphaCSR[ 115 ][ 315 ],
   alphaCSR[ 115 ][ 316 ],
   alphaCSR[ 115 ][ 317 ],
   alphaCSR[ 115 ][ 318 ],
   alphaCSR[ 115 ][ 319 ],
   alphaCSR[ 115 ][ 320 ],
   alphaCSR[ 115 ][ 321 ],
   alphaCSR[ 115 ][ 322 ],
   alphaCSR[ 115 ][ 323 ],
   alphaCSR[ 115 ][ 324 ],
   alphaCSR[ 115 ][ 325 ],
   alphaCSR[ 115 ][ 326 ],
   alphaCSR[ 115 ][ 327 ],
   alphaCSR[ 115 ][ 328 ],
   alphaCSR[ 115 ][ 329 ],
   alphaCSR[ 115 ][ 330 ],
   alphaCSR[ 115 ][ 331 ],
   alphaCSR[ 115 ][ 332 ],
   alphaCSR[ 115 ][ 333 ],
   alphaCSR[ 115 ][ 334 ],
   alphaCSR[ 115 ][ 335 ],
   alphaCSR[ 115 ][ 336 ],
   alphaCSR[ 115 ][ 337 ],
   alphaCSR[ 115 ][ 338 ],
   alphaCSR[ 115 ][ 339 ],
   alphaCSR[ 115 ][ 340 ],
   alphaCSR[ 115 ][ 341 ],
   alphaCSR[ 115 ][ 342 ],
   alphaCSR[ 115 ][ 343 ],
   alphaCSR[ 115 ][ 344 ],
   alphaCSR[ 115 ][ 345 ],
   alphaCSR[ 115 ][ 346 ],
   alphaCSR[ 115 ][ 347 ],
   alphaCSR[ 115 ][ 348 ],
   alphaCSR[ 115 ][ 349 ],
   alphaCSR[ 115 ][ 350 ],
   alphaCSR[ 115 ][ 351 ],
   alphaCSR[ 115 ][ 352 ],
   alphaCSR[ 115 ][ 353 ],
   alphaCSR[ 115 ][ 354 ],
   alphaCSR[ 115 ][ 355 ],
   alphaCSR[ 115 ][ 356 ],
   alphaCSR[ 115 ][ 357 ],
   alphaCSR[ 115 ][ 358 ],
   alphaCSR[ 115 ][ 359 ],
   alphaCSR[ 115 ][ 360 ],
   alphaCSR[ 115 ][ 361 ],
   alphaCSR[ 115 ][ 362 ],
   alphaCSR[ 115 ][ 363 ],
   alphaCSR[ 115 ][ 364 ],
   alphaCSR[ 115 ][ 365 ],
   alphaCSR[ 115 ][ 366 ],
   alphaCSR[ 115 ][ 367 ],
   alphaCSR[ 115 ][ 368 ],
   alphaCSR[ 115 ][ 369 ],
   alphaCSR[ 115 ][ 370 ],
   alphaCSR[ 115 ][ 371 ],
   alphaCSR[ 115 ][ 372 ],
   alphaCSR[ 115 ][ 373 ],
   alphaCSR[ 115 ][ 374 ],
   alphaCSR[ 115 ][ 375 ],
   alphaCSR[ 115 ][ 376 ],
   alphaCSR[ 115 ][ 377 ],
   alphaCSR[ 115 ][ 378 ],
   alphaCSR[ 115 ][ 379 ],
   alphaCSR[ 115 ][ 380 ],
   alphaCSR[ 115 ][ 381 ],
   alphaCSR[ 115 ][ 382 ],
   alphaCSR[ 115 ][ 383 ],
   alphaCSR[ 116 ][ 0 ],
   alphaCSR[ 116 ][ 1 ],
   alphaCSR[ 116 ][ 2 ],
   alphaCSR[ 116 ][ 3 ],
   alphaCSR[ 116 ][ 4 ],
   alphaCSR[ 116 ][ 5 ],
   alphaCSR[ 116 ][ 6 ],
   alphaCSR[ 116 ][ 7 ],
   alphaCSR[ 116 ][ 8 ],
   alphaCSR[ 116 ][ 9 ],
   alphaCSR[ 116 ][ 10 ],
   alphaCSR[ 116 ][ 11 ],
   alphaCSR[ 116 ][ 12 ],
   alphaCSR[ 116 ][ 13 ],
   alphaCSR[ 116 ][ 14 ],
   alphaCSR[ 116 ][ 15 ],
   alphaCSR[ 116 ][ 16 ],
   alphaCSR[ 116 ][ 17 ],
   alphaCSR[ 116 ][ 18 ],
   alphaCSR[ 116 ][ 19 ],
   alphaCSR[ 116 ][ 20 ],
   alphaCSR[ 116 ][ 21 ],
   alphaCSR[ 116 ][ 22 ],
   alphaCSR[ 116 ][ 23 ],
   alphaCSR[ 116 ][ 24 ],
   alphaCSR[ 116 ][ 25 ],
   alphaCSR[ 116 ][ 26 ],
   alphaCSR[ 116 ][ 27 ],
   alphaCSR[ 116 ][ 28 ],
   alphaCSR[ 116 ][ 29 ],
   alphaCSR[ 116 ][ 30 ],
   alphaCSR[ 116 ][ 31 ],
   alphaCSR[ 116 ][ 32 ],
   alphaCSR[ 116 ][ 33 ],
   alphaCSR[ 116 ][ 34 ],
   alphaCSR[ 116 ][ 35 ],
   alphaCSR[ 116 ][ 36 ],
   alphaCSR[ 116 ][ 37 ],
   alphaCSR[ 116 ][ 38 ],
   alphaCSR[ 116 ][ 39 ],
   alphaCSR[ 116 ][ 40 ],
   alphaCSR[ 116 ][ 41 ],
   alphaCSR[ 116 ][ 42 ],
   alphaCSR[ 116 ][ 43 ],
   alphaCSR[ 116 ][ 44 ],
   alphaCSR[ 116 ][ 45 ],
   alphaCSR[ 116 ][ 46 ],
   alphaCSR[ 116 ][ 47 ],
   alphaCSR[ 116 ][ 48 ],
   alphaCSR[ 116 ][ 49 ],
   alphaCSR[ 116 ][ 50 ],
   alphaCSR[ 116 ][ 51 ],
   alphaCSR[ 116 ][ 52 ],
   alphaCSR[ 116 ][ 53 ],
   alphaCSR[ 116 ][ 54 ],
   alphaCSR[ 116 ][ 55 ],
   alphaCSR[ 116 ][ 56 ],
   alphaCSR[ 116 ][ 57 ],
   alphaCSR[ 116 ][ 58 ],
   alphaCSR[ 116 ][ 59 ],
   alphaCSR[ 116 ][ 60 ],
   alphaCSR[ 116 ][ 61 ],
   alphaCSR[ 116 ][ 62 ],
   alphaCSR[ 116 ][ 63 ],
   alphaCSR[ 116 ][ 64 ],
   alphaCSR[ 116 ][ 65 ],
   alphaCSR[ 116 ][ 66 ],
   alphaCSR[ 116 ][ 67 ],
   alphaCSR[ 116 ][ 68 ],
   alphaCSR[ 116 ][ 69 ],
   alphaCSR[ 116 ][ 70 ],
   alphaCSR[ 116 ][ 71 ],
   alphaCSR[ 116 ][ 72 ],
   alphaCSR[ 116 ][ 73 ],
   alphaCSR[ 116 ][ 74 ],
   alphaCSR[ 116 ][ 75 ],
   alphaCSR[ 116 ][ 76 ],
   alphaCSR[ 116 ][ 77 ],
   alphaCSR[ 116 ][ 78 ],
   alphaCSR[ 116 ][ 79 ],
   alphaCSR[ 116 ][ 80 ],
   alphaCSR[ 116 ][ 81 ],
   alphaCSR[ 116 ][ 82 ],
   alphaCSR[ 116 ][ 83 ],
   alphaCSR[ 116 ][ 84 ],
   alphaCSR[ 116 ][ 85 ],
   alphaCSR[ 116 ][ 86 ],
   alphaCSR[ 116 ][ 87 ],
   alphaCSR[ 116 ][ 88 ],
   alphaCSR[ 116 ][ 89 ],
   alphaCSR[ 116 ][ 90 ],
   alphaCSR[ 116 ][ 91 ],
   alphaCSR[ 116 ][ 92 ],
   alphaCSR[ 116 ][ 93 ],
   alphaCSR[ 116 ][ 94 ],
   alphaCSR[ 116 ][ 95 ],
   alphaCSR[ 116 ][ 96 ],
   alphaCSR[ 116 ][ 97 ],
   alphaCSR[ 116 ][ 98 ],
   alphaCSR[ 116 ][ 99 ],
   alphaCSR[ 116 ][ 100 ],
   alphaCSR[ 116 ][ 101 ],
   alphaCSR[ 116 ][ 102 ],
   alphaCSR[ 116 ][ 103 ],
   alphaCSR[ 116 ][ 104 ],
   alphaCSR[ 116 ][ 105 ],
   alphaCSR[ 116 ][ 106 ],
   alphaCSR[ 116 ][ 107 ],
   alphaCSR[ 116 ][ 108 ],
   alphaCSR[ 116 ][ 109 ],
   alphaCSR[ 116 ][ 110 ],
   alphaCSR[ 116 ][ 111 ],
   alphaCSR[ 116 ][ 112 ],
   alphaCSR[ 116 ][ 113 ],
   alphaCSR[ 116 ][ 114 ],
   alphaCSR[ 116 ][ 115 ],
   alphaCSR[ 116 ][ 116 ],
   alphaCSR[ 116 ][ 117 ],
   alphaCSR[ 116 ][ 118 ],
   alphaCSR[ 116 ][ 119 ],
   alphaCSR[ 116 ][ 120 ],
   alphaCSR[ 116 ][ 121 ],
   alphaCSR[ 116 ][ 122 ],
   alphaCSR[ 116 ][ 123 ],
   alphaCSR[ 116 ][ 124 ],
   alphaCSR[ 116 ][ 125 ],
   alphaCSR[ 116 ][ 126 ],
   alphaCSR[ 116 ][ 127 ],
   alphaCSR[ 116 ][ 128 ],
   alphaCSR[ 116 ][ 129 ],
   alphaCSR[ 116 ][ 130 ],
   alphaCSR[ 116 ][ 131 ],
   alphaCSR[ 116 ][ 132 ],
   alphaCSR[ 116 ][ 133 ],
   alphaCSR[ 116 ][ 134 ],
   alphaCSR[ 116 ][ 135 ],
   alphaCSR[ 116 ][ 136 ],
   alphaCSR[ 116 ][ 137 ],
   alphaCSR[ 116 ][ 138 ],
   alphaCSR[ 116 ][ 139 ],
   alphaCSR[ 116 ][ 140 ],
   alphaCSR[ 116 ][ 141 ],
   alphaCSR[ 116 ][ 142 ],
   alphaCSR[ 116 ][ 143 ],
   alphaCSR[ 116 ][ 144 ],
   alphaCSR[ 116 ][ 145 ],
   alphaCSR[ 116 ][ 146 ],
   alphaCSR[ 116 ][ 147 ],
   alphaCSR[ 116 ][ 148 ],
   alphaCSR[ 116 ][ 149 ],
   alphaCSR[ 116 ][ 150 ],
   alphaCSR[ 116 ][ 151 ],
   alphaCSR[ 116 ][ 152 ],
   alphaCSR[ 116 ][ 153 ],
   alphaCSR[ 116 ][ 154 ],
   alphaCSR[ 116 ][ 155 ],
   alphaCSR[ 116 ][ 156 ],
   alphaCSR[ 116 ][ 157 ],
   alphaCSR[ 116 ][ 158 ],
   alphaCSR[ 116 ][ 159 ],
   alphaCSR[ 116 ][ 160 ],
   alphaCSR[ 116 ][ 161 ],
   alphaCSR[ 116 ][ 162 ],
   alphaCSR[ 116 ][ 163 ],
   alphaCSR[ 116 ][ 164 ],
   alphaCSR[ 116 ][ 165 ],
   alphaCSR[ 116 ][ 166 ],
   alphaCSR[ 116 ][ 167 ],
   alphaCSR[ 116 ][ 168 ],
   alphaCSR[ 116 ][ 169 ],
   alphaCSR[ 116 ][ 170 ],
   alphaCSR[ 116 ][ 171 ],
   alphaCSR[ 116 ][ 172 ],
   alphaCSR[ 116 ][ 173 ],
   alphaCSR[ 116 ][ 174 ],
   alphaCSR[ 116 ][ 175 ],
   alphaCSR[ 116 ][ 176 ],
   alphaCSR[ 116 ][ 177 ],
   alphaCSR[ 116 ][ 178 ],
   alphaCSR[ 116 ][ 179 ],
   alphaCSR[ 116 ][ 180 ],
   alphaCSR[ 116 ][ 181 ],
   alphaCSR[ 116 ][ 182 ],
   alphaCSR[ 116 ][ 183 ],
   alphaCSR[ 116 ][ 184 ],
   alphaCSR[ 116 ][ 185 ],
   alphaCSR[ 116 ][ 186 ],
   alphaCSR[ 116 ][ 187 ],
   alphaCSR[ 116 ][ 188 ],
   alphaCSR[ 116 ][ 189 ],
   alphaCSR[ 116 ][ 190 ],
   alphaCSR[ 116 ][ 191 ],
   alphaCSR[ 116 ][ 192 ],
   alphaCSR[ 116 ][ 193 ],
   alphaCSR[ 116 ][ 194 ],
   alphaCSR[ 116 ][ 195 ],
   alphaCSR[ 116 ][ 196 ],
   alphaCSR[ 116 ][ 197 ],
   alphaCSR[ 116 ][ 198 ],
   alphaCSR[ 116 ][ 199 ],
   alphaCSR[ 116 ][ 200 ],
   alphaCSR[ 116 ][ 201 ],
   alphaCSR[ 116 ][ 202 ],
   alphaCSR[ 116 ][ 203 ],
   alphaCSR[ 116 ][ 204 ],
   alphaCSR[ 116 ][ 205 ],
   alphaCSR[ 116 ][ 206 ],
   alphaCSR[ 116 ][ 207 ],
   alphaCSR[ 116 ][ 208 ],
   alphaCSR[ 116 ][ 209 ],
   alphaCSR[ 116 ][ 210 ],
   alphaCSR[ 116 ][ 211 ],
   alphaCSR[ 116 ][ 212 ],
   alphaCSR[ 116 ][ 213 ],
   alphaCSR[ 116 ][ 214 ],
   alphaCSR[ 116 ][ 215 ],
   alphaCSR[ 116 ][ 216 ],
   alphaCSR[ 116 ][ 217 ],
   alphaCSR[ 116 ][ 218 ],
   alphaCSR[ 116 ][ 219 ],
   alphaCSR[ 116 ][ 220 ],
   alphaCSR[ 116 ][ 221 ],
   alphaCSR[ 116 ][ 222 ],
   alphaCSR[ 116 ][ 223 ],
   alphaCSR[ 116 ][ 224 ],
   alphaCSR[ 116 ][ 225 ],
   alphaCSR[ 116 ][ 226 ],
   alphaCSR[ 116 ][ 227 ],
   alphaCSR[ 116 ][ 228 ],
   alphaCSR[ 116 ][ 229 ],
   alphaCSR[ 116 ][ 230 ],
   alphaCSR[ 116 ][ 231 ],
   alphaCSR[ 116 ][ 232 ],
   alphaCSR[ 116 ][ 233 ],
   alphaCSR[ 116 ][ 234 ],
   alphaCSR[ 116 ][ 235 ],
   alphaCSR[ 116 ][ 236 ],
   alphaCSR[ 116 ][ 237 ],
   alphaCSR[ 116 ][ 238 ],
   alphaCSR[ 116 ][ 239 ],
   alphaCSR[ 116 ][ 240 ],
   alphaCSR[ 116 ][ 241 ],
   alphaCSR[ 116 ][ 242 ],
   alphaCSR[ 116 ][ 243 ],
   alphaCSR[ 116 ][ 244 ],
   alphaCSR[ 116 ][ 245 ],
   alphaCSR[ 116 ][ 246 ],
   alphaCSR[ 116 ][ 247 ],
   alphaCSR[ 116 ][ 248 ],
   alphaCSR[ 116 ][ 249 ],
   alphaCSR[ 116 ][ 250 ],
   alphaCSR[ 116 ][ 251 ],
   alphaCSR[ 116 ][ 252 ],
   alphaCSR[ 116 ][ 253 ],
   alphaCSR[ 116 ][ 254 ],
   alphaCSR[ 116 ][ 255 ],
   alphaCSR[ 116 ][ 256 ],
   alphaCSR[ 116 ][ 257 ],
   alphaCSR[ 116 ][ 258 ],
   alphaCSR[ 116 ][ 259 ],
   alphaCSR[ 116 ][ 260 ],
   alphaCSR[ 116 ][ 261 ],
   alphaCSR[ 116 ][ 262 ],
   alphaCSR[ 116 ][ 263 ],
   alphaCSR[ 116 ][ 264 ],
   alphaCSR[ 116 ][ 265 ],
   alphaCSR[ 116 ][ 266 ],
   alphaCSR[ 116 ][ 267 ],
   alphaCSR[ 116 ][ 268 ],
   alphaCSR[ 116 ][ 269 ],
   alphaCSR[ 116 ][ 270 ],
   alphaCSR[ 116 ][ 271 ],
   alphaCSR[ 116 ][ 272 ],
   alphaCSR[ 116 ][ 273 ],
   alphaCSR[ 116 ][ 274 ],
   alphaCSR[ 116 ][ 275 ],
   alphaCSR[ 116 ][ 276 ],
   alphaCSR[ 116 ][ 277 ],
   alphaCSR[ 116 ][ 278 ],
   alphaCSR[ 116 ][ 279 ],
   alphaCSR[ 116 ][ 280 ],
   alphaCSR[ 116 ][ 281 ],
   alphaCSR[ 116 ][ 282 ],
   alphaCSR[ 116 ][ 283 ],
   alphaCSR[ 116 ][ 284 ],
   alphaCSR[ 116 ][ 285 ],
   alphaCSR[ 116 ][ 286 ],
   alphaCSR[ 116 ][ 287 ],
   alphaCSR[ 116 ][ 288 ],
   alphaCSR[ 116 ][ 289 ],
   alphaCSR[ 116 ][ 290 ],
   alphaCSR[ 116 ][ 291 ],
   alphaCSR[ 116 ][ 292 ],
   alphaCSR[ 116 ][ 293 ],
   alphaCSR[ 116 ][ 294 ],
   alphaCSR[ 116 ][ 295 ],
   alphaCSR[ 116 ][ 296 ],
   alphaCSR[ 116 ][ 297 ],
   alphaCSR[ 116 ][ 298 ],
   alphaCSR[ 116 ][ 299 ],
   alphaCSR[ 116 ][ 300 ],
   alphaCSR[ 116 ][ 301 ],
   alphaCSR[ 116 ][ 302 ],
   alphaCSR[ 116 ][ 303 ],
   alphaCSR[ 116 ][ 304 ],
   alphaCSR[ 116 ][ 305 ],
   alphaCSR[ 116 ][ 306 ],
   alphaCSR[ 116 ][ 307 ],
   alphaCSR[ 116 ][ 308 ],
   alphaCSR[ 116 ][ 309 ],
   alphaCSR[ 116 ][ 310 ],
   alphaCSR[ 116 ][ 311 ],
   alphaCSR[ 116 ][ 312 ],
   alphaCSR[ 116 ][ 313 ],
   alphaCSR[ 116 ][ 314 ],
   alphaCSR[ 116 ][ 315 ],
   alphaCSR[ 116 ][ 316 ],
   alphaCSR[ 116 ][ 317 ],
   alphaCSR[ 116 ][ 318 ],
   alphaCSR[ 116 ][ 319 ],
   alphaCSR[ 116 ][ 320 ],
   alphaCSR[ 116 ][ 321 ],
   alphaCSR[ 116 ][ 322 ],
   alphaCSR[ 116 ][ 323 ],
   alphaCSR[ 116 ][ 324 ],
   alphaCSR[ 116 ][ 325 ],
   alphaCSR[ 116 ][ 326 ],
   alphaCSR[ 116 ][ 327 ],
   alphaCSR[ 116 ][ 328 ],
   alphaCSR[ 116 ][ 329 ],
   alphaCSR[ 116 ][ 330 ],
   alphaCSR[ 116 ][ 331 ],
   alphaCSR[ 116 ][ 332 ],
   alphaCSR[ 116 ][ 333 ],
   alphaCSR[ 116 ][ 334 ],
   alphaCSR[ 116 ][ 335 ],
   alphaCSR[ 116 ][ 336 ],
   alphaCSR[ 116 ][ 337 ],
   alphaCSR[ 116 ][ 338 ],
   alphaCSR[ 116 ][ 339 ],
   alphaCSR[ 116 ][ 340 ],
   alphaCSR[ 116 ][ 341 ],
   alphaCSR[ 116 ][ 342 ],
   alphaCSR[ 116 ][ 343 ],
   alphaCSR[ 116 ][ 344 ],
   alphaCSR[ 116 ][ 345 ],
   alphaCSR[ 116 ][ 346 ],
   alphaCSR[ 116 ][ 347 ],
   alphaCSR[ 116 ][ 348 ],
   alphaCSR[ 116 ][ 349 ],
   alphaCSR[ 116 ][ 350 ],
   alphaCSR[ 116 ][ 351 ],
   alphaCSR[ 116 ][ 352 ],
   alphaCSR[ 116 ][ 353 ],
   alphaCSR[ 116 ][ 354 ],
   alphaCSR[ 116 ][ 355 ],
   alphaCSR[ 116 ][ 356 ],
   alphaCSR[ 116 ][ 357 ],
   alphaCSR[ 116 ][ 358 ],
   alphaCSR[ 116 ][ 359 ],
   alphaCSR[ 116 ][ 360 ],
   alphaCSR[ 116 ][ 361 ],
   alphaCSR[ 116 ][ 362 ],
   alphaCSR[ 116 ][ 363 ],
   alphaCSR[ 116 ][ 364 ],
   alphaCSR[ 116 ][ 365 ],
   alphaCSR[ 116 ][ 366 ],
   alphaCSR[ 116 ][ 367 ],
   alphaCSR[ 116 ][ 368 ],
   alphaCSR[ 116 ][ 369 ],
   alphaCSR[ 116 ][ 370 ],
   alphaCSR[ 116 ][ 371 ],
   alphaCSR[ 116 ][ 372 ],
   alphaCSR[ 116 ][ 373 ],
   alphaCSR[ 116 ][ 374 ],
   alphaCSR[ 116 ][ 375 ],
   alphaCSR[ 116 ][ 376 ],
   alphaCSR[ 116 ][ 377 ],
   alphaCSR[ 116 ][ 378 ],
   alphaCSR[ 116 ][ 379 ],
   alphaCSR[ 116 ][ 380 ],
   alphaCSR[ 116 ][ 381 ],
   alphaCSR[ 116 ][ 382 ],
   alphaCSR[ 116 ][ 383 ],
   alphaCSR[ 117 ][ 0 ],
   alphaCSR[ 117 ][ 1 ],
   alphaCSR[ 117 ][ 2 ],
   alphaCSR[ 117 ][ 3 ],
   alphaCSR[ 117 ][ 4 ],
   alphaCSR[ 117 ][ 5 ],
   alphaCSR[ 117 ][ 6 ],
   alphaCSR[ 117 ][ 7 ],
   alphaCSR[ 117 ][ 8 ],
   alphaCSR[ 117 ][ 9 ],
   alphaCSR[ 117 ][ 10 ],
   alphaCSR[ 117 ][ 11 ],
   alphaCSR[ 117 ][ 12 ],
   alphaCSR[ 117 ][ 13 ],
   alphaCSR[ 117 ][ 14 ],
   alphaCSR[ 117 ][ 15 ],
   alphaCSR[ 117 ][ 16 ],
   alphaCSR[ 117 ][ 17 ],
   alphaCSR[ 117 ][ 18 ],
   alphaCSR[ 117 ][ 19 ],
   alphaCSR[ 117 ][ 20 ],
   alphaCSR[ 117 ][ 21 ],
   alphaCSR[ 117 ][ 22 ],
   alphaCSR[ 117 ][ 23 ],
   alphaCSR[ 117 ][ 24 ],
   alphaCSR[ 117 ][ 25 ],
   alphaCSR[ 117 ][ 26 ],
   alphaCSR[ 117 ][ 27 ],
   alphaCSR[ 117 ][ 28 ],
   alphaCSR[ 117 ][ 29 ],
   alphaCSR[ 117 ][ 30 ],
   alphaCSR[ 117 ][ 31 ],
   alphaCSR[ 117 ][ 32 ],
   alphaCSR[ 117 ][ 33 ],
   alphaCSR[ 117 ][ 34 ],
   alphaCSR[ 117 ][ 35 ],
   alphaCSR[ 117 ][ 36 ],
   alphaCSR[ 117 ][ 37 ],
   alphaCSR[ 117 ][ 38 ],
   alphaCSR[ 117 ][ 39 ],
   alphaCSR[ 117 ][ 40 ],
   alphaCSR[ 117 ][ 41 ],
   alphaCSR[ 117 ][ 42 ],
   alphaCSR[ 117 ][ 43 ],
   alphaCSR[ 117 ][ 44 ],
   alphaCSR[ 117 ][ 45 ],
   alphaCSR[ 117 ][ 46 ],
   alphaCSR[ 117 ][ 47 ],
   alphaCSR[ 117 ][ 48 ],
   alphaCSR[ 117 ][ 49 ],
   alphaCSR[ 117 ][ 50 ],
   alphaCSR[ 117 ][ 51 ],
   alphaCSR[ 117 ][ 52 ],
   alphaCSR[ 117 ][ 53 ],
   alphaCSR[ 117 ][ 54 ],
   alphaCSR[ 117 ][ 55 ],
   alphaCSR[ 117 ][ 56 ],
   alphaCSR[ 117 ][ 57 ],
   alphaCSR[ 117 ][ 58 ],
   alphaCSR[ 117 ][ 59 ],
   alphaCSR[ 117 ][ 60 ],
   alphaCSR[ 117 ][ 61 ],
   alphaCSR[ 117 ][ 62 ],
   alphaCSR[ 117 ][ 63 ],
   alphaCSR[ 117 ][ 64 ],
   alphaCSR[ 117 ][ 65 ],
   alphaCSR[ 117 ][ 66 ],
   alphaCSR[ 117 ][ 67 ],
   alphaCSR[ 117 ][ 68 ],
   alphaCSR[ 117 ][ 69 ],
   alphaCSR[ 117 ][ 70 ],
   alphaCSR[ 117 ][ 71 ],
   alphaCSR[ 117 ][ 72 ],
   alphaCSR[ 117 ][ 73 ],
   alphaCSR[ 117 ][ 74 ],
   alphaCSR[ 117 ][ 75 ],
   alphaCSR[ 117 ][ 76 ],
   alphaCSR[ 117 ][ 77 ],
   alphaCSR[ 117 ][ 78 ],
   alphaCSR[ 117 ][ 79 ],
   alphaCSR[ 117 ][ 80 ],
   alphaCSR[ 117 ][ 81 ],
   alphaCSR[ 117 ][ 82 ],
   alphaCSR[ 117 ][ 83 ],
   alphaCSR[ 117 ][ 84 ],
   alphaCSR[ 117 ][ 85 ],
   alphaCSR[ 117 ][ 86 ],
   alphaCSR[ 117 ][ 87 ],
   alphaCSR[ 117 ][ 88 ],
   alphaCSR[ 117 ][ 89 ],
   alphaCSR[ 117 ][ 90 ],
   alphaCSR[ 117 ][ 91 ],
   alphaCSR[ 117 ][ 92 ],
   alphaCSR[ 117 ][ 93 ],
   alphaCSR[ 117 ][ 94 ],
   alphaCSR[ 117 ][ 95 ],
   alphaCSR[ 117 ][ 96 ],
   alphaCSR[ 117 ][ 97 ],
   alphaCSR[ 117 ][ 98 ],
   alphaCSR[ 117 ][ 99 ],
   alphaCSR[ 117 ][ 100 ],
   alphaCSR[ 117 ][ 101 ],
   alphaCSR[ 117 ][ 102 ],
   alphaCSR[ 117 ][ 103 ],
   alphaCSR[ 117 ][ 104 ],
   alphaCSR[ 117 ][ 105 ],
   alphaCSR[ 117 ][ 106 ],
   alphaCSR[ 117 ][ 107 ],
   alphaCSR[ 117 ][ 108 ],
   alphaCSR[ 117 ][ 109 ],
   alphaCSR[ 117 ][ 110 ],
   alphaCSR[ 117 ][ 111 ],
   alphaCSR[ 117 ][ 112 ],
   alphaCSR[ 117 ][ 113 ],
   alphaCSR[ 117 ][ 114 ],
   alphaCSR[ 117 ][ 115 ],
   alphaCSR[ 117 ][ 116 ],
   alphaCSR[ 117 ][ 117 ],
   alphaCSR[ 117 ][ 118 ],
   alphaCSR[ 117 ][ 119 ],
   alphaCSR[ 117 ][ 120 ],
   alphaCSR[ 117 ][ 121 ],
   alphaCSR[ 117 ][ 122 ],
   alphaCSR[ 117 ][ 123 ],
   alphaCSR[ 117 ][ 124 ],
   alphaCSR[ 117 ][ 125 ],
   alphaCSR[ 117 ][ 126 ],
   alphaCSR[ 117 ][ 127 ],
   alphaCSR[ 117 ][ 128 ],
   alphaCSR[ 117 ][ 129 ],
   alphaCSR[ 117 ][ 130 ],
   alphaCSR[ 117 ][ 131 ],
   alphaCSR[ 117 ][ 132 ],
   alphaCSR[ 117 ][ 133 ],
   alphaCSR[ 117 ][ 134 ],
   alphaCSR[ 117 ][ 135 ],
   alphaCSR[ 117 ][ 136 ],
   alphaCSR[ 117 ][ 137 ],
   alphaCSR[ 117 ][ 138 ],
   alphaCSR[ 117 ][ 139 ],
   alphaCSR[ 117 ][ 140 ],
   alphaCSR[ 117 ][ 141 ],
   alphaCSR[ 117 ][ 142 ],
   alphaCSR[ 117 ][ 143 ],
   alphaCSR[ 117 ][ 144 ],
   alphaCSR[ 117 ][ 145 ],
   alphaCSR[ 117 ][ 146 ],
   alphaCSR[ 117 ][ 147 ],
   alphaCSR[ 117 ][ 148 ],
   alphaCSR[ 117 ][ 149 ],
   alphaCSR[ 117 ][ 150 ],
   alphaCSR[ 117 ][ 151 ],
   alphaCSR[ 117 ][ 152 ],
   alphaCSR[ 117 ][ 153 ],
   alphaCSR[ 117 ][ 154 ],
   alphaCSR[ 117 ][ 155 ],
   alphaCSR[ 117 ][ 156 ],
   alphaCSR[ 117 ][ 157 ],
   alphaCSR[ 117 ][ 158 ],
   alphaCSR[ 117 ][ 159 ],
   alphaCSR[ 117 ][ 160 ],
   alphaCSR[ 117 ][ 161 ],
   alphaCSR[ 117 ][ 162 ],
   alphaCSR[ 117 ][ 163 ],
   alphaCSR[ 117 ][ 164 ],
   alphaCSR[ 117 ][ 165 ],
   alphaCSR[ 117 ][ 166 ],
   alphaCSR[ 117 ][ 167 ],
   alphaCSR[ 117 ][ 168 ],
   alphaCSR[ 117 ][ 169 ],
   alphaCSR[ 117 ][ 170 ],
   alphaCSR[ 117 ][ 171 ],
   alphaCSR[ 117 ][ 172 ],
   alphaCSR[ 117 ][ 173 ],
   alphaCSR[ 117 ][ 174 ],
   alphaCSR[ 117 ][ 175 ],
   alphaCSR[ 117 ][ 176 ],
   alphaCSR[ 117 ][ 177 ],
   alphaCSR[ 117 ][ 178 ],
   alphaCSR[ 117 ][ 179 ],
   alphaCSR[ 117 ][ 180 ],
   alphaCSR[ 117 ][ 181 ],
   alphaCSR[ 117 ][ 182 ],
   alphaCSR[ 117 ][ 183 ],
   alphaCSR[ 117 ][ 184 ],
   alphaCSR[ 117 ][ 185 ],
   alphaCSR[ 117 ][ 186 ],
   alphaCSR[ 117 ][ 187 ],
   alphaCSR[ 117 ][ 188 ],
   alphaCSR[ 117 ][ 189 ],
   alphaCSR[ 117 ][ 190 ],
   alphaCSR[ 117 ][ 191 ],
   alphaCSR[ 117 ][ 192 ],
   alphaCSR[ 117 ][ 193 ],
   alphaCSR[ 117 ][ 194 ],
   alphaCSR[ 117 ][ 195 ],
   alphaCSR[ 117 ][ 196 ],
   alphaCSR[ 117 ][ 197 ],
   alphaCSR[ 117 ][ 198 ],
   alphaCSR[ 117 ][ 199 ],
   alphaCSR[ 117 ][ 200 ],
   alphaCSR[ 117 ][ 201 ],
   alphaCSR[ 117 ][ 202 ],
   alphaCSR[ 117 ][ 203 ],
   alphaCSR[ 117 ][ 204 ],
   alphaCSR[ 117 ][ 205 ],
   alphaCSR[ 117 ][ 206 ],
   alphaCSR[ 117 ][ 207 ],
   alphaCSR[ 117 ][ 208 ],
   alphaCSR[ 117 ][ 209 ],
   alphaCSR[ 117 ][ 210 ],
   alphaCSR[ 117 ][ 211 ],
   alphaCSR[ 117 ][ 212 ],
   alphaCSR[ 117 ][ 213 ],
   alphaCSR[ 117 ][ 214 ],
   alphaCSR[ 117 ][ 215 ],
   alphaCSR[ 117 ][ 216 ],
   alphaCSR[ 117 ][ 217 ],
   alphaCSR[ 117 ][ 218 ],
   alphaCSR[ 117 ][ 219 ],
   alphaCSR[ 117 ][ 220 ],
   alphaCSR[ 117 ][ 221 ],
   alphaCSR[ 117 ][ 222 ],
   alphaCSR[ 117 ][ 223 ],
   alphaCSR[ 117 ][ 224 ],
   alphaCSR[ 117 ][ 225 ],
   alphaCSR[ 117 ][ 226 ],
   alphaCSR[ 117 ][ 227 ],
   alphaCSR[ 117 ][ 228 ],
   alphaCSR[ 117 ][ 229 ],
   alphaCSR[ 117 ][ 230 ],
   alphaCSR[ 117 ][ 231 ],
   alphaCSR[ 117 ][ 232 ],
   alphaCSR[ 117 ][ 233 ],
   alphaCSR[ 117 ][ 234 ],
   alphaCSR[ 117 ][ 235 ],
   alphaCSR[ 117 ][ 236 ],
   alphaCSR[ 117 ][ 237 ],
   alphaCSR[ 117 ][ 238 ],
   alphaCSR[ 117 ][ 239 ],
   alphaCSR[ 117 ][ 240 ],
   alphaCSR[ 117 ][ 241 ],
   alphaCSR[ 117 ][ 242 ],
   alphaCSR[ 117 ][ 243 ],
   alphaCSR[ 117 ][ 244 ],
   alphaCSR[ 117 ][ 245 ],
   alphaCSR[ 117 ][ 246 ],
   alphaCSR[ 117 ][ 247 ],
   alphaCSR[ 117 ][ 248 ],
   alphaCSR[ 117 ][ 249 ],
   alphaCSR[ 117 ][ 250 ],
   alphaCSR[ 117 ][ 251 ],
   alphaCSR[ 117 ][ 252 ],
   alphaCSR[ 117 ][ 253 ],
   alphaCSR[ 117 ][ 254 ],
   alphaCSR[ 117 ][ 255 ],
   alphaCSR[ 117 ][ 256 ],
   alphaCSR[ 117 ][ 257 ],
   alphaCSR[ 117 ][ 258 ],
   alphaCSR[ 117 ][ 259 ],
   alphaCSR[ 117 ][ 260 ],
   alphaCSR[ 117 ][ 261 ],
   alphaCSR[ 117 ][ 262 ],
   alphaCSR[ 117 ][ 263 ],
   alphaCSR[ 117 ][ 264 ],
   alphaCSR[ 117 ][ 265 ],
   alphaCSR[ 117 ][ 266 ],
   alphaCSR[ 117 ][ 267 ],
   alphaCSR[ 117 ][ 268 ],
   alphaCSR[ 117 ][ 269 ],
   alphaCSR[ 117 ][ 270 ],
   alphaCSR[ 117 ][ 271 ],
   alphaCSR[ 117 ][ 272 ],
   alphaCSR[ 117 ][ 273 ],
   alphaCSR[ 117 ][ 274 ],
   alphaCSR[ 117 ][ 275 ],
   alphaCSR[ 117 ][ 276 ],
   alphaCSR[ 117 ][ 277 ],
   alphaCSR[ 117 ][ 278 ],
   alphaCSR[ 117 ][ 279 ],
   alphaCSR[ 117 ][ 280 ],
   alphaCSR[ 117 ][ 281 ],
   alphaCSR[ 117 ][ 282 ],
   alphaCSR[ 117 ][ 283 ],
   alphaCSR[ 117 ][ 284 ],
   alphaCSR[ 117 ][ 285 ],
   alphaCSR[ 117 ][ 286 ],
   alphaCSR[ 117 ][ 287 ],
   alphaCSR[ 117 ][ 288 ],
   alphaCSR[ 117 ][ 289 ],
   alphaCSR[ 117 ][ 290 ],
   alphaCSR[ 117 ][ 291 ],
   alphaCSR[ 117 ][ 292 ],
   alphaCSR[ 117 ][ 293 ],
   alphaCSR[ 117 ][ 294 ],
   alphaCSR[ 117 ][ 295 ],
   alphaCSR[ 117 ][ 296 ],
   alphaCSR[ 117 ][ 297 ],
   alphaCSR[ 117 ][ 298 ],
   alphaCSR[ 117 ][ 299 ],
   alphaCSR[ 117 ][ 300 ],
   alphaCSR[ 117 ][ 301 ],
   alphaCSR[ 117 ][ 302 ],
   alphaCSR[ 117 ][ 303 ],
   alphaCSR[ 117 ][ 304 ],
   alphaCSR[ 117 ][ 305 ],
   alphaCSR[ 117 ][ 306 ],
   alphaCSR[ 117 ][ 307 ],
   alphaCSR[ 117 ][ 308 ],
   alphaCSR[ 117 ][ 309 ],
   alphaCSR[ 117 ][ 310 ],
   alphaCSR[ 117 ][ 311 ],
   alphaCSR[ 117 ][ 312 ],
   alphaCSR[ 117 ][ 313 ],
   alphaCSR[ 117 ][ 314 ],
   alphaCSR[ 117 ][ 315 ],
   alphaCSR[ 117 ][ 316 ],
   alphaCSR[ 117 ][ 317 ],
   alphaCSR[ 117 ][ 318 ],
   alphaCSR[ 117 ][ 319 ],
   alphaCSR[ 117 ][ 320 ],
   alphaCSR[ 117 ][ 321 ],
   alphaCSR[ 117 ][ 322 ],
   alphaCSR[ 117 ][ 323 ],
   alphaCSR[ 117 ][ 324 ],
   alphaCSR[ 117 ][ 325 ],
   alphaCSR[ 117 ][ 326 ],
   alphaCSR[ 117 ][ 327 ],
   alphaCSR[ 117 ][ 328 ],
   alphaCSR[ 117 ][ 329 ],
   alphaCSR[ 117 ][ 330 ],
   alphaCSR[ 117 ][ 331 ],
   alphaCSR[ 117 ][ 332 ],
   alphaCSR[ 117 ][ 333 ],
   alphaCSR[ 117 ][ 334 ],
   alphaCSR[ 117 ][ 335 ],
   alphaCSR[ 117 ][ 336 ],
   alphaCSR[ 117 ][ 337 ],
   alphaCSR[ 117 ][ 338 ],
   alphaCSR[ 117 ][ 339 ],
   alphaCSR[ 117 ][ 340 ],
   alphaCSR[ 117 ][ 341 ],
   alphaCSR[ 117 ][ 342 ],
   alphaCSR[ 117 ][ 343 ],
   alphaCSR[ 117 ][ 344 ],
   alphaCSR[ 117 ][ 345 ],
   alphaCSR[ 117 ][ 346 ],
   alphaCSR[ 117 ][ 347 ],
   alphaCSR[ 117 ][ 348 ],
   alphaCSR[ 117 ][ 349 ],
   alphaCSR[ 117 ][ 350 ],
   alphaCSR[ 117 ][ 351 ],
   alphaCSR[ 117 ][ 352 ],
   alphaCSR[ 117 ][ 353 ],
   alphaCSR[ 117 ][ 354 ],
   alphaCSR[ 117 ][ 355 ],
   alphaCSR[ 117 ][ 356 ],
   alphaCSR[ 117 ][ 357 ],
   alphaCSR[ 117 ][ 358 ],
   alphaCSR[ 117 ][ 359 ],
   alphaCSR[ 117 ][ 360 ],
   alphaCSR[ 117 ][ 361 ],
   alphaCSR[ 117 ][ 362 ],
   alphaCSR[ 117 ][ 363 ],
   alphaCSR[ 117 ][ 364 ],
   alphaCSR[ 117 ][ 365 ],
   alphaCSR[ 117 ][ 366 ],
   alphaCSR[ 117 ][ 367 ],
   alphaCSR[ 117 ][ 368 ],
   alphaCSR[ 117 ][ 369 ],
   alphaCSR[ 117 ][ 370 ],
   alphaCSR[ 117 ][ 371 ],
   alphaCSR[ 117 ][ 372 ],
   alphaCSR[ 117 ][ 373 ],
   alphaCSR[ 117 ][ 374 ],
   alphaCSR[ 117 ][ 375 ],
   alphaCSR[ 117 ][ 376 ],
   alphaCSR[ 117 ][ 377 ],
   alphaCSR[ 117 ][ 378 ],
   alphaCSR[ 117 ][ 379 ],
   alphaCSR[ 117 ][ 380 ],
   alphaCSR[ 117 ][ 381 ],
   alphaCSR[ 117 ][ 382 ],
   alphaCSR[ 117 ][ 383 ],
   alphaCSR[ 118 ][ 0 ],
   alphaCSR[ 118 ][ 1 ],
   alphaCSR[ 118 ][ 2 ],
   alphaCSR[ 118 ][ 3 ],
   alphaCSR[ 118 ][ 4 ],
   alphaCSR[ 118 ][ 5 ],
   alphaCSR[ 118 ][ 6 ],
   alphaCSR[ 118 ][ 7 ],
   alphaCSR[ 118 ][ 8 ],
   alphaCSR[ 118 ][ 9 ],
   alphaCSR[ 118 ][ 10 ],
   alphaCSR[ 118 ][ 11 ],
   alphaCSR[ 118 ][ 12 ],
   alphaCSR[ 118 ][ 13 ],
   alphaCSR[ 118 ][ 14 ],
   alphaCSR[ 118 ][ 15 ],
   alphaCSR[ 118 ][ 16 ],
   alphaCSR[ 118 ][ 17 ],
   alphaCSR[ 118 ][ 18 ],
   alphaCSR[ 118 ][ 19 ],
   alphaCSR[ 118 ][ 20 ],
   alphaCSR[ 118 ][ 21 ],
   alphaCSR[ 118 ][ 22 ],
   alphaCSR[ 118 ][ 23 ],
   alphaCSR[ 118 ][ 24 ],
   alphaCSR[ 118 ][ 25 ],
   alphaCSR[ 118 ][ 26 ],
   alphaCSR[ 118 ][ 27 ],
   alphaCSR[ 118 ][ 28 ],
   alphaCSR[ 118 ][ 29 ],
   alphaCSR[ 118 ][ 30 ],
   alphaCSR[ 118 ][ 31 ],
   alphaCSR[ 118 ][ 32 ],
   alphaCSR[ 118 ][ 33 ],
   alphaCSR[ 118 ][ 34 ],
   alphaCSR[ 118 ][ 35 ],
   alphaCSR[ 118 ][ 36 ],
   alphaCSR[ 118 ][ 37 ],
   alphaCSR[ 118 ][ 38 ],
   alphaCSR[ 118 ][ 39 ],
   alphaCSR[ 118 ][ 40 ],
   alphaCSR[ 118 ][ 41 ],
   alphaCSR[ 118 ][ 42 ],
   alphaCSR[ 118 ][ 43 ],
   alphaCSR[ 118 ][ 44 ],
   alphaCSR[ 118 ][ 45 ],
   alphaCSR[ 118 ][ 46 ],
   alphaCSR[ 118 ][ 47 ],
   alphaCSR[ 118 ][ 48 ],
   alphaCSR[ 118 ][ 49 ],
   alphaCSR[ 118 ][ 50 ],
   alphaCSR[ 118 ][ 51 ],
   alphaCSR[ 118 ][ 52 ],
   alphaCSR[ 118 ][ 53 ],
   alphaCSR[ 118 ][ 54 ],
   alphaCSR[ 118 ][ 55 ],
   alphaCSR[ 118 ][ 56 ],
   alphaCSR[ 118 ][ 57 ],
   alphaCSR[ 118 ][ 58 ],
   alphaCSR[ 118 ][ 59 ],
   alphaCSR[ 118 ][ 60 ],
   alphaCSR[ 118 ][ 61 ],
   alphaCSR[ 118 ][ 62 ],
   alphaCSR[ 118 ][ 63 ],
   alphaCSR[ 118 ][ 64 ],
   alphaCSR[ 118 ][ 65 ],
   alphaCSR[ 118 ][ 66 ],
   alphaCSR[ 118 ][ 67 ],
   alphaCSR[ 118 ][ 68 ],
   alphaCSR[ 118 ][ 69 ],
   alphaCSR[ 118 ][ 70 ],
   alphaCSR[ 118 ][ 71 ],
   alphaCSR[ 118 ][ 72 ],
   alphaCSR[ 118 ][ 73 ],
   alphaCSR[ 118 ][ 74 ],
   alphaCSR[ 118 ][ 75 ],
   alphaCSR[ 118 ][ 76 ],
   alphaCSR[ 118 ][ 77 ],
   alphaCSR[ 118 ][ 78 ],
   alphaCSR[ 118 ][ 79 ],
   alphaCSR[ 118 ][ 80 ],
   alphaCSR[ 118 ][ 81 ],
   alphaCSR[ 118 ][ 82 ],
   alphaCSR[ 118 ][ 83 ],
   alphaCSR[ 118 ][ 84 ],
   alphaCSR[ 118 ][ 85 ],
   alphaCSR[ 118 ][ 86 ],
   alphaCSR[ 118 ][ 87 ],
   alphaCSR[ 118 ][ 88 ],
   alphaCSR[ 118 ][ 89 ],
   alphaCSR[ 118 ][ 90 ],
   alphaCSR[ 118 ][ 91 ],
   alphaCSR[ 118 ][ 92 ],
   alphaCSR[ 118 ][ 93 ],
   alphaCSR[ 118 ][ 94 ],
   alphaCSR[ 118 ][ 95 ],
   alphaCSR[ 118 ][ 96 ],
   alphaCSR[ 118 ][ 97 ],
   alphaCSR[ 118 ][ 98 ],
   alphaCSR[ 118 ][ 99 ],
   alphaCSR[ 118 ][ 100 ],
   alphaCSR[ 118 ][ 101 ],
   alphaCSR[ 118 ][ 102 ],
   alphaCSR[ 118 ][ 103 ],
   alphaCSR[ 118 ][ 104 ],
   alphaCSR[ 118 ][ 105 ],
   alphaCSR[ 118 ][ 106 ],
   alphaCSR[ 118 ][ 107 ],
   alphaCSR[ 118 ][ 108 ],
   alphaCSR[ 118 ][ 109 ],
   alphaCSR[ 118 ][ 110 ],
   alphaCSR[ 118 ][ 111 ],
   alphaCSR[ 118 ][ 112 ],
   alphaCSR[ 118 ][ 113 ],
   alphaCSR[ 118 ][ 114 ],
   alphaCSR[ 118 ][ 115 ],
   alphaCSR[ 118 ][ 116 ],
   alphaCSR[ 118 ][ 117 ],
   alphaCSR[ 118 ][ 118 ],
   alphaCSR[ 118 ][ 119 ],
   alphaCSR[ 118 ][ 120 ],
   alphaCSR[ 118 ][ 121 ],
   alphaCSR[ 118 ][ 122 ],
   alphaCSR[ 118 ][ 123 ],
   alphaCSR[ 118 ][ 124 ],
   alphaCSR[ 118 ][ 125 ],
   alphaCSR[ 118 ][ 126 ],
   alphaCSR[ 118 ][ 127 ],
   alphaCSR[ 118 ][ 128 ],
   alphaCSR[ 118 ][ 129 ],
   alphaCSR[ 118 ][ 130 ],
   alphaCSR[ 118 ][ 131 ],
   alphaCSR[ 118 ][ 132 ],
   alphaCSR[ 118 ][ 133 ],
   alphaCSR[ 118 ][ 134 ],
   alphaCSR[ 118 ][ 135 ],
   alphaCSR[ 118 ][ 136 ],
   alphaCSR[ 118 ][ 137 ],
   alphaCSR[ 118 ][ 138 ],
   alphaCSR[ 118 ][ 139 ],
   alphaCSR[ 118 ][ 140 ],
   alphaCSR[ 118 ][ 141 ],
   alphaCSR[ 118 ][ 142 ],
   alphaCSR[ 118 ][ 143 ],
   alphaCSR[ 118 ][ 144 ],
   alphaCSR[ 118 ][ 145 ],
   alphaCSR[ 118 ][ 146 ],
   alphaCSR[ 118 ][ 147 ],
   alphaCSR[ 118 ][ 148 ],
   alphaCSR[ 118 ][ 149 ],
   alphaCSR[ 118 ][ 150 ],
   alphaCSR[ 118 ][ 151 ],
   alphaCSR[ 118 ][ 152 ],
   alphaCSR[ 118 ][ 153 ],
   alphaCSR[ 118 ][ 154 ],
   alphaCSR[ 118 ][ 155 ],
   alphaCSR[ 118 ][ 156 ],
   alphaCSR[ 118 ][ 157 ],
   alphaCSR[ 118 ][ 158 ],
   alphaCSR[ 118 ][ 159 ],
   alphaCSR[ 118 ][ 160 ],
   alphaCSR[ 118 ][ 161 ],
   alphaCSR[ 118 ][ 162 ],
   alphaCSR[ 118 ][ 163 ],
   alphaCSR[ 118 ][ 164 ],
   alphaCSR[ 118 ][ 165 ],
   alphaCSR[ 118 ][ 166 ],
   alphaCSR[ 118 ][ 167 ],
   alphaCSR[ 118 ][ 168 ],
   alphaCSR[ 118 ][ 169 ],
   alphaCSR[ 118 ][ 170 ],
   alphaCSR[ 118 ][ 171 ],
   alphaCSR[ 118 ][ 172 ],
   alphaCSR[ 118 ][ 173 ],
   alphaCSR[ 118 ][ 174 ],
   alphaCSR[ 118 ][ 175 ],
   alphaCSR[ 118 ][ 176 ],
   alphaCSR[ 118 ][ 177 ],
   alphaCSR[ 118 ][ 178 ],
   alphaCSR[ 118 ][ 179 ],
   alphaCSR[ 118 ][ 180 ],
   alphaCSR[ 118 ][ 181 ],
   alphaCSR[ 118 ][ 182 ],
   alphaCSR[ 118 ][ 183 ],
   alphaCSR[ 118 ][ 184 ],
   alphaCSR[ 118 ][ 185 ],
   alphaCSR[ 118 ][ 186 ],
   alphaCSR[ 118 ][ 187 ],
   alphaCSR[ 118 ][ 188 ],
   alphaCSR[ 118 ][ 189 ],
   alphaCSR[ 118 ][ 190 ],
   alphaCSR[ 118 ][ 191 ],
   alphaCSR[ 118 ][ 192 ],
   alphaCSR[ 118 ][ 193 ],
   alphaCSR[ 118 ][ 194 ],
   alphaCSR[ 118 ][ 195 ],
   alphaCSR[ 118 ][ 196 ],
   alphaCSR[ 118 ][ 197 ],
   alphaCSR[ 118 ][ 198 ],
   alphaCSR[ 118 ][ 199 ],
   alphaCSR[ 118 ][ 200 ],
   alphaCSR[ 118 ][ 201 ],
   alphaCSR[ 118 ][ 202 ],
   alphaCSR[ 118 ][ 203 ],
   alphaCSR[ 118 ][ 204 ],
   alphaCSR[ 118 ][ 205 ],
   alphaCSR[ 118 ][ 206 ],
   alphaCSR[ 118 ][ 207 ],
   alphaCSR[ 118 ][ 208 ],
   alphaCSR[ 118 ][ 209 ],
   alphaCSR[ 118 ][ 210 ],
   alphaCSR[ 118 ][ 211 ],
   alphaCSR[ 118 ][ 212 ],
   alphaCSR[ 118 ][ 213 ],
   alphaCSR[ 118 ][ 214 ],
   alphaCSR[ 118 ][ 215 ],
   alphaCSR[ 118 ][ 216 ],
   alphaCSR[ 118 ][ 217 ],
   alphaCSR[ 118 ][ 218 ],
   alphaCSR[ 118 ][ 219 ],
   alphaCSR[ 118 ][ 220 ],
   alphaCSR[ 118 ][ 221 ],
   alphaCSR[ 118 ][ 222 ],
   alphaCSR[ 118 ][ 223 ],
   alphaCSR[ 118 ][ 224 ],
   alphaCSR[ 118 ][ 225 ],
   alphaCSR[ 118 ][ 226 ],
   alphaCSR[ 118 ][ 227 ],
   alphaCSR[ 118 ][ 228 ],
   alphaCSR[ 118 ][ 229 ],
   alphaCSR[ 118 ][ 230 ],
   alphaCSR[ 118 ][ 231 ],
   alphaCSR[ 118 ][ 232 ],
   alphaCSR[ 118 ][ 233 ],
   alphaCSR[ 118 ][ 234 ],
   alphaCSR[ 118 ][ 235 ],
   alphaCSR[ 118 ][ 236 ],
   alphaCSR[ 118 ][ 237 ],
   alphaCSR[ 118 ][ 238 ],
   alphaCSR[ 118 ][ 239 ],
   alphaCSR[ 118 ][ 240 ],
   alphaCSR[ 118 ][ 241 ],
   alphaCSR[ 118 ][ 242 ],
   alphaCSR[ 118 ][ 243 ],
   alphaCSR[ 118 ][ 244 ],
   alphaCSR[ 118 ][ 245 ],
   alphaCSR[ 118 ][ 246 ],
   alphaCSR[ 118 ][ 247 ],
   alphaCSR[ 118 ][ 248 ],
   alphaCSR[ 118 ][ 249 ],
   alphaCSR[ 118 ][ 250 ],
   alphaCSR[ 118 ][ 251 ],
   alphaCSR[ 118 ][ 252 ],
   alphaCSR[ 118 ][ 253 ],
   alphaCSR[ 118 ][ 254 ],
   alphaCSR[ 118 ][ 255 ],
   alphaCSR[ 118 ][ 256 ],
   alphaCSR[ 118 ][ 257 ],
   alphaCSR[ 118 ][ 258 ],
   alphaCSR[ 118 ][ 259 ],
   alphaCSR[ 118 ][ 260 ],
   alphaCSR[ 118 ][ 261 ],
   alphaCSR[ 118 ][ 262 ],
   alphaCSR[ 118 ][ 263 ],
   alphaCSR[ 118 ][ 264 ],
   alphaCSR[ 118 ][ 265 ],
   alphaCSR[ 118 ][ 266 ],
   alphaCSR[ 118 ][ 267 ],
   alphaCSR[ 118 ][ 268 ],
   alphaCSR[ 118 ][ 269 ],
   alphaCSR[ 118 ][ 270 ],
   alphaCSR[ 118 ][ 271 ],
   alphaCSR[ 118 ][ 272 ],
   alphaCSR[ 118 ][ 273 ],
   alphaCSR[ 118 ][ 274 ],
   alphaCSR[ 118 ][ 275 ],
   alphaCSR[ 118 ][ 276 ],
   alphaCSR[ 118 ][ 277 ],
   alphaCSR[ 118 ][ 278 ],
   alphaCSR[ 118 ][ 279 ],
   alphaCSR[ 118 ][ 280 ],
   alphaCSR[ 118 ][ 281 ],
   alphaCSR[ 118 ][ 282 ],
   alphaCSR[ 118 ][ 283 ],
   alphaCSR[ 118 ][ 284 ],
   alphaCSR[ 118 ][ 285 ],
   alphaCSR[ 118 ][ 286 ],
   alphaCSR[ 118 ][ 287 ],
   alphaCSR[ 118 ][ 288 ],
   alphaCSR[ 118 ][ 289 ],
   alphaCSR[ 118 ][ 290 ],
   alphaCSR[ 118 ][ 291 ],
   alphaCSR[ 118 ][ 292 ],
   alphaCSR[ 118 ][ 293 ],
   alphaCSR[ 118 ][ 294 ],
   alphaCSR[ 118 ][ 295 ],
   alphaCSR[ 118 ][ 296 ],
   alphaCSR[ 118 ][ 297 ],
   alphaCSR[ 118 ][ 298 ],
   alphaCSR[ 118 ][ 299 ],
   alphaCSR[ 118 ][ 300 ],
   alphaCSR[ 118 ][ 301 ],
   alphaCSR[ 118 ][ 302 ],
   alphaCSR[ 118 ][ 303 ],
   alphaCSR[ 118 ][ 304 ],
   alphaCSR[ 118 ][ 305 ],
   alphaCSR[ 118 ][ 306 ],
   alphaCSR[ 118 ][ 307 ],
   alphaCSR[ 118 ][ 308 ],
   alphaCSR[ 118 ][ 309 ],
   alphaCSR[ 118 ][ 310 ],
   alphaCSR[ 118 ][ 311 ],
   alphaCSR[ 118 ][ 312 ],
   alphaCSR[ 118 ][ 313 ],
   alphaCSR[ 118 ][ 314 ],
   alphaCSR[ 118 ][ 315 ],
   alphaCSR[ 118 ][ 316 ],
   alphaCSR[ 118 ][ 317 ],
   alphaCSR[ 118 ][ 318 ],
   alphaCSR[ 118 ][ 319 ],
   alphaCSR[ 118 ][ 320 ],
   alphaCSR[ 118 ][ 321 ],
   alphaCSR[ 118 ][ 322 ],
   alphaCSR[ 118 ][ 323 ],
   alphaCSR[ 118 ][ 324 ],
   alphaCSR[ 118 ][ 325 ],
   alphaCSR[ 118 ][ 326 ],
   alphaCSR[ 118 ][ 327 ],
   alphaCSR[ 118 ][ 328 ],
   alphaCSR[ 118 ][ 329 ],
   alphaCSR[ 118 ][ 330 ],
   alphaCSR[ 118 ][ 331 ],
   alphaCSR[ 118 ][ 332 ],
   alphaCSR[ 118 ][ 333 ],
   alphaCSR[ 118 ][ 334 ],
   alphaCSR[ 118 ][ 335 ],
   alphaCSR[ 118 ][ 336 ],
   alphaCSR[ 118 ][ 337 ],
   alphaCSR[ 118 ][ 338 ],
   alphaCSR[ 118 ][ 339 ],
   alphaCSR[ 118 ][ 340 ],
   alphaCSR[ 118 ][ 341 ],
   alphaCSR[ 118 ][ 342 ],
   alphaCSR[ 118 ][ 343 ],
   alphaCSR[ 118 ][ 344 ],
   alphaCSR[ 118 ][ 345 ],
   alphaCSR[ 118 ][ 346 ],
   alphaCSR[ 118 ][ 347 ],
   alphaCSR[ 118 ][ 348 ],
   alphaCSR[ 118 ][ 349 ],
   alphaCSR[ 118 ][ 350 ],
   alphaCSR[ 118 ][ 351 ],
   alphaCSR[ 118 ][ 352 ],
   alphaCSR[ 118 ][ 353 ],
   alphaCSR[ 118 ][ 354 ],
   alphaCSR[ 118 ][ 355 ],
   alphaCSR[ 118 ][ 356 ],
   alphaCSR[ 118 ][ 357 ],
   alphaCSR[ 118 ][ 358 ],
   alphaCSR[ 118 ][ 359 ],
   alphaCSR[ 118 ][ 360 ],
   alphaCSR[ 118 ][ 361 ],
   alphaCSR[ 118 ][ 362 ],
   alphaCSR[ 118 ][ 363 ],
   alphaCSR[ 118 ][ 364 ],
   alphaCSR[ 118 ][ 365 ],
   alphaCSR[ 118 ][ 366 ],
   alphaCSR[ 118 ][ 367 ],
   alphaCSR[ 118 ][ 368 ],
   alphaCSR[ 118 ][ 369 ],
   alphaCSR[ 118 ][ 370 ],
   alphaCSR[ 118 ][ 371 ],
   alphaCSR[ 118 ][ 372 ],
   alphaCSR[ 118 ][ 373 ],
   alphaCSR[ 118 ][ 374 ],
   alphaCSR[ 118 ][ 375 ],
   alphaCSR[ 118 ][ 376 ],
   alphaCSR[ 118 ][ 377 ],
   alphaCSR[ 118 ][ 378 ],
   alphaCSR[ 118 ][ 379 ],
   alphaCSR[ 118 ][ 380 ],
   alphaCSR[ 118 ][ 381 ],
   alphaCSR[ 118 ][ 382 ],
   alphaCSR[ 118 ][ 383 ],
   alphaCSR[ 119 ][ 0 ],
   alphaCSR[ 119 ][ 1 ],
   alphaCSR[ 119 ][ 2 ],
   alphaCSR[ 119 ][ 3 ],
   alphaCSR[ 119 ][ 4 ],
   alphaCSR[ 119 ][ 5 ],
   alphaCSR[ 119 ][ 6 ],
   alphaCSR[ 119 ][ 7 ],
   alphaCSR[ 119 ][ 8 ],
   alphaCSR[ 119 ][ 9 ],
   alphaCSR[ 119 ][ 10 ],
   alphaCSR[ 119 ][ 11 ],
   alphaCSR[ 119 ][ 12 ],
   alphaCSR[ 119 ][ 13 ],
   alphaCSR[ 119 ][ 14 ],
   alphaCSR[ 119 ][ 15 ],
   alphaCSR[ 119 ][ 16 ],
   alphaCSR[ 119 ][ 17 ],
   alphaCSR[ 119 ][ 18 ],
   alphaCSR[ 119 ][ 19 ],
   alphaCSR[ 119 ][ 20 ],
   alphaCSR[ 119 ][ 21 ],
   alphaCSR[ 119 ][ 22 ],
   alphaCSR[ 119 ][ 23 ],
   alphaCSR[ 119 ][ 24 ],
   alphaCSR[ 119 ][ 25 ],
   alphaCSR[ 119 ][ 26 ],
   alphaCSR[ 119 ][ 27 ],
   alphaCSR[ 119 ][ 28 ],
   alphaCSR[ 119 ][ 29 ],
   alphaCSR[ 119 ][ 30 ],
   alphaCSR[ 119 ][ 31 ],
   alphaCSR[ 119 ][ 32 ],
   alphaCSR[ 119 ][ 33 ],
   alphaCSR[ 119 ][ 34 ],
   alphaCSR[ 119 ][ 35 ],
   alphaCSR[ 119 ][ 36 ],
   alphaCSR[ 119 ][ 37 ],
   alphaCSR[ 119 ][ 38 ],
   alphaCSR[ 119 ][ 39 ],
   alphaCSR[ 119 ][ 40 ],
   alphaCSR[ 119 ][ 41 ],
   alphaCSR[ 119 ][ 42 ],
   alphaCSR[ 119 ][ 43 ],
   alphaCSR[ 119 ][ 44 ],
   alphaCSR[ 119 ][ 45 ],
   alphaCSR[ 119 ][ 46 ],
   alphaCSR[ 119 ][ 47 ],
   alphaCSR[ 119 ][ 48 ],
   alphaCSR[ 119 ][ 49 ],
   alphaCSR[ 119 ][ 50 ],
   alphaCSR[ 119 ][ 51 ],
   alphaCSR[ 119 ][ 52 ],
   alphaCSR[ 119 ][ 53 ],
   alphaCSR[ 119 ][ 54 ],
   alphaCSR[ 119 ][ 55 ],
   alphaCSR[ 119 ][ 56 ],
   alphaCSR[ 119 ][ 57 ],
   alphaCSR[ 119 ][ 58 ],
   alphaCSR[ 119 ][ 59 ],
   alphaCSR[ 119 ][ 60 ],
   alphaCSR[ 119 ][ 61 ],
   alphaCSR[ 119 ][ 62 ],
   alphaCSR[ 119 ][ 63 ],
   alphaCSR[ 119 ][ 64 ],
   alphaCSR[ 119 ][ 65 ],
   alphaCSR[ 119 ][ 66 ],
   alphaCSR[ 119 ][ 67 ],
   alphaCSR[ 119 ][ 68 ],
   alphaCSR[ 119 ][ 69 ],
   alphaCSR[ 119 ][ 70 ],
   alphaCSR[ 119 ][ 71 ],
   alphaCSR[ 119 ][ 72 ],
   alphaCSR[ 119 ][ 73 ],
   alphaCSR[ 119 ][ 74 ],
   alphaCSR[ 119 ][ 75 ],
   alphaCSR[ 119 ][ 76 ],
   alphaCSR[ 119 ][ 77 ],
   alphaCSR[ 119 ][ 78 ],
   alphaCSR[ 119 ][ 79 ],
   alphaCSR[ 119 ][ 80 ],
   alphaCSR[ 119 ][ 81 ],
   alphaCSR[ 119 ][ 82 ],
   alphaCSR[ 119 ][ 83 ],
   alphaCSR[ 119 ][ 84 ],
   alphaCSR[ 119 ][ 85 ],
   alphaCSR[ 119 ][ 86 ],
   alphaCSR[ 119 ][ 87 ],
   alphaCSR[ 119 ][ 88 ],
   alphaCSR[ 119 ][ 89 ],
   alphaCSR[ 119 ][ 90 ],
   alphaCSR[ 119 ][ 91 ],
   alphaCSR[ 119 ][ 92 ],
   alphaCSR[ 119 ][ 93 ],
   alphaCSR[ 119 ][ 94 ],
   alphaCSR[ 119 ][ 95 ],
   alphaCSR[ 119 ][ 96 ],
   alphaCSR[ 119 ][ 97 ],
   alphaCSR[ 119 ][ 98 ],
   alphaCSR[ 119 ][ 99 ],
   alphaCSR[ 119 ][ 100 ],
   alphaCSR[ 119 ][ 101 ],
   alphaCSR[ 119 ][ 102 ],
   alphaCSR[ 119 ][ 103 ],
   alphaCSR[ 119 ][ 104 ],
   alphaCSR[ 119 ][ 105 ],
   alphaCSR[ 119 ][ 106 ],
   alphaCSR[ 119 ][ 107 ],
   alphaCSR[ 119 ][ 108 ],
   alphaCSR[ 119 ][ 109 ],
   alphaCSR[ 119 ][ 110 ],
   alphaCSR[ 119 ][ 111 ],
   alphaCSR[ 119 ][ 112 ],
   alphaCSR[ 119 ][ 113 ],
   alphaCSR[ 119 ][ 114 ],
   alphaCSR[ 119 ][ 115 ],
   alphaCSR[ 119 ][ 116 ],
   alphaCSR[ 119 ][ 117 ],
   alphaCSR[ 119 ][ 118 ],
   alphaCSR[ 119 ][ 119 ],
   alphaCSR[ 119 ][ 120 ],
   alphaCSR[ 119 ][ 121 ],
   alphaCSR[ 119 ][ 122 ],
   alphaCSR[ 119 ][ 123 ],
   alphaCSR[ 119 ][ 124 ],
   alphaCSR[ 119 ][ 125 ],
   alphaCSR[ 119 ][ 126 ],
   alphaCSR[ 119 ][ 127 ],
   alphaCSR[ 119 ][ 128 ],
   alphaCSR[ 119 ][ 129 ],
   alphaCSR[ 119 ][ 130 ],
   alphaCSR[ 119 ][ 131 ],
   alphaCSR[ 119 ][ 132 ],
   alphaCSR[ 119 ][ 133 ],
   alphaCSR[ 119 ][ 134 ],
   alphaCSR[ 119 ][ 135 ],
   alphaCSR[ 119 ][ 136 ],
   alphaCSR[ 119 ][ 137 ],
   alphaCSR[ 119 ][ 138 ],
   alphaCSR[ 119 ][ 139 ],
   alphaCSR[ 119 ][ 140 ],
   alphaCSR[ 119 ][ 141 ],
   alphaCSR[ 119 ][ 142 ],
   alphaCSR[ 119 ][ 143 ],
   alphaCSR[ 119 ][ 144 ],
   alphaCSR[ 119 ][ 145 ],
   alphaCSR[ 119 ][ 146 ],
   alphaCSR[ 119 ][ 147 ],
   alphaCSR[ 119 ][ 148 ],
   alphaCSR[ 119 ][ 149 ],
   alphaCSR[ 119 ][ 150 ],
   alphaCSR[ 119 ][ 151 ],
   alphaCSR[ 119 ][ 152 ],
   alphaCSR[ 119 ][ 153 ],
   alphaCSR[ 119 ][ 154 ],
   alphaCSR[ 119 ][ 155 ],
   alphaCSR[ 119 ][ 156 ],
   alphaCSR[ 119 ][ 157 ],
   alphaCSR[ 119 ][ 158 ],
   alphaCSR[ 119 ][ 159 ],
   alphaCSR[ 119 ][ 160 ],
   alphaCSR[ 119 ][ 161 ],
   alphaCSR[ 119 ][ 162 ],
   alphaCSR[ 119 ][ 163 ],
   alphaCSR[ 119 ][ 164 ],
   alphaCSR[ 119 ][ 165 ],
   alphaCSR[ 119 ][ 166 ],
   alphaCSR[ 119 ][ 167 ],
   alphaCSR[ 119 ][ 168 ],
   alphaCSR[ 119 ][ 169 ],
   alphaCSR[ 119 ][ 170 ],
   alphaCSR[ 119 ][ 171 ],
   alphaCSR[ 119 ][ 172 ],
   alphaCSR[ 119 ][ 173 ],
   alphaCSR[ 119 ][ 174 ],
   alphaCSR[ 119 ][ 175 ],
   alphaCSR[ 119 ][ 176 ],
   alphaCSR[ 119 ][ 177 ],
   alphaCSR[ 119 ][ 178 ],
   alphaCSR[ 119 ][ 179 ],
   alphaCSR[ 119 ][ 180 ],
   alphaCSR[ 119 ][ 181 ],
   alphaCSR[ 119 ][ 182 ],
   alphaCSR[ 119 ][ 183 ],
   alphaCSR[ 119 ][ 184 ],
   alphaCSR[ 119 ][ 185 ],
   alphaCSR[ 119 ][ 186 ],
   alphaCSR[ 119 ][ 187 ],
   alphaCSR[ 119 ][ 188 ],
   alphaCSR[ 119 ][ 189 ],
   alphaCSR[ 119 ][ 190 ],
   alphaCSR[ 119 ][ 191 ],
   alphaCSR[ 119 ][ 192 ],
   alphaCSR[ 119 ][ 193 ],
   alphaCSR[ 119 ][ 194 ],
   alphaCSR[ 119 ][ 195 ],
   alphaCSR[ 119 ][ 196 ],
   alphaCSR[ 119 ][ 197 ],
   alphaCSR[ 119 ][ 198 ],
   alphaCSR[ 119 ][ 199 ],
   alphaCSR[ 119 ][ 200 ],
   alphaCSR[ 119 ][ 201 ],
   alphaCSR[ 119 ][ 202 ],
   alphaCSR[ 119 ][ 203 ],
   alphaCSR[ 119 ][ 204 ],
   alphaCSR[ 119 ][ 205 ],
   alphaCSR[ 119 ][ 206 ],
   alphaCSR[ 119 ][ 207 ],
   alphaCSR[ 119 ][ 208 ],
   alphaCSR[ 119 ][ 209 ],
   alphaCSR[ 119 ][ 210 ],
   alphaCSR[ 119 ][ 211 ],
   alphaCSR[ 119 ][ 212 ],
   alphaCSR[ 119 ][ 213 ],
   alphaCSR[ 119 ][ 214 ],
   alphaCSR[ 119 ][ 215 ],
   alphaCSR[ 119 ][ 216 ],
   alphaCSR[ 119 ][ 217 ],
   alphaCSR[ 119 ][ 218 ],
   alphaCSR[ 119 ][ 219 ],
   alphaCSR[ 119 ][ 220 ],
   alphaCSR[ 119 ][ 221 ],
   alphaCSR[ 119 ][ 222 ],
   alphaCSR[ 119 ][ 223 ],
   alphaCSR[ 119 ][ 224 ],
   alphaCSR[ 119 ][ 225 ],
   alphaCSR[ 119 ][ 226 ],
   alphaCSR[ 119 ][ 227 ],
   alphaCSR[ 119 ][ 228 ],
   alphaCSR[ 119 ][ 229 ],
   alphaCSR[ 119 ][ 230 ],
   alphaCSR[ 119 ][ 231 ],
   alphaCSR[ 119 ][ 232 ],
   alphaCSR[ 119 ][ 233 ],
   alphaCSR[ 119 ][ 234 ],
   alphaCSR[ 119 ][ 235 ],
   alphaCSR[ 119 ][ 236 ],
   alphaCSR[ 119 ][ 237 ],
   alphaCSR[ 119 ][ 238 ],
   alphaCSR[ 119 ][ 239 ],
   alphaCSR[ 119 ][ 240 ],
   alphaCSR[ 119 ][ 241 ],
   alphaCSR[ 119 ][ 242 ],
   alphaCSR[ 119 ][ 243 ],
   alphaCSR[ 119 ][ 244 ],
   alphaCSR[ 119 ][ 245 ],
   alphaCSR[ 119 ][ 246 ],
   alphaCSR[ 119 ][ 247 ],
   alphaCSR[ 119 ][ 248 ],
   alphaCSR[ 119 ][ 249 ],
   alphaCSR[ 119 ][ 250 ],
   alphaCSR[ 119 ][ 251 ],
   alphaCSR[ 119 ][ 252 ],
   alphaCSR[ 119 ][ 253 ],
   alphaCSR[ 119 ][ 254 ],
   alphaCSR[ 119 ][ 255 ],
   alphaCSR[ 119 ][ 256 ],
   alphaCSR[ 119 ][ 257 ],
   alphaCSR[ 119 ][ 258 ],
   alphaCSR[ 119 ][ 259 ],
   alphaCSR[ 119 ][ 260 ],
   alphaCSR[ 119 ][ 261 ],
   alphaCSR[ 119 ][ 262 ],
   alphaCSR[ 119 ][ 263 ],
   alphaCSR[ 119 ][ 264 ],
   alphaCSR[ 119 ][ 265 ],
   alphaCSR[ 119 ][ 266 ],
   alphaCSR[ 119 ][ 267 ],
   alphaCSR[ 119 ][ 268 ],
   alphaCSR[ 119 ][ 269 ],
   alphaCSR[ 119 ][ 270 ],
   alphaCSR[ 119 ][ 271 ],
   alphaCSR[ 119 ][ 272 ],
   alphaCSR[ 119 ][ 273 ],
   alphaCSR[ 119 ][ 274 ],
   alphaCSR[ 119 ][ 275 ],
   alphaCSR[ 119 ][ 276 ],
   alphaCSR[ 119 ][ 277 ],
   alphaCSR[ 119 ][ 278 ],
   alphaCSR[ 119 ][ 279 ],
   alphaCSR[ 119 ][ 280 ],
   alphaCSR[ 119 ][ 281 ],
   alphaCSR[ 119 ][ 282 ],
   alphaCSR[ 119 ][ 283 ],
   alphaCSR[ 119 ][ 284 ],
   alphaCSR[ 119 ][ 285 ],
   alphaCSR[ 119 ][ 286 ],
   alphaCSR[ 119 ][ 287 ],
   alphaCSR[ 119 ][ 288 ],
   alphaCSR[ 119 ][ 289 ],
   alphaCSR[ 119 ][ 290 ],
   alphaCSR[ 119 ][ 291 ],
   alphaCSR[ 119 ][ 292 ],
   alphaCSR[ 119 ][ 293 ],
   alphaCSR[ 119 ][ 294 ],
   alphaCSR[ 119 ][ 295 ],
   alphaCSR[ 119 ][ 296 ],
   alphaCSR[ 119 ][ 297 ],
   alphaCSR[ 119 ][ 298 ],
   alphaCSR[ 119 ][ 299 ],
   alphaCSR[ 119 ][ 300 ],
   alphaCSR[ 119 ][ 301 ],
   alphaCSR[ 119 ][ 302 ],
   alphaCSR[ 119 ][ 303 ],
   alphaCSR[ 119 ][ 304 ],
   alphaCSR[ 119 ][ 305 ],
   alphaCSR[ 119 ][ 306 ],
   alphaCSR[ 119 ][ 307 ],
   alphaCSR[ 119 ][ 308 ],
   alphaCSR[ 119 ][ 309 ],
   alphaCSR[ 119 ][ 310 ],
   alphaCSR[ 119 ][ 311 ],
   alphaCSR[ 119 ][ 312 ],
   alphaCSR[ 119 ][ 313 ],
   alphaCSR[ 119 ][ 314 ],
   alphaCSR[ 119 ][ 315 ],
   alphaCSR[ 119 ][ 316 ],
   alphaCSR[ 119 ][ 317 ],
   alphaCSR[ 119 ][ 318 ],
   alphaCSR[ 119 ][ 319 ],
   alphaCSR[ 119 ][ 320 ],
   alphaCSR[ 119 ][ 321 ],
   alphaCSR[ 119 ][ 322 ],
   alphaCSR[ 119 ][ 323 ],
   alphaCSR[ 119 ][ 324 ],
   alphaCSR[ 119 ][ 325 ],
   alphaCSR[ 119 ][ 326 ],
   alphaCSR[ 119 ][ 327 ],
   alphaCSR[ 119 ][ 328 ],
   alphaCSR[ 119 ][ 329 ],
   alphaCSR[ 119 ][ 330 ],
   alphaCSR[ 119 ][ 331 ],
   alphaCSR[ 119 ][ 332 ],
   alphaCSR[ 119 ][ 333 ],
   alphaCSR[ 119 ][ 334 ],
   alphaCSR[ 119 ][ 335 ],
   alphaCSR[ 119 ][ 336 ],
   alphaCSR[ 119 ][ 337 ],
   alphaCSR[ 119 ][ 338 ],
   alphaCSR[ 119 ][ 339 ],
   alphaCSR[ 119 ][ 340 ],
   alphaCSR[ 119 ][ 341 ],
   alphaCSR[ 119 ][ 342 ],
   alphaCSR[ 119 ][ 343 ],
   alphaCSR[ 119 ][ 344 ],
   alphaCSR[ 119 ][ 345 ],
   alphaCSR[ 119 ][ 346 ],
   alphaCSR[ 119 ][ 347 ],
   alphaCSR[ 119 ][ 348 ],
   alphaCSR[ 119 ][ 349 ],
   alphaCSR[ 119 ][ 350 ],
   alphaCSR[ 119 ][ 351 ],
   alphaCSR[ 119 ][ 352 ],
   alphaCSR[ 119 ][ 353 ],
   alphaCSR[ 119 ][ 354 ],
   alphaCSR[ 119 ][ 355 ],
   alphaCSR[ 119 ][ 356 ],
   alphaCSR[ 119 ][ 357 ],
   alphaCSR[ 119 ][ 358 ],
   alphaCSR[ 119 ][ 359 ],
   alphaCSR[ 119 ][ 360 ],
   alphaCSR[ 119 ][ 361 ],
   alphaCSR[ 119 ][ 362 ],
   alphaCSR[ 119 ][ 363 ],
   alphaCSR[ 119 ][ 364 ],
   alphaCSR[ 119 ][ 365 ],
   alphaCSR[ 119 ][ 366 ],
   alphaCSR[ 119 ][ 367 ],
   alphaCSR[ 119 ][ 368 ],
   alphaCSR[ 119 ][ 369 ],
   alphaCSR[ 119 ][ 370 ],
   alphaCSR[ 119 ][ 371 ],
   alphaCSR[ 119 ][ 372 ],
   alphaCSR[ 119 ][ 373 ],
   alphaCSR[ 119 ][ 374 ],
   alphaCSR[ 119 ][ 375 ],
   alphaCSR[ 119 ][ 376 ],
   alphaCSR[ 119 ][ 377 ],
   alphaCSR[ 119 ][ 378 ],
   alphaCSR[ 119 ][ 379 ],
   alphaCSR[ 119 ][ 380 ],
   alphaCSR[ 119 ][ 381 ],
   alphaCSR[ 119 ][ 382 ],
   alphaCSR[ 119 ][ 383 ],
   alphaCSR[ 120 ][ 0 ],
   alphaCSR[ 120 ][ 1 ],
   alphaCSR[ 120 ][ 2 ],
   alphaCSR[ 120 ][ 3 ],
   alphaCSR[ 120 ][ 4 ],
   alphaCSR[ 120 ][ 5 ],
   alphaCSR[ 120 ][ 6 ],
   alphaCSR[ 120 ][ 7 ],
   alphaCSR[ 120 ][ 8 ],
   alphaCSR[ 120 ][ 9 ],
   alphaCSR[ 120 ][ 10 ],
   alphaCSR[ 120 ][ 11 ],
   alphaCSR[ 120 ][ 12 ],
   alphaCSR[ 120 ][ 13 ],
   alphaCSR[ 120 ][ 14 ],
   alphaCSR[ 120 ][ 15 ],
   alphaCSR[ 120 ][ 16 ],
   alphaCSR[ 120 ][ 17 ],
   alphaCSR[ 120 ][ 18 ],
   alphaCSR[ 120 ][ 19 ],
   alphaCSR[ 120 ][ 20 ],
   alphaCSR[ 120 ][ 21 ],
   alphaCSR[ 120 ][ 22 ],
   alphaCSR[ 120 ][ 23 ],
   alphaCSR[ 120 ][ 24 ],
   alphaCSR[ 120 ][ 25 ],
   alphaCSR[ 120 ][ 26 ],
   alphaCSR[ 120 ][ 27 ],
   alphaCSR[ 120 ][ 28 ],
   alphaCSR[ 120 ][ 29 ],
   alphaCSR[ 120 ][ 30 ],
   alphaCSR[ 120 ][ 31 ],
   alphaCSR[ 120 ][ 32 ],
   alphaCSR[ 120 ][ 33 ],
   alphaCSR[ 120 ][ 34 ],
   alphaCSR[ 120 ][ 35 ],
   alphaCSR[ 120 ][ 36 ],
   alphaCSR[ 120 ][ 37 ],
   alphaCSR[ 120 ][ 38 ],
   alphaCSR[ 120 ][ 39 ],
   alphaCSR[ 120 ][ 40 ],
   alphaCSR[ 120 ][ 41 ],
   alphaCSR[ 120 ][ 42 ],
   alphaCSR[ 120 ][ 43 ],
   alphaCSR[ 120 ][ 44 ],
   alphaCSR[ 120 ][ 45 ],
   alphaCSR[ 120 ][ 46 ],
   alphaCSR[ 120 ][ 47 ],
   alphaCSR[ 120 ][ 48 ],
   alphaCSR[ 120 ][ 49 ],
   alphaCSR[ 120 ][ 50 ],
   alphaCSR[ 120 ][ 51 ],
   alphaCSR[ 120 ][ 52 ],
   alphaCSR[ 120 ][ 53 ],
   alphaCSR[ 120 ][ 54 ],
   alphaCSR[ 120 ][ 55 ],
   alphaCSR[ 120 ][ 56 ],
   alphaCSR[ 120 ][ 57 ],
   alphaCSR[ 120 ][ 58 ],
   alphaCSR[ 120 ][ 59 ],
   alphaCSR[ 120 ][ 60 ],
   alphaCSR[ 120 ][ 61 ],
   alphaCSR[ 120 ][ 62 ],
   alphaCSR[ 120 ][ 63 ],
   alphaCSR[ 120 ][ 64 ],
   alphaCSR[ 120 ][ 65 ],
   alphaCSR[ 120 ][ 66 ],
   alphaCSR[ 120 ][ 67 ],
   alphaCSR[ 120 ][ 68 ],
   alphaCSR[ 120 ][ 69 ],
   alphaCSR[ 120 ][ 70 ],
   alphaCSR[ 120 ][ 71 ],
   alphaCSR[ 120 ][ 72 ],
   alphaCSR[ 120 ][ 73 ],
   alphaCSR[ 120 ][ 74 ],
   alphaCSR[ 120 ][ 75 ],
   alphaCSR[ 120 ][ 76 ],
   alphaCSR[ 120 ][ 77 ],
   alphaCSR[ 120 ][ 78 ],
   alphaCSR[ 120 ][ 79 ],
   alphaCSR[ 120 ][ 80 ],
   alphaCSR[ 120 ][ 81 ],
   alphaCSR[ 120 ][ 82 ],
   alphaCSR[ 120 ][ 83 ],
   alphaCSR[ 120 ][ 84 ],
   alphaCSR[ 120 ][ 85 ],
   alphaCSR[ 120 ][ 86 ],
   alphaCSR[ 120 ][ 87 ],
   alphaCSR[ 120 ][ 88 ],
   alphaCSR[ 120 ][ 89 ],
   alphaCSR[ 120 ][ 90 ],
   alphaCSR[ 120 ][ 91 ],
   alphaCSR[ 120 ][ 92 ],
   alphaCSR[ 120 ][ 93 ],
   alphaCSR[ 120 ][ 94 ],
   alphaCSR[ 120 ][ 95 ],
   alphaCSR[ 120 ][ 96 ],
   alphaCSR[ 120 ][ 97 ],
   alphaCSR[ 120 ][ 98 ],
   alphaCSR[ 120 ][ 99 ],
   alphaCSR[ 120 ][ 100 ],
   alphaCSR[ 120 ][ 101 ],
   alphaCSR[ 120 ][ 102 ],
   alphaCSR[ 120 ][ 103 ],
   alphaCSR[ 120 ][ 104 ],
   alphaCSR[ 120 ][ 105 ],
   alphaCSR[ 120 ][ 106 ],
   alphaCSR[ 120 ][ 107 ],
   alphaCSR[ 120 ][ 108 ],
   alphaCSR[ 120 ][ 109 ],
   alphaCSR[ 120 ][ 110 ],
   alphaCSR[ 120 ][ 111 ],
   alphaCSR[ 120 ][ 112 ],
   alphaCSR[ 120 ][ 113 ],
   alphaCSR[ 120 ][ 114 ],
   alphaCSR[ 120 ][ 115 ],
   alphaCSR[ 120 ][ 116 ],
   alphaCSR[ 120 ][ 117 ],
   alphaCSR[ 120 ][ 118 ],
   alphaCSR[ 120 ][ 119 ],
   alphaCSR[ 120 ][ 120 ],
   alphaCSR[ 120 ][ 121 ],
   alphaCSR[ 120 ][ 122 ],
   alphaCSR[ 120 ][ 123 ],
   alphaCSR[ 120 ][ 124 ],
   alphaCSR[ 120 ][ 125 ],
   alphaCSR[ 120 ][ 126 ],
   alphaCSR[ 120 ][ 127 ],
   alphaCSR[ 120 ][ 128 ],
   alphaCSR[ 120 ][ 129 ],
   alphaCSR[ 120 ][ 130 ],
   alphaCSR[ 120 ][ 131 ],
   alphaCSR[ 120 ][ 132 ],
   alphaCSR[ 120 ][ 133 ],
   alphaCSR[ 120 ][ 134 ],
   alphaCSR[ 120 ][ 135 ],
   alphaCSR[ 120 ][ 136 ],
   alphaCSR[ 120 ][ 137 ],
   alphaCSR[ 120 ][ 138 ],
   alphaCSR[ 120 ][ 139 ],
   alphaCSR[ 120 ][ 140 ],
   alphaCSR[ 120 ][ 141 ],
   alphaCSR[ 120 ][ 142 ],
   alphaCSR[ 120 ][ 143 ],
   alphaCSR[ 120 ][ 144 ],
   alphaCSR[ 120 ][ 145 ],
   alphaCSR[ 120 ][ 146 ],
   alphaCSR[ 120 ][ 147 ],
   alphaCSR[ 120 ][ 148 ],
   alphaCSR[ 120 ][ 149 ],
   alphaCSR[ 120 ][ 150 ],
   alphaCSR[ 120 ][ 151 ],
   alphaCSR[ 120 ][ 152 ],
   alphaCSR[ 120 ][ 153 ],
   alphaCSR[ 120 ][ 154 ],
   alphaCSR[ 120 ][ 155 ],
   alphaCSR[ 120 ][ 156 ],
   alphaCSR[ 120 ][ 157 ],
   alphaCSR[ 120 ][ 158 ],
   alphaCSR[ 120 ][ 159 ],
   alphaCSR[ 120 ][ 160 ],
   alphaCSR[ 120 ][ 161 ],
   alphaCSR[ 120 ][ 162 ],
   alphaCSR[ 120 ][ 163 ],
   alphaCSR[ 120 ][ 164 ],
   alphaCSR[ 120 ][ 165 ],
   alphaCSR[ 120 ][ 166 ],
   alphaCSR[ 120 ][ 167 ],
   alphaCSR[ 120 ][ 168 ],
   alphaCSR[ 120 ][ 169 ],
   alphaCSR[ 120 ][ 170 ],
   alphaCSR[ 120 ][ 171 ],
   alphaCSR[ 120 ][ 172 ],
   alphaCSR[ 120 ][ 173 ],
   alphaCSR[ 120 ][ 174 ],
   alphaCSR[ 120 ][ 175 ],
   alphaCSR[ 120 ][ 176 ],
   alphaCSR[ 120 ][ 177 ],
   alphaCSR[ 120 ][ 178 ],
   alphaCSR[ 120 ][ 179 ],
   alphaCSR[ 120 ][ 180 ],
   alphaCSR[ 120 ][ 181 ],
   alphaCSR[ 120 ][ 182 ],
   alphaCSR[ 120 ][ 183 ],
   alphaCSR[ 120 ][ 184 ],
   alphaCSR[ 120 ][ 185 ],
   alphaCSR[ 120 ][ 186 ],
   alphaCSR[ 120 ][ 187 ],
   alphaCSR[ 120 ][ 188 ],
   alphaCSR[ 120 ][ 189 ],
   alphaCSR[ 120 ][ 190 ],
   alphaCSR[ 120 ][ 191 ],
   alphaCSR[ 120 ][ 192 ],
   alphaCSR[ 120 ][ 193 ],
   alphaCSR[ 120 ][ 194 ],
   alphaCSR[ 120 ][ 195 ],
   alphaCSR[ 120 ][ 196 ],
   alphaCSR[ 120 ][ 197 ],
   alphaCSR[ 120 ][ 198 ],
   alphaCSR[ 120 ][ 199 ],
   alphaCSR[ 120 ][ 200 ],
   alphaCSR[ 120 ][ 201 ],
   alphaCSR[ 120 ][ 202 ],
   alphaCSR[ 120 ][ 203 ],
   alphaCSR[ 120 ][ 204 ],
   alphaCSR[ 120 ][ 205 ],
   alphaCSR[ 120 ][ 206 ],
   alphaCSR[ 120 ][ 207 ],
   alphaCSR[ 120 ][ 208 ],
   alphaCSR[ 120 ][ 209 ],
   alphaCSR[ 120 ][ 210 ],
   alphaCSR[ 120 ][ 211 ],
   alphaCSR[ 120 ][ 212 ],
   alphaCSR[ 120 ][ 213 ],
   alphaCSR[ 120 ][ 214 ],
   alphaCSR[ 120 ][ 215 ],
   alphaCSR[ 120 ][ 216 ],
   alphaCSR[ 120 ][ 217 ],
   alphaCSR[ 120 ][ 218 ],
   alphaCSR[ 120 ][ 219 ],
   alphaCSR[ 120 ][ 220 ],
   alphaCSR[ 120 ][ 221 ],
   alphaCSR[ 120 ][ 222 ],
   alphaCSR[ 120 ][ 223 ],
   alphaCSR[ 120 ][ 224 ],
   alphaCSR[ 120 ][ 225 ],
   alphaCSR[ 120 ][ 226 ],
   alphaCSR[ 120 ][ 227 ],
   alphaCSR[ 120 ][ 228 ],
   alphaCSR[ 120 ][ 229 ],
   alphaCSR[ 120 ][ 230 ],
   alphaCSR[ 120 ][ 231 ],
   alphaCSR[ 120 ][ 232 ],
   alphaCSR[ 120 ][ 233 ],
   alphaCSR[ 120 ][ 234 ],
   alphaCSR[ 120 ][ 235 ],
   alphaCSR[ 120 ][ 236 ],
   alphaCSR[ 120 ][ 237 ],
   alphaCSR[ 120 ][ 238 ],
   alphaCSR[ 120 ][ 239 ],
   alphaCSR[ 120 ][ 240 ],
   alphaCSR[ 120 ][ 241 ],
   alphaCSR[ 120 ][ 242 ],
   alphaCSR[ 120 ][ 243 ],
   alphaCSR[ 120 ][ 244 ],
   alphaCSR[ 120 ][ 245 ],
   alphaCSR[ 120 ][ 246 ],
   alphaCSR[ 120 ][ 247 ],
   alphaCSR[ 120 ][ 248 ],
   alphaCSR[ 120 ][ 249 ],
   alphaCSR[ 120 ][ 250 ],
   alphaCSR[ 120 ][ 251 ],
   alphaCSR[ 120 ][ 252 ],
   alphaCSR[ 120 ][ 253 ],
   alphaCSR[ 120 ][ 254 ],
   alphaCSR[ 120 ][ 255 ],
   alphaCSR[ 120 ][ 256 ],
   alphaCSR[ 120 ][ 257 ],
   alphaCSR[ 120 ][ 258 ],
   alphaCSR[ 120 ][ 259 ],
   alphaCSR[ 120 ][ 260 ],
   alphaCSR[ 120 ][ 261 ],
   alphaCSR[ 120 ][ 262 ],
   alphaCSR[ 120 ][ 263 ],
   alphaCSR[ 120 ][ 264 ],
   alphaCSR[ 120 ][ 265 ],
   alphaCSR[ 120 ][ 266 ],
   alphaCSR[ 120 ][ 267 ],
   alphaCSR[ 120 ][ 268 ],
   alphaCSR[ 120 ][ 269 ],
   alphaCSR[ 120 ][ 270 ],
   alphaCSR[ 120 ][ 271 ],
   alphaCSR[ 120 ][ 272 ],
   alphaCSR[ 120 ][ 273 ],
   alphaCSR[ 120 ][ 274 ],
   alphaCSR[ 120 ][ 275 ],
   alphaCSR[ 120 ][ 276 ],
   alphaCSR[ 120 ][ 277 ],
   alphaCSR[ 120 ][ 278 ],
   alphaCSR[ 120 ][ 279 ],
   alphaCSR[ 120 ][ 280 ],
   alphaCSR[ 120 ][ 281 ],
   alphaCSR[ 120 ][ 282 ],
   alphaCSR[ 120 ][ 283 ],
   alphaCSR[ 120 ][ 284 ],
   alphaCSR[ 120 ][ 285 ],
   alphaCSR[ 120 ][ 286 ],
   alphaCSR[ 120 ][ 287 ],
   alphaCSR[ 120 ][ 288 ],
   alphaCSR[ 120 ][ 289 ],
   alphaCSR[ 120 ][ 290 ],
   alphaCSR[ 120 ][ 291 ],
   alphaCSR[ 120 ][ 292 ],
   alphaCSR[ 120 ][ 293 ],
   alphaCSR[ 120 ][ 294 ],
   alphaCSR[ 120 ][ 295 ],
   alphaCSR[ 120 ][ 296 ],
   alphaCSR[ 120 ][ 297 ],
   alphaCSR[ 120 ][ 298 ],
   alphaCSR[ 120 ][ 299 ],
   alphaCSR[ 120 ][ 300 ],
   alphaCSR[ 120 ][ 301 ],
   alphaCSR[ 120 ][ 302 ],
   alphaCSR[ 120 ][ 303 ],
   alphaCSR[ 120 ][ 304 ],
   alphaCSR[ 120 ][ 305 ],
   alphaCSR[ 120 ][ 306 ],
   alphaCSR[ 120 ][ 307 ],
   alphaCSR[ 120 ][ 308 ],
   alphaCSR[ 120 ][ 309 ],
   alphaCSR[ 120 ][ 310 ],
   alphaCSR[ 120 ][ 311 ],
   alphaCSR[ 120 ][ 312 ],
   alphaCSR[ 120 ][ 313 ],
   alphaCSR[ 120 ][ 314 ],
   alphaCSR[ 120 ][ 315 ],
   alphaCSR[ 120 ][ 316 ],
   alphaCSR[ 120 ][ 317 ],
   alphaCSR[ 120 ][ 318 ],
   alphaCSR[ 120 ][ 319 ],
   alphaCSR[ 120 ][ 320 ],
   alphaCSR[ 120 ][ 321 ],
   alphaCSR[ 120 ][ 322 ],
   alphaCSR[ 120 ][ 323 ],
   alphaCSR[ 120 ][ 324 ],
   alphaCSR[ 120 ][ 325 ],
   alphaCSR[ 120 ][ 326 ],
   alphaCSR[ 120 ][ 327 ],
   alphaCSR[ 120 ][ 328 ],
   alphaCSR[ 120 ][ 329 ],
   alphaCSR[ 120 ][ 330 ],
   alphaCSR[ 120 ][ 331 ],
   alphaCSR[ 120 ][ 332 ],
   alphaCSR[ 120 ][ 333 ],
   alphaCSR[ 120 ][ 334 ],
   alphaCSR[ 120 ][ 335 ],
   alphaCSR[ 120 ][ 336 ],
   alphaCSR[ 120 ][ 337 ],
   alphaCSR[ 120 ][ 338 ],
   alphaCSR[ 120 ][ 339 ],
   alphaCSR[ 120 ][ 340 ],
   alphaCSR[ 120 ][ 341 ],
   alphaCSR[ 120 ][ 342 ],
   alphaCSR[ 120 ][ 343 ],
   alphaCSR[ 120 ][ 344 ],
   alphaCSR[ 120 ][ 345 ],
   alphaCSR[ 120 ][ 346 ],
   alphaCSR[ 120 ][ 347 ],
   alphaCSR[ 120 ][ 348 ],
   alphaCSR[ 120 ][ 349 ],
   alphaCSR[ 120 ][ 350 ],
   alphaCSR[ 120 ][ 351 ],
   alphaCSR[ 120 ][ 352 ],
   alphaCSR[ 120 ][ 353 ],
   alphaCSR[ 120 ][ 354 ],
   alphaCSR[ 120 ][ 355 ],
   alphaCSR[ 120 ][ 356 ],
   alphaCSR[ 120 ][ 357 ],
   alphaCSR[ 120 ][ 358 ],
   alphaCSR[ 120 ][ 359 ],
   alphaCSR[ 120 ][ 360 ],
   alphaCSR[ 120 ][ 361 ],
   alphaCSR[ 120 ][ 362 ],
   alphaCSR[ 120 ][ 363 ],
   alphaCSR[ 120 ][ 364 ],
   alphaCSR[ 120 ][ 365 ],
   alphaCSR[ 120 ][ 366 ],
   alphaCSR[ 120 ][ 367 ],
   alphaCSR[ 120 ][ 368 ],
   alphaCSR[ 120 ][ 369 ],
   alphaCSR[ 120 ][ 370 ],
   alphaCSR[ 120 ][ 371 ],
   alphaCSR[ 120 ][ 372 ],
   alphaCSR[ 120 ][ 373 ],
   alphaCSR[ 120 ][ 374 ],
   alphaCSR[ 120 ][ 375 ],
   alphaCSR[ 120 ][ 376 ],
   alphaCSR[ 120 ][ 377 ],
   alphaCSR[ 120 ][ 378 ],
   alphaCSR[ 120 ][ 379 ],
   alphaCSR[ 120 ][ 380 ],
   alphaCSR[ 120 ][ 381 ],
   alphaCSR[ 120 ][ 382 ],
   alphaCSR[ 120 ][ 383 ],
   alphaCSR[ 121 ][ 0 ],
   alphaCSR[ 121 ][ 1 ],
   alphaCSR[ 121 ][ 2 ],
   alphaCSR[ 121 ][ 3 ],
   alphaCSR[ 121 ][ 4 ],
   alphaCSR[ 121 ][ 5 ],
   alphaCSR[ 121 ][ 6 ],
   alphaCSR[ 121 ][ 7 ],
   alphaCSR[ 121 ][ 8 ],
   alphaCSR[ 121 ][ 9 ],
   alphaCSR[ 121 ][ 10 ],
   alphaCSR[ 121 ][ 11 ],
   alphaCSR[ 121 ][ 12 ],
   alphaCSR[ 121 ][ 13 ],
   alphaCSR[ 121 ][ 14 ],
   alphaCSR[ 121 ][ 15 ],
   alphaCSR[ 121 ][ 16 ],
   alphaCSR[ 121 ][ 17 ],
   alphaCSR[ 121 ][ 18 ],
   alphaCSR[ 121 ][ 19 ],
   alphaCSR[ 121 ][ 20 ],
   alphaCSR[ 121 ][ 21 ],
   alphaCSR[ 121 ][ 22 ],
   alphaCSR[ 121 ][ 23 ],
   alphaCSR[ 121 ][ 24 ],
   alphaCSR[ 121 ][ 25 ],
   alphaCSR[ 121 ][ 26 ],
   alphaCSR[ 121 ][ 27 ],
   alphaCSR[ 121 ][ 28 ],
   alphaCSR[ 121 ][ 29 ],
   alphaCSR[ 121 ][ 30 ],
   alphaCSR[ 121 ][ 31 ],
   alphaCSR[ 121 ][ 32 ],
   alphaCSR[ 121 ][ 33 ],
   alphaCSR[ 121 ][ 34 ],
   alphaCSR[ 121 ][ 35 ],
   alphaCSR[ 121 ][ 36 ],
   alphaCSR[ 121 ][ 37 ],
   alphaCSR[ 121 ][ 38 ],
   alphaCSR[ 121 ][ 39 ],
   alphaCSR[ 121 ][ 40 ],
   alphaCSR[ 121 ][ 41 ],
   alphaCSR[ 121 ][ 42 ],
   alphaCSR[ 121 ][ 43 ],
   alphaCSR[ 121 ][ 44 ],
   alphaCSR[ 121 ][ 45 ],
   alphaCSR[ 121 ][ 46 ],
   alphaCSR[ 121 ][ 47 ],
   alphaCSR[ 121 ][ 48 ],
   alphaCSR[ 121 ][ 49 ],
   alphaCSR[ 121 ][ 50 ],
   alphaCSR[ 121 ][ 51 ],
   alphaCSR[ 121 ][ 52 ],
   alphaCSR[ 121 ][ 53 ],
   alphaCSR[ 121 ][ 54 ],
   alphaCSR[ 121 ][ 55 ],
   alphaCSR[ 121 ][ 56 ],
   alphaCSR[ 121 ][ 57 ],
   alphaCSR[ 121 ][ 58 ],
   alphaCSR[ 121 ][ 59 ],
   alphaCSR[ 121 ][ 60 ],
   alphaCSR[ 121 ][ 61 ],
   alphaCSR[ 121 ][ 62 ],
   alphaCSR[ 121 ][ 63 ],
   alphaCSR[ 121 ][ 64 ],
   alphaCSR[ 121 ][ 65 ],
   alphaCSR[ 121 ][ 66 ],
   alphaCSR[ 121 ][ 67 ],
   alphaCSR[ 121 ][ 68 ],
   alphaCSR[ 121 ][ 69 ],
   alphaCSR[ 121 ][ 70 ],
   alphaCSR[ 121 ][ 71 ],
   alphaCSR[ 121 ][ 72 ],
   alphaCSR[ 121 ][ 73 ],
   alphaCSR[ 121 ][ 74 ],
   alphaCSR[ 121 ][ 75 ],
   alphaCSR[ 121 ][ 76 ],
   alphaCSR[ 121 ][ 77 ],
   alphaCSR[ 121 ][ 78 ],
   alphaCSR[ 121 ][ 79 ],
   alphaCSR[ 121 ][ 80 ],
   alphaCSR[ 121 ][ 81 ],
   alphaCSR[ 121 ][ 82 ],
   alphaCSR[ 121 ][ 83 ],
   alphaCSR[ 121 ][ 84 ],
   alphaCSR[ 121 ][ 85 ],
   alphaCSR[ 121 ][ 86 ],
   alphaCSR[ 121 ][ 87 ],
   alphaCSR[ 121 ][ 88 ],
   alphaCSR[ 121 ][ 89 ],
   alphaCSR[ 121 ][ 90 ],
   alphaCSR[ 121 ][ 91 ],
   alphaCSR[ 121 ][ 92 ],
   alphaCSR[ 121 ][ 93 ],
   alphaCSR[ 121 ][ 94 ],
   alphaCSR[ 121 ][ 95 ],
   alphaCSR[ 121 ][ 96 ],
   alphaCSR[ 121 ][ 97 ],
   alphaCSR[ 121 ][ 98 ],
   alphaCSR[ 121 ][ 99 ],
   alphaCSR[ 121 ][ 100 ],
   alphaCSR[ 121 ][ 101 ],
   alphaCSR[ 121 ][ 102 ],
   alphaCSR[ 121 ][ 103 ],
   alphaCSR[ 121 ][ 104 ],
   alphaCSR[ 121 ][ 105 ],
   alphaCSR[ 121 ][ 106 ],
   alphaCSR[ 121 ][ 107 ],
   alphaCSR[ 121 ][ 108 ],
   alphaCSR[ 121 ][ 109 ],
   alphaCSR[ 121 ][ 110 ],
   alphaCSR[ 121 ][ 111 ],
   alphaCSR[ 121 ][ 112 ],
   alphaCSR[ 121 ][ 113 ],
   alphaCSR[ 121 ][ 114 ],
   alphaCSR[ 121 ][ 115 ],
   alphaCSR[ 121 ][ 116 ],
   alphaCSR[ 121 ][ 117 ],
   alphaCSR[ 121 ][ 118 ],
   alphaCSR[ 121 ][ 119 ],
   alphaCSR[ 121 ][ 120 ],
   alphaCSR[ 121 ][ 121 ],
   alphaCSR[ 121 ][ 122 ],
   alphaCSR[ 121 ][ 123 ],
   alphaCSR[ 121 ][ 124 ],
   alphaCSR[ 121 ][ 125 ],
   alphaCSR[ 121 ][ 126 ],
   alphaCSR[ 121 ][ 127 ],
   alphaCSR[ 121 ][ 128 ],
   alphaCSR[ 121 ][ 129 ],
   alphaCSR[ 121 ][ 130 ],
   alphaCSR[ 121 ][ 131 ],
   alphaCSR[ 121 ][ 132 ],
   alphaCSR[ 121 ][ 133 ],
   alphaCSR[ 121 ][ 134 ],
   alphaCSR[ 121 ][ 135 ],
   alphaCSR[ 121 ][ 136 ],
   alphaCSR[ 121 ][ 137 ],
   alphaCSR[ 121 ][ 138 ],
   alphaCSR[ 121 ][ 139 ],
   alphaCSR[ 121 ][ 140 ],
   alphaCSR[ 121 ][ 141 ],
   alphaCSR[ 121 ][ 142 ],
   alphaCSR[ 121 ][ 143 ],
   alphaCSR[ 121 ][ 144 ],
   alphaCSR[ 121 ][ 145 ],
   alphaCSR[ 121 ][ 146 ],
   alphaCSR[ 121 ][ 147 ],
   alphaCSR[ 121 ][ 148 ],
   alphaCSR[ 121 ][ 149 ],
   alphaCSR[ 121 ][ 150 ],
   alphaCSR[ 121 ][ 151 ],
   alphaCSR[ 121 ][ 152 ],
   alphaCSR[ 121 ][ 153 ],
   alphaCSR[ 121 ][ 154 ],
   alphaCSR[ 121 ][ 155 ],
   alphaCSR[ 121 ][ 156 ],
   alphaCSR[ 121 ][ 157 ],
   alphaCSR[ 121 ][ 158 ],
   alphaCSR[ 121 ][ 159 ],
   alphaCSR[ 121 ][ 160 ],
   alphaCSR[ 121 ][ 161 ],
   alphaCSR[ 121 ][ 162 ],
   alphaCSR[ 121 ][ 163 ],
   alphaCSR[ 121 ][ 164 ],
   alphaCSR[ 121 ][ 165 ],
   alphaCSR[ 121 ][ 166 ],
   alphaCSR[ 121 ][ 167 ],
   alphaCSR[ 121 ][ 168 ],
   alphaCSR[ 121 ][ 169 ],
   alphaCSR[ 121 ][ 170 ],
   alphaCSR[ 121 ][ 171 ],
   alphaCSR[ 121 ][ 172 ],
   alphaCSR[ 121 ][ 173 ],
   alphaCSR[ 121 ][ 174 ],
   alphaCSR[ 121 ][ 175 ],
   alphaCSR[ 121 ][ 176 ],
   alphaCSR[ 121 ][ 177 ],
   alphaCSR[ 121 ][ 178 ],
   alphaCSR[ 121 ][ 179 ],
   alphaCSR[ 121 ][ 180 ],
   alphaCSR[ 121 ][ 181 ],
   alphaCSR[ 121 ][ 182 ],
   alphaCSR[ 121 ][ 183 ],
   alphaCSR[ 121 ][ 184 ],
   alphaCSR[ 121 ][ 185 ],
   alphaCSR[ 121 ][ 186 ],
   alphaCSR[ 121 ][ 187 ],
   alphaCSR[ 121 ][ 188 ],
   alphaCSR[ 121 ][ 189 ],
   alphaCSR[ 121 ][ 190 ],
   alphaCSR[ 121 ][ 191 ],
   alphaCSR[ 121 ][ 192 ],
   alphaCSR[ 121 ][ 193 ],
   alphaCSR[ 121 ][ 194 ],
   alphaCSR[ 121 ][ 195 ],
   alphaCSR[ 121 ][ 196 ],
   alphaCSR[ 121 ][ 197 ],
   alphaCSR[ 121 ][ 198 ],
   alphaCSR[ 121 ][ 199 ],
   alphaCSR[ 121 ][ 200 ],
   alphaCSR[ 121 ][ 201 ],
   alphaCSR[ 121 ][ 202 ],
   alphaCSR[ 121 ][ 203 ],
   alphaCSR[ 121 ][ 204 ],
   alphaCSR[ 121 ][ 205 ],
   alphaCSR[ 121 ][ 206 ],
   alphaCSR[ 121 ][ 207 ],
   alphaCSR[ 121 ][ 208 ],
   alphaCSR[ 121 ][ 209 ],
   alphaCSR[ 121 ][ 210 ],
   alphaCSR[ 121 ][ 211 ],
   alphaCSR[ 121 ][ 212 ],
   alphaCSR[ 121 ][ 213 ],
   alphaCSR[ 121 ][ 214 ],
   alphaCSR[ 121 ][ 215 ],
   alphaCSR[ 121 ][ 216 ],
   alphaCSR[ 121 ][ 217 ],
   alphaCSR[ 121 ][ 218 ],
   alphaCSR[ 121 ][ 219 ],
   alphaCSR[ 121 ][ 220 ],
   alphaCSR[ 121 ][ 221 ],
   alphaCSR[ 121 ][ 222 ],
   alphaCSR[ 121 ][ 223 ],
   alphaCSR[ 121 ][ 224 ],
   alphaCSR[ 121 ][ 225 ],
   alphaCSR[ 121 ][ 226 ],
   alphaCSR[ 121 ][ 227 ],
   alphaCSR[ 121 ][ 228 ],
   alphaCSR[ 121 ][ 229 ],
   alphaCSR[ 121 ][ 230 ],
   alphaCSR[ 121 ][ 231 ],
   alphaCSR[ 121 ][ 232 ],
   alphaCSR[ 121 ][ 233 ],
   alphaCSR[ 121 ][ 234 ],
   alphaCSR[ 121 ][ 235 ],
   alphaCSR[ 121 ][ 236 ],
   alphaCSR[ 121 ][ 237 ],
   alphaCSR[ 121 ][ 238 ],
   alphaCSR[ 121 ][ 239 ],
   alphaCSR[ 121 ][ 240 ],
   alphaCSR[ 121 ][ 241 ],
   alphaCSR[ 121 ][ 242 ],
   alphaCSR[ 121 ][ 243 ],
   alphaCSR[ 121 ][ 244 ],
   alphaCSR[ 121 ][ 245 ],
   alphaCSR[ 121 ][ 246 ],
   alphaCSR[ 121 ][ 247 ],
   alphaCSR[ 121 ][ 248 ],
   alphaCSR[ 121 ][ 249 ],
   alphaCSR[ 121 ][ 250 ],
   alphaCSR[ 121 ][ 251 ],
   alphaCSR[ 121 ][ 252 ],
   alphaCSR[ 121 ][ 253 ],
   alphaCSR[ 121 ][ 254 ],
   alphaCSR[ 121 ][ 255 ],
   alphaCSR[ 121 ][ 256 ],
   alphaCSR[ 121 ][ 257 ],
   alphaCSR[ 121 ][ 258 ],
   alphaCSR[ 121 ][ 259 ],
   alphaCSR[ 121 ][ 260 ],
   alphaCSR[ 121 ][ 261 ],
   alphaCSR[ 121 ][ 262 ],
   alphaCSR[ 121 ][ 263 ],
   alphaCSR[ 121 ][ 264 ],
   alphaCSR[ 121 ][ 265 ],
   alphaCSR[ 121 ][ 266 ],
   alphaCSR[ 121 ][ 267 ],
   alphaCSR[ 121 ][ 268 ],
   alphaCSR[ 121 ][ 269 ],
   alphaCSR[ 121 ][ 270 ],
   alphaCSR[ 121 ][ 271 ],
   alphaCSR[ 121 ][ 272 ],
   alphaCSR[ 121 ][ 273 ],
   alphaCSR[ 121 ][ 274 ],
   alphaCSR[ 121 ][ 275 ],
   alphaCSR[ 121 ][ 276 ],
   alphaCSR[ 121 ][ 277 ],
   alphaCSR[ 121 ][ 278 ],
   alphaCSR[ 121 ][ 279 ],
   alphaCSR[ 121 ][ 280 ],
   alphaCSR[ 121 ][ 281 ],
   alphaCSR[ 121 ][ 282 ],
   alphaCSR[ 121 ][ 283 ],
   alphaCSR[ 121 ][ 284 ],
   alphaCSR[ 121 ][ 285 ],
   alphaCSR[ 121 ][ 286 ],
   alphaCSR[ 121 ][ 287 ],
   alphaCSR[ 121 ][ 288 ],
   alphaCSR[ 121 ][ 289 ],
   alphaCSR[ 121 ][ 290 ],
   alphaCSR[ 121 ][ 291 ],
   alphaCSR[ 121 ][ 292 ],
   alphaCSR[ 121 ][ 293 ],
   alphaCSR[ 121 ][ 294 ],
   alphaCSR[ 121 ][ 295 ],
   alphaCSR[ 121 ][ 296 ],
   alphaCSR[ 121 ][ 297 ],
   alphaCSR[ 121 ][ 298 ],
   alphaCSR[ 121 ][ 299 ],
   alphaCSR[ 121 ][ 300 ],
   alphaCSR[ 121 ][ 301 ],
   alphaCSR[ 121 ][ 302 ],
   alphaCSR[ 121 ][ 303 ],
   alphaCSR[ 121 ][ 304 ],
   alphaCSR[ 121 ][ 305 ],
   alphaCSR[ 121 ][ 306 ],
   alphaCSR[ 121 ][ 307 ],
   alphaCSR[ 121 ][ 308 ],
   alphaCSR[ 121 ][ 309 ],
   alphaCSR[ 121 ][ 310 ],
   alphaCSR[ 121 ][ 311 ],
   alphaCSR[ 121 ][ 312 ],
   alphaCSR[ 121 ][ 313 ],
   alphaCSR[ 121 ][ 314 ],
   alphaCSR[ 121 ][ 315 ],
   alphaCSR[ 121 ][ 316 ],
   alphaCSR[ 121 ][ 317 ],
   alphaCSR[ 121 ][ 318 ],
   alphaCSR[ 121 ][ 319 ],
   alphaCSR[ 121 ][ 320 ],
   alphaCSR[ 121 ][ 321 ],
   alphaCSR[ 121 ][ 322 ],
   alphaCSR[ 121 ][ 323 ],
   alphaCSR[ 121 ][ 324 ],
   alphaCSR[ 121 ][ 325 ],
   alphaCSR[ 121 ][ 326 ],
   alphaCSR[ 121 ][ 327 ],
   alphaCSR[ 121 ][ 328 ],
   alphaCSR[ 121 ][ 329 ],
   alphaCSR[ 121 ][ 330 ],
   alphaCSR[ 121 ][ 331 ],
   alphaCSR[ 121 ][ 332 ],
   alphaCSR[ 121 ][ 333 ],
   alphaCSR[ 121 ][ 334 ],
   alphaCSR[ 121 ][ 335 ],
   alphaCSR[ 121 ][ 336 ],
   alphaCSR[ 121 ][ 337 ],
   alphaCSR[ 121 ][ 338 ],
   alphaCSR[ 121 ][ 339 ],
   alphaCSR[ 121 ][ 340 ],
   alphaCSR[ 121 ][ 341 ],
   alphaCSR[ 121 ][ 342 ],
   alphaCSR[ 121 ][ 343 ],
   alphaCSR[ 121 ][ 344 ],
   alphaCSR[ 121 ][ 345 ],
   alphaCSR[ 121 ][ 346 ],
   alphaCSR[ 121 ][ 347 ],
   alphaCSR[ 121 ][ 348 ],
   alphaCSR[ 121 ][ 349 ],
   alphaCSR[ 121 ][ 350 ],
   alphaCSR[ 121 ][ 351 ],
   alphaCSR[ 121 ][ 352 ],
   alphaCSR[ 121 ][ 353 ],
   alphaCSR[ 121 ][ 354 ],
   alphaCSR[ 121 ][ 355 ],
   alphaCSR[ 121 ][ 356 ],
   alphaCSR[ 121 ][ 357 ],
   alphaCSR[ 121 ][ 358 ],
   alphaCSR[ 121 ][ 359 ],
   alphaCSR[ 121 ][ 360 ],
   alphaCSR[ 121 ][ 361 ],
   alphaCSR[ 121 ][ 362 ],
   alphaCSR[ 121 ][ 363 ],
   alphaCSR[ 121 ][ 364 ],
   alphaCSR[ 121 ][ 365 ],
   alphaCSR[ 121 ][ 366 ],
   alphaCSR[ 121 ][ 367 ],
   alphaCSR[ 121 ][ 368 ],
   alphaCSR[ 121 ][ 369 ],
   alphaCSR[ 121 ][ 370 ],
   alphaCSR[ 121 ][ 371 ],
   alphaCSR[ 121 ][ 372 ],
   alphaCSR[ 121 ][ 373 ],
   alphaCSR[ 121 ][ 374 ],
   alphaCSR[ 121 ][ 375 ],
   alphaCSR[ 121 ][ 376 ],
   alphaCSR[ 121 ][ 377 ],
   alphaCSR[ 121 ][ 378 ],
   alphaCSR[ 121 ][ 379 ],
   alphaCSR[ 121 ][ 380 ],
   alphaCSR[ 121 ][ 381 ],
   alphaCSR[ 121 ][ 382 ],
   alphaCSR[ 121 ][ 383 ],
   alphaCSR[ 122 ][ 0 ],
   alphaCSR[ 122 ][ 1 ],
   alphaCSR[ 122 ][ 2 ],
   alphaCSR[ 122 ][ 3 ],
   alphaCSR[ 122 ][ 4 ],
   alphaCSR[ 122 ][ 5 ],
   alphaCSR[ 122 ][ 6 ],
   alphaCSR[ 122 ][ 7 ],
   alphaCSR[ 122 ][ 8 ],
   alphaCSR[ 122 ][ 9 ],
   alphaCSR[ 122 ][ 10 ],
   alphaCSR[ 122 ][ 11 ],
   alphaCSR[ 122 ][ 12 ],
   alphaCSR[ 122 ][ 13 ],
   alphaCSR[ 122 ][ 14 ],
   alphaCSR[ 122 ][ 15 ],
   alphaCSR[ 122 ][ 16 ],
   alphaCSR[ 122 ][ 17 ],
   alphaCSR[ 122 ][ 18 ],
   alphaCSR[ 122 ][ 19 ],
   alphaCSR[ 122 ][ 20 ],
   alphaCSR[ 122 ][ 21 ],
   alphaCSR[ 122 ][ 22 ],
   alphaCSR[ 122 ][ 23 ],
   alphaCSR[ 122 ][ 24 ],
   alphaCSR[ 122 ][ 25 ],
   alphaCSR[ 122 ][ 26 ],
   alphaCSR[ 122 ][ 27 ],
   alphaCSR[ 122 ][ 28 ],
   alphaCSR[ 122 ][ 29 ],
   alphaCSR[ 122 ][ 30 ],
   alphaCSR[ 122 ][ 31 ],
   alphaCSR[ 122 ][ 32 ],
   alphaCSR[ 122 ][ 33 ],
   alphaCSR[ 122 ][ 34 ],
   alphaCSR[ 122 ][ 35 ],
   alphaCSR[ 122 ][ 36 ],
   alphaCSR[ 122 ][ 37 ],
   alphaCSR[ 122 ][ 38 ],
   alphaCSR[ 122 ][ 39 ],
   alphaCSR[ 122 ][ 40 ],
   alphaCSR[ 122 ][ 41 ],
   alphaCSR[ 122 ][ 42 ],
   alphaCSR[ 122 ][ 43 ],
   alphaCSR[ 122 ][ 44 ],
   alphaCSR[ 122 ][ 45 ],
   alphaCSR[ 122 ][ 46 ],
   alphaCSR[ 122 ][ 47 ],
   alphaCSR[ 122 ][ 48 ],
   alphaCSR[ 122 ][ 49 ],
   alphaCSR[ 122 ][ 50 ],
   alphaCSR[ 122 ][ 51 ],
   alphaCSR[ 122 ][ 52 ],
   alphaCSR[ 122 ][ 53 ],
   alphaCSR[ 122 ][ 54 ],
   alphaCSR[ 122 ][ 55 ],
   alphaCSR[ 122 ][ 56 ],
   alphaCSR[ 122 ][ 57 ],
   alphaCSR[ 122 ][ 58 ],
   alphaCSR[ 122 ][ 59 ],
   alphaCSR[ 122 ][ 60 ],
   alphaCSR[ 122 ][ 61 ],
   alphaCSR[ 122 ][ 62 ],
   alphaCSR[ 122 ][ 63 ],
   alphaCSR[ 122 ][ 64 ],
   alphaCSR[ 122 ][ 65 ],
   alphaCSR[ 122 ][ 66 ],
   alphaCSR[ 122 ][ 67 ],
   alphaCSR[ 122 ][ 68 ],
   alphaCSR[ 122 ][ 69 ],
   alphaCSR[ 122 ][ 70 ],
   alphaCSR[ 122 ][ 71 ],
   alphaCSR[ 122 ][ 72 ],
   alphaCSR[ 122 ][ 73 ],
   alphaCSR[ 122 ][ 74 ],
   alphaCSR[ 122 ][ 75 ],
   alphaCSR[ 122 ][ 76 ],
   alphaCSR[ 122 ][ 77 ],
   alphaCSR[ 122 ][ 78 ],
   alphaCSR[ 122 ][ 79 ],
   alphaCSR[ 122 ][ 80 ],
   alphaCSR[ 122 ][ 81 ],
   alphaCSR[ 122 ][ 82 ],
   alphaCSR[ 122 ][ 83 ],
   alphaCSR[ 122 ][ 84 ],
   alphaCSR[ 122 ][ 85 ],
   alphaCSR[ 122 ][ 86 ],
   alphaCSR[ 122 ][ 87 ],
   alphaCSR[ 122 ][ 88 ],
   alphaCSR[ 122 ][ 89 ],
   alphaCSR[ 122 ][ 90 ],
   alphaCSR[ 122 ][ 91 ],
   alphaCSR[ 122 ][ 92 ],
   alphaCSR[ 122 ][ 93 ],
   alphaCSR[ 122 ][ 94 ],
   alphaCSR[ 122 ][ 95 ],
   alphaCSR[ 122 ][ 96 ],
   alphaCSR[ 122 ][ 97 ],
   alphaCSR[ 122 ][ 98 ],
   alphaCSR[ 122 ][ 99 ],
   alphaCSR[ 122 ][ 100 ],
   alphaCSR[ 122 ][ 101 ],
   alphaCSR[ 122 ][ 102 ],
   alphaCSR[ 122 ][ 103 ],
   alphaCSR[ 122 ][ 104 ],
   alphaCSR[ 122 ][ 105 ],
   alphaCSR[ 122 ][ 106 ],
   alphaCSR[ 122 ][ 107 ],
   alphaCSR[ 122 ][ 108 ],
   alphaCSR[ 122 ][ 109 ],
   alphaCSR[ 122 ][ 110 ],
   alphaCSR[ 122 ][ 111 ],
   alphaCSR[ 122 ][ 112 ],
   alphaCSR[ 122 ][ 113 ],
   alphaCSR[ 122 ][ 114 ],
   alphaCSR[ 122 ][ 115 ],
   alphaCSR[ 122 ][ 116 ],
   alphaCSR[ 122 ][ 117 ],
   alphaCSR[ 122 ][ 118 ],
   alphaCSR[ 122 ][ 119 ],
   alphaCSR[ 122 ][ 120 ],
   alphaCSR[ 122 ][ 121 ],
   alphaCSR[ 122 ][ 122 ],
   alphaCSR[ 122 ][ 123 ],
   alphaCSR[ 122 ][ 124 ],
   alphaCSR[ 122 ][ 125 ],
   alphaCSR[ 122 ][ 126 ],
   alphaCSR[ 122 ][ 127 ],
   alphaCSR[ 122 ][ 128 ],
   alphaCSR[ 122 ][ 129 ],
   alphaCSR[ 122 ][ 130 ],
   alphaCSR[ 122 ][ 131 ],
   alphaCSR[ 122 ][ 132 ],
   alphaCSR[ 122 ][ 133 ],
   alphaCSR[ 122 ][ 134 ],
   alphaCSR[ 122 ][ 135 ],
   alphaCSR[ 122 ][ 136 ],
   alphaCSR[ 122 ][ 137 ],
   alphaCSR[ 122 ][ 138 ],
   alphaCSR[ 122 ][ 139 ],
   alphaCSR[ 122 ][ 140 ],
   alphaCSR[ 122 ][ 141 ],
   alphaCSR[ 122 ][ 142 ],
   alphaCSR[ 122 ][ 143 ],
   alphaCSR[ 122 ][ 144 ],
   alphaCSR[ 122 ][ 145 ],
   alphaCSR[ 122 ][ 146 ],
   alphaCSR[ 122 ][ 147 ],
   alphaCSR[ 122 ][ 148 ],
   alphaCSR[ 122 ][ 149 ],
   alphaCSR[ 122 ][ 150 ],
   alphaCSR[ 122 ][ 151 ],
   alphaCSR[ 122 ][ 152 ],
   alphaCSR[ 122 ][ 153 ],
   alphaCSR[ 122 ][ 154 ],
   alphaCSR[ 122 ][ 155 ],
   alphaCSR[ 122 ][ 156 ],
   alphaCSR[ 122 ][ 157 ],
   alphaCSR[ 122 ][ 158 ],
   alphaCSR[ 122 ][ 159 ],
   alphaCSR[ 122 ][ 160 ],
   alphaCSR[ 122 ][ 161 ],
   alphaCSR[ 122 ][ 162 ],
   alphaCSR[ 122 ][ 163 ],
   alphaCSR[ 122 ][ 164 ],
   alphaCSR[ 122 ][ 165 ],
   alphaCSR[ 122 ][ 166 ],
   alphaCSR[ 122 ][ 167 ],
   alphaCSR[ 122 ][ 168 ],
   alphaCSR[ 122 ][ 169 ],
   alphaCSR[ 122 ][ 170 ],
   alphaCSR[ 122 ][ 171 ],
   alphaCSR[ 122 ][ 172 ],
   alphaCSR[ 122 ][ 173 ],
   alphaCSR[ 122 ][ 174 ],
   alphaCSR[ 122 ][ 175 ],
   alphaCSR[ 122 ][ 176 ],
   alphaCSR[ 122 ][ 177 ],
   alphaCSR[ 122 ][ 178 ],
   alphaCSR[ 122 ][ 179 ],
   alphaCSR[ 122 ][ 180 ],
   alphaCSR[ 122 ][ 181 ],
   alphaCSR[ 122 ][ 182 ],
   alphaCSR[ 122 ][ 183 ],
   alphaCSR[ 122 ][ 184 ],
   alphaCSR[ 122 ][ 185 ],
   alphaCSR[ 122 ][ 186 ],
   alphaCSR[ 122 ][ 187 ],
   alphaCSR[ 122 ][ 188 ],
   alphaCSR[ 122 ][ 189 ],
   alphaCSR[ 122 ][ 190 ],
   alphaCSR[ 122 ][ 191 ],
   alphaCSR[ 122 ][ 192 ],
   alphaCSR[ 122 ][ 193 ],
   alphaCSR[ 122 ][ 194 ],
   alphaCSR[ 122 ][ 195 ],
   alphaCSR[ 122 ][ 196 ],
   alphaCSR[ 122 ][ 197 ],
   alphaCSR[ 122 ][ 198 ],
   alphaCSR[ 122 ][ 199 ],
   alphaCSR[ 122 ][ 200 ],
   alphaCSR[ 122 ][ 201 ],
   alphaCSR[ 122 ][ 202 ],
   alphaCSR[ 122 ][ 203 ],
   alphaCSR[ 122 ][ 204 ],
   alphaCSR[ 122 ][ 205 ],
   alphaCSR[ 122 ][ 206 ],
   alphaCSR[ 122 ][ 207 ],
   alphaCSR[ 122 ][ 208 ],
   alphaCSR[ 122 ][ 209 ],
   alphaCSR[ 122 ][ 210 ],
   alphaCSR[ 122 ][ 211 ],
   alphaCSR[ 122 ][ 212 ],
   alphaCSR[ 122 ][ 213 ],
   alphaCSR[ 122 ][ 214 ],
   alphaCSR[ 122 ][ 215 ],
   alphaCSR[ 122 ][ 216 ],
   alphaCSR[ 122 ][ 217 ],
   alphaCSR[ 122 ][ 218 ],
   alphaCSR[ 122 ][ 219 ],
   alphaCSR[ 122 ][ 220 ],
   alphaCSR[ 122 ][ 221 ],
   alphaCSR[ 122 ][ 222 ],
   alphaCSR[ 122 ][ 223 ],
   alphaCSR[ 122 ][ 224 ],
   alphaCSR[ 122 ][ 225 ],
   alphaCSR[ 122 ][ 226 ],
   alphaCSR[ 122 ][ 227 ],
   alphaCSR[ 122 ][ 228 ],
   alphaCSR[ 122 ][ 229 ],
   alphaCSR[ 122 ][ 230 ],
   alphaCSR[ 122 ][ 231 ],
   alphaCSR[ 122 ][ 232 ],
   alphaCSR[ 122 ][ 233 ],
   alphaCSR[ 122 ][ 234 ],
   alphaCSR[ 122 ][ 235 ],
   alphaCSR[ 122 ][ 236 ],
   alphaCSR[ 122 ][ 237 ],
   alphaCSR[ 122 ][ 238 ],
   alphaCSR[ 122 ][ 239 ],
   alphaCSR[ 122 ][ 240 ],
   alphaCSR[ 122 ][ 241 ],
   alphaCSR[ 122 ][ 242 ],
   alphaCSR[ 122 ][ 243 ],
   alphaCSR[ 122 ][ 244 ],
   alphaCSR[ 122 ][ 245 ],
   alphaCSR[ 122 ][ 246 ],
   alphaCSR[ 122 ][ 247 ],
   alphaCSR[ 122 ][ 248 ],
   alphaCSR[ 122 ][ 249 ],
   alphaCSR[ 122 ][ 250 ],
   alphaCSR[ 122 ][ 251 ],
   alphaCSR[ 122 ][ 252 ],
   alphaCSR[ 122 ][ 253 ],
   alphaCSR[ 122 ][ 254 ],
   alphaCSR[ 122 ][ 255 ],
   alphaCSR[ 122 ][ 256 ],
   alphaCSR[ 122 ][ 257 ],
   alphaCSR[ 122 ][ 258 ],
   alphaCSR[ 122 ][ 259 ],
   alphaCSR[ 122 ][ 260 ],
   alphaCSR[ 122 ][ 261 ],
   alphaCSR[ 122 ][ 262 ],
   alphaCSR[ 122 ][ 263 ],
   alphaCSR[ 122 ][ 264 ],
   alphaCSR[ 122 ][ 265 ],
   alphaCSR[ 122 ][ 266 ],
   alphaCSR[ 122 ][ 267 ],
   alphaCSR[ 122 ][ 268 ],
   alphaCSR[ 122 ][ 269 ],
   alphaCSR[ 122 ][ 270 ],
   alphaCSR[ 122 ][ 271 ],
   alphaCSR[ 122 ][ 272 ],
   alphaCSR[ 122 ][ 273 ],
   alphaCSR[ 122 ][ 274 ],
   alphaCSR[ 122 ][ 275 ],
   alphaCSR[ 122 ][ 276 ],
   alphaCSR[ 122 ][ 277 ],
   alphaCSR[ 122 ][ 278 ],
   alphaCSR[ 122 ][ 279 ],
   alphaCSR[ 122 ][ 280 ],
   alphaCSR[ 122 ][ 281 ],
   alphaCSR[ 122 ][ 282 ],
   alphaCSR[ 122 ][ 283 ],
   alphaCSR[ 122 ][ 284 ],
   alphaCSR[ 122 ][ 285 ],
   alphaCSR[ 122 ][ 286 ],
   alphaCSR[ 122 ][ 287 ],
   alphaCSR[ 122 ][ 288 ],
   alphaCSR[ 122 ][ 289 ],
   alphaCSR[ 122 ][ 290 ],
   alphaCSR[ 122 ][ 291 ],
   alphaCSR[ 122 ][ 292 ],
   alphaCSR[ 122 ][ 293 ],
   alphaCSR[ 122 ][ 294 ],
   alphaCSR[ 122 ][ 295 ],
   alphaCSR[ 122 ][ 296 ],
   alphaCSR[ 122 ][ 297 ],
   alphaCSR[ 122 ][ 298 ],
   alphaCSR[ 122 ][ 299 ],
   alphaCSR[ 122 ][ 300 ],
   alphaCSR[ 122 ][ 301 ],
   alphaCSR[ 122 ][ 302 ],
   alphaCSR[ 122 ][ 303 ],
   alphaCSR[ 122 ][ 304 ],
   alphaCSR[ 122 ][ 305 ],
   alphaCSR[ 122 ][ 306 ],
   alphaCSR[ 122 ][ 307 ],
   alphaCSR[ 122 ][ 308 ],
   alphaCSR[ 122 ][ 309 ],
   alphaCSR[ 122 ][ 310 ],
   alphaCSR[ 122 ][ 311 ],
   alphaCSR[ 122 ][ 312 ],
   alphaCSR[ 122 ][ 313 ],
   alphaCSR[ 122 ][ 314 ],
   alphaCSR[ 122 ][ 315 ],
   alphaCSR[ 122 ][ 316 ],
   alphaCSR[ 122 ][ 317 ],
   alphaCSR[ 122 ][ 318 ],
   alphaCSR[ 122 ][ 319 ],
   alphaCSR[ 122 ][ 320 ],
   alphaCSR[ 122 ][ 321 ],
   alphaCSR[ 122 ][ 322 ],
   alphaCSR[ 122 ][ 323 ],
   alphaCSR[ 122 ][ 324 ],
   alphaCSR[ 122 ][ 325 ],
   alphaCSR[ 122 ][ 326 ],
   alphaCSR[ 122 ][ 327 ],
   alphaCSR[ 122 ][ 328 ],
   alphaCSR[ 122 ][ 329 ],
   alphaCSR[ 122 ][ 330 ],
   alphaCSR[ 122 ][ 331 ],
   alphaCSR[ 122 ][ 332 ],
   alphaCSR[ 122 ][ 333 ],
   alphaCSR[ 122 ][ 334 ],
   alphaCSR[ 122 ][ 335 ],
   alphaCSR[ 122 ][ 336 ],
   alphaCSR[ 122 ][ 337 ],
   alphaCSR[ 122 ][ 338 ],
   alphaCSR[ 122 ][ 339 ],
   alphaCSR[ 122 ][ 340 ],
   alphaCSR[ 122 ][ 341 ],
   alphaCSR[ 122 ][ 342 ],
   alphaCSR[ 122 ][ 343 ],
   alphaCSR[ 122 ][ 344 ],
   alphaCSR[ 122 ][ 345 ],
   alphaCSR[ 122 ][ 346 ],
   alphaCSR[ 122 ][ 347 ],
   alphaCSR[ 122 ][ 348 ],
   alphaCSR[ 122 ][ 349 ],
   alphaCSR[ 122 ][ 350 ],
   alphaCSR[ 122 ][ 351 ],
   alphaCSR[ 122 ][ 352 ],
   alphaCSR[ 122 ][ 353 ],
   alphaCSR[ 122 ][ 354 ],
   alphaCSR[ 122 ][ 355 ],
   alphaCSR[ 122 ][ 356 ],
   alphaCSR[ 122 ][ 357 ],
   alphaCSR[ 122 ][ 358 ],
   alphaCSR[ 122 ][ 359 ],
   alphaCSR[ 122 ][ 360 ],
   alphaCSR[ 122 ][ 361 ],
   alphaCSR[ 122 ][ 362 ],
   alphaCSR[ 122 ][ 363 ],
   alphaCSR[ 122 ][ 364 ],
   alphaCSR[ 122 ][ 365 ],
   alphaCSR[ 122 ][ 366 ],
   alphaCSR[ 122 ][ 367 ],
   alphaCSR[ 122 ][ 368 ],
   alphaCSR[ 122 ][ 369 ],
   alphaCSR[ 122 ][ 370 ],
   alphaCSR[ 122 ][ 371 ],
   alphaCSR[ 122 ][ 372 ],
   alphaCSR[ 122 ][ 373 ],
   alphaCSR[ 122 ][ 374 ],
   alphaCSR[ 122 ][ 375 ],
   alphaCSR[ 122 ][ 376 ],
   alphaCSR[ 122 ][ 377 ],
   alphaCSR[ 122 ][ 378 ],
   alphaCSR[ 122 ][ 379 ],
   alphaCSR[ 122 ][ 380 ],
   alphaCSR[ 122 ][ 381 ],
   alphaCSR[ 122 ][ 382 ],
   alphaCSR[ 122 ][ 383 ],
   alphaCSR[ 123 ][ 0 ],
   alphaCSR[ 123 ][ 1 ],
   alphaCSR[ 123 ][ 2 ],
   alphaCSR[ 123 ][ 3 ],
   alphaCSR[ 123 ][ 4 ],
   alphaCSR[ 123 ][ 5 ],
   alphaCSR[ 123 ][ 6 ],
   alphaCSR[ 123 ][ 7 ],
   alphaCSR[ 123 ][ 8 ],
   alphaCSR[ 123 ][ 9 ],
   alphaCSR[ 123 ][ 10 ],
   alphaCSR[ 123 ][ 11 ],
   alphaCSR[ 123 ][ 12 ],
   alphaCSR[ 123 ][ 13 ],
   alphaCSR[ 123 ][ 14 ],
   alphaCSR[ 123 ][ 15 ],
   alphaCSR[ 123 ][ 16 ],
   alphaCSR[ 123 ][ 17 ],
   alphaCSR[ 123 ][ 18 ],
   alphaCSR[ 123 ][ 19 ],
   alphaCSR[ 123 ][ 20 ],
   alphaCSR[ 123 ][ 21 ],
   alphaCSR[ 123 ][ 22 ],
   alphaCSR[ 123 ][ 23 ],
   alphaCSR[ 123 ][ 24 ],
   alphaCSR[ 123 ][ 25 ],
   alphaCSR[ 123 ][ 26 ],
   alphaCSR[ 123 ][ 27 ],
   alphaCSR[ 123 ][ 28 ],
   alphaCSR[ 123 ][ 29 ],
   alphaCSR[ 123 ][ 30 ],
   alphaCSR[ 123 ][ 31 ],
   alphaCSR[ 123 ][ 32 ],
   alphaCSR[ 123 ][ 33 ],
   alphaCSR[ 123 ][ 34 ],
   alphaCSR[ 123 ][ 35 ],
   alphaCSR[ 123 ][ 36 ],
   alphaCSR[ 123 ][ 37 ],
   alphaCSR[ 123 ][ 38 ],
   alphaCSR[ 123 ][ 39 ],
   alphaCSR[ 123 ][ 40 ],
   alphaCSR[ 123 ][ 41 ],
   alphaCSR[ 123 ][ 42 ],
   alphaCSR[ 123 ][ 43 ],
   alphaCSR[ 123 ][ 44 ],
   alphaCSR[ 123 ][ 45 ],
   alphaCSR[ 123 ][ 46 ],
   alphaCSR[ 123 ][ 47 ],
   alphaCSR[ 123 ][ 48 ],
   alphaCSR[ 123 ][ 49 ],
   alphaCSR[ 123 ][ 50 ],
   alphaCSR[ 123 ][ 51 ],
   alphaCSR[ 123 ][ 52 ],
   alphaCSR[ 123 ][ 53 ],
   alphaCSR[ 123 ][ 54 ],
   alphaCSR[ 123 ][ 55 ],
   alphaCSR[ 123 ][ 56 ],
   alphaCSR[ 123 ][ 57 ],
   alphaCSR[ 123 ][ 58 ],
   alphaCSR[ 123 ][ 59 ],
   alphaCSR[ 123 ][ 60 ],
   alphaCSR[ 123 ][ 61 ],
   alphaCSR[ 123 ][ 62 ],
   alphaCSR[ 123 ][ 63 ],
   alphaCSR[ 123 ][ 64 ],
   alphaCSR[ 123 ][ 65 ],
   alphaCSR[ 123 ][ 66 ],
   alphaCSR[ 123 ][ 67 ],
   alphaCSR[ 123 ][ 68 ],
   alphaCSR[ 123 ][ 69 ],
   alphaCSR[ 123 ][ 70 ],
   alphaCSR[ 123 ][ 71 ],
   alphaCSR[ 123 ][ 72 ],
   alphaCSR[ 123 ][ 73 ],
   alphaCSR[ 123 ][ 74 ],
   alphaCSR[ 123 ][ 75 ],
   alphaCSR[ 123 ][ 76 ],
   alphaCSR[ 123 ][ 77 ],
   alphaCSR[ 123 ][ 78 ],
   alphaCSR[ 123 ][ 79 ],
   alphaCSR[ 123 ][ 80 ],
   alphaCSR[ 123 ][ 81 ],
   alphaCSR[ 123 ][ 82 ],
   alphaCSR[ 123 ][ 83 ],
   alphaCSR[ 123 ][ 84 ],
   alphaCSR[ 123 ][ 85 ],
   alphaCSR[ 123 ][ 86 ],
   alphaCSR[ 123 ][ 87 ],
   alphaCSR[ 123 ][ 88 ],
   alphaCSR[ 123 ][ 89 ],
   alphaCSR[ 123 ][ 90 ],
   alphaCSR[ 123 ][ 91 ],
   alphaCSR[ 123 ][ 92 ],
   alphaCSR[ 123 ][ 93 ],
   alphaCSR[ 123 ][ 94 ],
   alphaCSR[ 123 ][ 95 ],
   alphaCSR[ 123 ][ 96 ],
   alphaCSR[ 123 ][ 97 ],
   alphaCSR[ 123 ][ 98 ],
   alphaCSR[ 123 ][ 99 ],
   alphaCSR[ 123 ][ 100 ],
   alphaCSR[ 123 ][ 101 ],
   alphaCSR[ 123 ][ 102 ],
   alphaCSR[ 123 ][ 103 ],
   alphaCSR[ 123 ][ 104 ],
   alphaCSR[ 123 ][ 105 ],
   alphaCSR[ 123 ][ 106 ],
   alphaCSR[ 123 ][ 107 ],
   alphaCSR[ 123 ][ 108 ],
   alphaCSR[ 123 ][ 109 ],
   alphaCSR[ 123 ][ 110 ],
   alphaCSR[ 123 ][ 111 ],
   alphaCSR[ 123 ][ 112 ],
   alphaCSR[ 123 ][ 113 ],
   alphaCSR[ 123 ][ 114 ],
   alphaCSR[ 123 ][ 115 ],
   alphaCSR[ 123 ][ 116 ],
   alphaCSR[ 123 ][ 117 ],
   alphaCSR[ 123 ][ 118 ],
   alphaCSR[ 123 ][ 119 ],
   alphaCSR[ 123 ][ 120 ],
   alphaCSR[ 123 ][ 121 ],
   alphaCSR[ 123 ][ 122 ],
   alphaCSR[ 123 ][ 123 ],
   alphaCSR[ 123 ][ 124 ],
   alphaCSR[ 123 ][ 125 ],
   alphaCSR[ 123 ][ 126 ],
   alphaCSR[ 123 ][ 127 ],
   alphaCSR[ 123 ][ 128 ],
   alphaCSR[ 123 ][ 129 ],
   alphaCSR[ 123 ][ 130 ],
   alphaCSR[ 123 ][ 131 ],
   alphaCSR[ 123 ][ 132 ],
   alphaCSR[ 123 ][ 133 ],
   alphaCSR[ 123 ][ 134 ],
   alphaCSR[ 123 ][ 135 ],
   alphaCSR[ 123 ][ 136 ],
   alphaCSR[ 123 ][ 137 ],
   alphaCSR[ 123 ][ 138 ],
   alphaCSR[ 123 ][ 139 ],
   alphaCSR[ 123 ][ 140 ],
   alphaCSR[ 123 ][ 141 ],
   alphaCSR[ 123 ][ 142 ],
   alphaCSR[ 123 ][ 143 ],
   alphaCSR[ 123 ][ 144 ],
   alphaCSR[ 123 ][ 145 ],
   alphaCSR[ 123 ][ 146 ],
   alphaCSR[ 123 ][ 147 ],
   alphaCSR[ 123 ][ 148 ],
   alphaCSR[ 123 ][ 149 ],
   alphaCSR[ 123 ][ 150 ],
   alphaCSR[ 123 ][ 151 ],
   alphaCSR[ 123 ][ 152 ],
   alphaCSR[ 123 ][ 153 ],
   alphaCSR[ 123 ][ 154 ],
   alphaCSR[ 123 ][ 155 ],
   alphaCSR[ 123 ][ 156 ],
   alphaCSR[ 123 ][ 157 ],
   alphaCSR[ 123 ][ 158 ],
   alphaCSR[ 123 ][ 159 ],
   alphaCSR[ 123 ][ 160 ],
   alphaCSR[ 123 ][ 161 ],
   alphaCSR[ 123 ][ 162 ],
   alphaCSR[ 123 ][ 163 ],
   alphaCSR[ 123 ][ 164 ],
   alphaCSR[ 123 ][ 165 ],
   alphaCSR[ 123 ][ 166 ],
   alphaCSR[ 123 ][ 167 ],
   alphaCSR[ 123 ][ 168 ],
   alphaCSR[ 123 ][ 169 ],
   alphaCSR[ 123 ][ 170 ],
   alphaCSR[ 123 ][ 171 ],
   alphaCSR[ 123 ][ 172 ],
   alphaCSR[ 123 ][ 173 ],
   alphaCSR[ 123 ][ 174 ],
   alphaCSR[ 123 ][ 175 ],
   alphaCSR[ 123 ][ 176 ],
   alphaCSR[ 123 ][ 177 ],
   alphaCSR[ 123 ][ 178 ],
   alphaCSR[ 123 ][ 179 ],
   alphaCSR[ 123 ][ 180 ],
   alphaCSR[ 123 ][ 181 ],
   alphaCSR[ 123 ][ 182 ],
   alphaCSR[ 123 ][ 183 ],
   alphaCSR[ 123 ][ 184 ],
   alphaCSR[ 123 ][ 185 ],
   alphaCSR[ 123 ][ 186 ],
   alphaCSR[ 123 ][ 187 ],
   alphaCSR[ 123 ][ 188 ],
   alphaCSR[ 123 ][ 189 ],
   alphaCSR[ 123 ][ 190 ],
   alphaCSR[ 123 ][ 191 ],
   alphaCSR[ 123 ][ 192 ],
   alphaCSR[ 123 ][ 193 ],
   alphaCSR[ 123 ][ 194 ],
   alphaCSR[ 123 ][ 195 ],
   alphaCSR[ 123 ][ 196 ],
   alphaCSR[ 123 ][ 197 ],
   alphaCSR[ 123 ][ 198 ],
   alphaCSR[ 123 ][ 199 ],
   alphaCSR[ 123 ][ 200 ],
   alphaCSR[ 123 ][ 201 ],
   alphaCSR[ 123 ][ 202 ],
   alphaCSR[ 123 ][ 203 ],
   alphaCSR[ 123 ][ 204 ],
   alphaCSR[ 123 ][ 205 ],
   alphaCSR[ 123 ][ 206 ],
   alphaCSR[ 123 ][ 207 ],
   alphaCSR[ 123 ][ 208 ],
   alphaCSR[ 123 ][ 209 ],
   alphaCSR[ 123 ][ 210 ],
   alphaCSR[ 123 ][ 211 ],
   alphaCSR[ 123 ][ 212 ],
   alphaCSR[ 123 ][ 213 ],
   alphaCSR[ 123 ][ 214 ],
   alphaCSR[ 123 ][ 215 ],
   alphaCSR[ 123 ][ 216 ],
   alphaCSR[ 123 ][ 217 ],
   alphaCSR[ 123 ][ 218 ],
   alphaCSR[ 123 ][ 219 ],
   alphaCSR[ 123 ][ 220 ],
   alphaCSR[ 123 ][ 221 ],
   alphaCSR[ 123 ][ 222 ],
   alphaCSR[ 123 ][ 223 ],
   alphaCSR[ 123 ][ 224 ],
   alphaCSR[ 123 ][ 225 ],
   alphaCSR[ 123 ][ 226 ],
   alphaCSR[ 123 ][ 227 ],
   alphaCSR[ 123 ][ 228 ],
   alphaCSR[ 123 ][ 229 ],
   alphaCSR[ 123 ][ 230 ],
   alphaCSR[ 123 ][ 231 ],
   alphaCSR[ 123 ][ 232 ],
   alphaCSR[ 123 ][ 233 ],
   alphaCSR[ 123 ][ 234 ],
   alphaCSR[ 123 ][ 235 ],
   alphaCSR[ 123 ][ 236 ],
   alphaCSR[ 123 ][ 237 ],
   alphaCSR[ 123 ][ 238 ],
   alphaCSR[ 123 ][ 239 ],
   alphaCSR[ 123 ][ 240 ],
   alphaCSR[ 123 ][ 241 ],
   alphaCSR[ 123 ][ 242 ],
   alphaCSR[ 123 ][ 243 ],
   alphaCSR[ 123 ][ 244 ],
   alphaCSR[ 123 ][ 245 ],
   alphaCSR[ 123 ][ 246 ],
   alphaCSR[ 123 ][ 247 ],
   alphaCSR[ 123 ][ 248 ],
   alphaCSR[ 123 ][ 249 ],
   alphaCSR[ 123 ][ 250 ],
   alphaCSR[ 123 ][ 251 ],
   alphaCSR[ 123 ][ 252 ],
   alphaCSR[ 123 ][ 253 ],
   alphaCSR[ 123 ][ 254 ],
   alphaCSR[ 123 ][ 255 ],
   alphaCSR[ 123 ][ 256 ],
   alphaCSR[ 123 ][ 257 ],
   alphaCSR[ 123 ][ 258 ],
   alphaCSR[ 123 ][ 259 ],
   alphaCSR[ 123 ][ 260 ],
   alphaCSR[ 123 ][ 261 ],
   alphaCSR[ 123 ][ 262 ],
   alphaCSR[ 123 ][ 263 ],
   alphaCSR[ 123 ][ 264 ],
   alphaCSR[ 123 ][ 265 ],
   alphaCSR[ 123 ][ 266 ],
   alphaCSR[ 123 ][ 267 ],
   alphaCSR[ 123 ][ 268 ],
   alphaCSR[ 123 ][ 269 ],
   alphaCSR[ 123 ][ 270 ],
   alphaCSR[ 123 ][ 271 ],
   alphaCSR[ 123 ][ 272 ],
   alphaCSR[ 123 ][ 273 ],
   alphaCSR[ 123 ][ 274 ],
   alphaCSR[ 123 ][ 275 ],
   alphaCSR[ 123 ][ 276 ],
   alphaCSR[ 123 ][ 277 ],
   alphaCSR[ 123 ][ 278 ],
   alphaCSR[ 123 ][ 279 ],
   alphaCSR[ 123 ][ 280 ],
   alphaCSR[ 123 ][ 281 ],
   alphaCSR[ 123 ][ 282 ],
   alphaCSR[ 123 ][ 283 ],
   alphaCSR[ 123 ][ 284 ],
   alphaCSR[ 123 ][ 285 ],
   alphaCSR[ 123 ][ 286 ],
   alphaCSR[ 123 ][ 287 ],
   alphaCSR[ 123 ][ 288 ],
   alphaCSR[ 123 ][ 289 ],
   alphaCSR[ 123 ][ 290 ],
   alphaCSR[ 123 ][ 291 ],
   alphaCSR[ 123 ][ 292 ],
   alphaCSR[ 123 ][ 293 ],
   alphaCSR[ 123 ][ 294 ],
   alphaCSR[ 123 ][ 295 ],
   alphaCSR[ 123 ][ 296 ],
   alphaCSR[ 123 ][ 297 ],
   alphaCSR[ 123 ][ 298 ],
   alphaCSR[ 123 ][ 299 ],
   alphaCSR[ 123 ][ 300 ],
   alphaCSR[ 123 ][ 301 ],
   alphaCSR[ 123 ][ 302 ],
   alphaCSR[ 123 ][ 303 ],
   alphaCSR[ 123 ][ 304 ],
   alphaCSR[ 123 ][ 305 ],
   alphaCSR[ 123 ][ 306 ],
   alphaCSR[ 123 ][ 307 ],
   alphaCSR[ 123 ][ 308 ],
   alphaCSR[ 123 ][ 309 ],
   alphaCSR[ 123 ][ 310 ],
   alphaCSR[ 123 ][ 311 ],
   alphaCSR[ 123 ][ 312 ],
   alphaCSR[ 123 ][ 313 ],
   alphaCSR[ 123 ][ 314 ],
   alphaCSR[ 123 ][ 315 ],
   alphaCSR[ 123 ][ 316 ],
   alphaCSR[ 123 ][ 317 ],
   alphaCSR[ 123 ][ 318 ],
   alphaCSR[ 123 ][ 319 ],
   alphaCSR[ 123 ][ 320 ],
   alphaCSR[ 123 ][ 321 ],
   alphaCSR[ 123 ][ 322 ],
   alphaCSR[ 123 ][ 323 ],
   alphaCSR[ 123 ][ 324 ],
   alphaCSR[ 123 ][ 325 ],
   alphaCSR[ 123 ][ 326 ],
   alphaCSR[ 123 ][ 327 ],
   alphaCSR[ 123 ][ 328 ],
   alphaCSR[ 123 ][ 329 ],
   alphaCSR[ 123 ][ 330 ],
   alphaCSR[ 123 ][ 331 ],
   alphaCSR[ 123 ][ 332 ],
   alphaCSR[ 123 ][ 333 ],
   alphaCSR[ 123 ][ 334 ],
   alphaCSR[ 123 ][ 335 ],
   alphaCSR[ 123 ][ 336 ],
   alphaCSR[ 123 ][ 337 ],
   alphaCSR[ 123 ][ 338 ],
   alphaCSR[ 123 ][ 339 ],
   alphaCSR[ 123 ][ 340 ],
   alphaCSR[ 123 ][ 341 ],
   alphaCSR[ 123 ][ 342 ],
   alphaCSR[ 123 ][ 343 ],
   alphaCSR[ 123 ][ 344 ],
   alphaCSR[ 123 ][ 345 ],
   alphaCSR[ 123 ][ 346 ],
   alphaCSR[ 123 ][ 347 ],
   alphaCSR[ 123 ][ 348 ],
   alphaCSR[ 123 ][ 349 ],
   alphaCSR[ 123 ][ 350 ],
   alphaCSR[ 123 ][ 351 ],
   alphaCSR[ 123 ][ 352 ],
   alphaCSR[ 123 ][ 353 ],
   alphaCSR[ 123 ][ 354 ],
   alphaCSR[ 123 ][ 355 ],
   alphaCSR[ 123 ][ 356 ],
   alphaCSR[ 123 ][ 357 ],
   alphaCSR[ 123 ][ 358 ],
   alphaCSR[ 123 ][ 359 ],
   alphaCSR[ 123 ][ 360 ],
   alphaCSR[ 123 ][ 361 ],
   alphaCSR[ 123 ][ 362 ],
   alphaCSR[ 123 ][ 363 ],
   alphaCSR[ 123 ][ 364 ],
   alphaCSR[ 123 ][ 365 ],
   alphaCSR[ 123 ][ 366 ],
   alphaCSR[ 123 ][ 367 ],
   alphaCSR[ 123 ][ 368 ],
   alphaCSR[ 123 ][ 369 ],
   alphaCSR[ 123 ][ 370 ],
   alphaCSR[ 123 ][ 371 ],
   alphaCSR[ 123 ][ 372 ],
   alphaCSR[ 123 ][ 373 ],
   alphaCSR[ 123 ][ 374 ],
   alphaCSR[ 123 ][ 375 ],
   alphaCSR[ 123 ][ 376 ],
   alphaCSR[ 123 ][ 377 ],
   alphaCSR[ 123 ][ 378 ],
   alphaCSR[ 123 ][ 379 ],
   alphaCSR[ 123 ][ 380 ],
   alphaCSR[ 123 ][ 381 ],
   alphaCSR[ 123 ][ 382 ],
   alphaCSR[ 123 ][ 383 ],
   alphaCSR[ 124 ][ 0 ],
   alphaCSR[ 124 ][ 1 ],
   alphaCSR[ 124 ][ 2 ],
   alphaCSR[ 124 ][ 3 ],
   alphaCSR[ 124 ][ 4 ],
   alphaCSR[ 124 ][ 5 ],
   alphaCSR[ 124 ][ 6 ],
   alphaCSR[ 124 ][ 7 ],
   alphaCSR[ 124 ][ 8 ],
   alphaCSR[ 124 ][ 9 ],
   alphaCSR[ 124 ][ 10 ],
   alphaCSR[ 124 ][ 11 ],
   alphaCSR[ 124 ][ 12 ],
   alphaCSR[ 124 ][ 13 ],
   alphaCSR[ 124 ][ 14 ],
   alphaCSR[ 124 ][ 15 ],
   alphaCSR[ 124 ][ 16 ],
   alphaCSR[ 124 ][ 17 ],
   alphaCSR[ 124 ][ 18 ],
   alphaCSR[ 124 ][ 19 ],
   alphaCSR[ 124 ][ 20 ],
   alphaCSR[ 124 ][ 21 ],
   alphaCSR[ 124 ][ 22 ],
   alphaCSR[ 124 ][ 23 ],
   alphaCSR[ 124 ][ 24 ],
   alphaCSR[ 124 ][ 25 ],
   alphaCSR[ 124 ][ 26 ],
   alphaCSR[ 124 ][ 27 ],
   alphaCSR[ 124 ][ 28 ],
   alphaCSR[ 124 ][ 29 ],
   alphaCSR[ 124 ][ 30 ],
   alphaCSR[ 124 ][ 31 ],
   alphaCSR[ 124 ][ 32 ],
   alphaCSR[ 124 ][ 33 ],
   alphaCSR[ 124 ][ 34 ],
   alphaCSR[ 124 ][ 35 ],
   alphaCSR[ 124 ][ 36 ],
   alphaCSR[ 124 ][ 37 ],
   alphaCSR[ 124 ][ 38 ],
   alphaCSR[ 124 ][ 39 ],
   alphaCSR[ 124 ][ 40 ],
   alphaCSR[ 124 ][ 41 ],
   alphaCSR[ 124 ][ 42 ],
   alphaCSR[ 124 ][ 43 ],
   alphaCSR[ 124 ][ 44 ],
   alphaCSR[ 124 ][ 45 ],
   alphaCSR[ 124 ][ 46 ],
   alphaCSR[ 124 ][ 47 ],
   alphaCSR[ 124 ][ 48 ],
   alphaCSR[ 124 ][ 49 ],
   alphaCSR[ 124 ][ 50 ],
   alphaCSR[ 124 ][ 51 ],
   alphaCSR[ 124 ][ 52 ],
   alphaCSR[ 124 ][ 53 ],
   alphaCSR[ 124 ][ 54 ],
   alphaCSR[ 124 ][ 55 ],
   alphaCSR[ 124 ][ 56 ],
   alphaCSR[ 124 ][ 57 ],
   alphaCSR[ 124 ][ 58 ],
   alphaCSR[ 124 ][ 59 ],
   alphaCSR[ 124 ][ 60 ],
   alphaCSR[ 124 ][ 61 ],
   alphaCSR[ 124 ][ 62 ],
   alphaCSR[ 124 ][ 63 ],
   alphaCSR[ 124 ][ 64 ],
   alphaCSR[ 124 ][ 65 ],
   alphaCSR[ 124 ][ 66 ],
   alphaCSR[ 124 ][ 67 ],
   alphaCSR[ 124 ][ 68 ],
   alphaCSR[ 124 ][ 69 ],
   alphaCSR[ 124 ][ 70 ],
   alphaCSR[ 124 ][ 71 ],
   alphaCSR[ 124 ][ 72 ],
   alphaCSR[ 124 ][ 73 ],
   alphaCSR[ 124 ][ 74 ],
   alphaCSR[ 124 ][ 75 ],
   alphaCSR[ 124 ][ 76 ],
   alphaCSR[ 124 ][ 77 ],
   alphaCSR[ 124 ][ 78 ],
   alphaCSR[ 124 ][ 79 ],
   alphaCSR[ 124 ][ 80 ],
   alphaCSR[ 124 ][ 81 ],
   alphaCSR[ 124 ][ 82 ],
   alphaCSR[ 124 ][ 83 ],
   alphaCSR[ 124 ][ 84 ],
   alphaCSR[ 124 ][ 85 ],
   alphaCSR[ 124 ][ 86 ],
   alphaCSR[ 124 ][ 87 ],
   alphaCSR[ 124 ][ 88 ],
   alphaCSR[ 124 ][ 89 ],
   alphaCSR[ 124 ][ 90 ],
   alphaCSR[ 124 ][ 91 ],
   alphaCSR[ 124 ][ 92 ],
   alphaCSR[ 124 ][ 93 ],
   alphaCSR[ 124 ][ 94 ],
   alphaCSR[ 124 ][ 95 ],
   alphaCSR[ 124 ][ 96 ],
   alphaCSR[ 124 ][ 97 ],
   alphaCSR[ 124 ][ 98 ],
   alphaCSR[ 124 ][ 99 ],
   alphaCSR[ 124 ][ 100 ],
   alphaCSR[ 124 ][ 101 ],
   alphaCSR[ 124 ][ 102 ],
   alphaCSR[ 124 ][ 103 ],
   alphaCSR[ 124 ][ 104 ],
   alphaCSR[ 124 ][ 105 ],
   alphaCSR[ 124 ][ 106 ],
   alphaCSR[ 124 ][ 107 ],
   alphaCSR[ 124 ][ 108 ],
   alphaCSR[ 124 ][ 109 ],
   alphaCSR[ 124 ][ 110 ],
   alphaCSR[ 124 ][ 111 ],
   alphaCSR[ 124 ][ 112 ],
   alphaCSR[ 124 ][ 113 ],
   alphaCSR[ 124 ][ 114 ],
   alphaCSR[ 124 ][ 115 ],
   alphaCSR[ 124 ][ 116 ],
   alphaCSR[ 124 ][ 117 ],
   alphaCSR[ 124 ][ 118 ],
   alphaCSR[ 124 ][ 119 ],
   alphaCSR[ 124 ][ 120 ],
   alphaCSR[ 124 ][ 121 ],
   alphaCSR[ 124 ][ 122 ],
   alphaCSR[ 124 ][ 123 ],
   alphaCSR[ 124 ][ 124 ],
   alphaCSR[ 124 ][ 125 ],
   alphaCSR[ 124 ][ 126 ],
   alphaCSR[ 124 ][ 127 ],
   alphaCSR[ 124 ][ 128 ],
   alphaCSR[ 124 ][ 129 ],
   alphaCSR[ 124 ][ 130 ],
   alphaCSR[ 124 ][ 131 ],
   alphaCSR[ 124 ][ 132 ],
   alphaCSR[ 124 ][ 133 ],
   alphaCSR[ 124 ][ 134 ],
   alphaCSR[ 124 ][ 135 ],
   alphaCSR[ 124 ][ 136 ],
   alphaCSR[ 124 ][ 137 ],
   alphaCSR[ 124 ][ 138 ],
   alphaCSR[ 124 ][ 139 ],
   alphaCSR[ 124 ][ 140 ],
   alphaCSR[ 124 ][ 141 ],
   alphaCSR[ 124 ][ 142 ],
   alphaCSR[ 124 ][ 143 ],
   alphaCSR[ 124 ][ 144 ],
   alphaCSR[ 124 ][ 145 ],
   alphaCSR[ 124 ][ 146 ],
   alphaCSR[ 124 ][ 147 ],
   alphaCSR[ 124 ][ 148 ],
   alphaCSR[ 124 ][ 149 ],
   alphaCSR[ 124 ][ 150 ],
   alphaCSR[ 124 ][ 151 ],
   alphaCSR[ 124 ][ 152 ],
   alphaCSR[ 124 ][ 153 ],
   alphaCSR[ 124 ][ 154 ],
   alphaCSR[ 124 ][ 155 ],
   alphaCSR[ 124 ][ 156 ],
   alphaCSR[ 124 ][ 157 ],
   alphaCSR[ 124 ][ 158 ],
   alphaCSR[ 124 ][ 159 ],
   alphaCSR[ 124 ][ 160 ],
   alphaCSR[ 124 ][ 161 ],
   alphaCSR[ 124 ][ 162 ],
   alphaCSR[ 124 ][ 163 ],
   alphaCSR[ 124 ][ 164 ],
   alphaCSR[ 124 ][ 165 ],
   alphaCSR[ 124 ][ 166 ],
   alphaCSR[ 124 ][ 167 ],
   alphaCSR[ 124 ][ 168 ],
   alphaCSR[ 124 ][ 169 ],
   alphaCSR[ 124 ][ 170 ],
   alphaCSR[ 124 ][ 171 ],
   alphaCSR[ 124 ][ 172 ],
   alphaCSR[ 124 ][ 173 ],
   alphaCSR[ 124 ][ 174 ],
   alphaCSR[ 124 ][ 175 ],
   alphaCSR[ 124 ][ 176 ],
   alphaCSR[ 124 ][ 177 ],
   alphaCSR[ 124 ][ 178 ],
   alphaCSR[ 124 ][ 179 ],
   alphaCSR[ 124 ][ 180 ],
   alphaCSR[ 124 ][ 181 ],
   alphaCSR[ 124 ][ 182 ],
   alphaCSR[ 124 ][ 183 ],
   alphaCSR[ 124 ][ 184 ],
   alphaCSR[ 124 ][ 185 ],
   alphaCSR[ 124 ][ 186 ],
   alphaCSR[ 124 ][ 187 ],
   alphaCSR[ 124 ][ 188 ],
   alphaCSR[ 124 ][ 189 ],
   alphaCSR[ 124 ][ 190 ],
   alphaCSR[ 124 ][ 191 ],
   alphaCSR[ 124 ][ 192 ],
   alphaCSR[ 124 ][ 193 ],
   alphaCSR[ 124 ][ 194 ],
   alphaCSR[ 124 ][ 195 ],
   alphaCSR[ 124 ][ 196 ],
   alphaCSR[ 124 ][ 197 ],
   alphaCSR[ 124 ][ 198 ],
   alphaCSR[ 124 ][ 199 ],
   alphaCSR[ 124 ][ 200 ],
   alphaCSR[ 124 ][ 201 ],
   alphaCSR[ 124 ][ 202 ],
   alphaCSR[ 124 ][ 203 ],
   alphaCSR[ 124 ][ 204 ],
   alphaCSR[ 124 ][ 205 ],
   alphaCSR[ 124 ][ 206 ],
   alphaCSR[ 124 ][ 207 ],
   alphaCSR[ 124 ][ 208 ],
   alphaCSR[ 124 ][ 209 ],
   alphaCSR[ 124 ][ 210 ],
   alphaCSR[ 124 ][ 211 ],
   alphaCSR[ 124 ][ 212 ],
   alphaCSR[ 124 ][ 213 ],
   alphaCSR[ 124 ][ 214 ],
   alphaCSR[ 124 ][ 215 ],
   alphaCSR[ 124 ][ 216 ],
   alphaCSR[ 124 ][ 217 ],
   alphaCSR[ 124 ][ 218 ],
   alphaCSR[ 124 ][ 219 ],
   alphaCSR[ 124 ][ 220 ],
   alphaCSR[ 124 ][ 221 ],
   alphaCSR[ 124 ][ 222 ],
   alphaCSR[ 124 ][ 223 ],
   alphaCSR[ 124 ][ 224 ],
   alphaCSR[ 124 ][ 225 ],
   alphaCSR[ 124 ][ 226 ],
   alphaCSR[ 124 ][ 227 ],
   alphaCSR[ 124 ][ 228 ],
   alphaCSR[ 124 ][ 229 ],
   alphaCSR[ 124 ][ 230 ],
   alphaCSR[ 124 ][ 231 ],
   alphaCSR[ 124 ][ 232 ],
   alphaCSR[ 124 ][ 233 ],
   alphaCSR[ 124 ][ 234 ],
   alphaCSR[ 124 ][ 235 ],
   alphaCSR[ 124 ][ 236 ],
   alphaCSR[ 124 ][ 237 ],
   alphaCSR[ 124 ][ 238 ],
   alphaCSR[ 124 ][ 239 ],
   alphaCSR[ 124 ][ 240 ],
   alphaCSR[ 124 ][ 241 ],
   alphaCSR[ 124 ][ 242 ],
   alphaCSR[ 124 ][ 243 ],
   alphaCSR[ 124 ][ 244 ],
   alphaCSR[ 124 ][ 245 ],
   alphaCSR[ 124 ][ 246 ],
   alphaCSR[ 124 ][ 247 ],
   alphaCSR[ 124 ][ 248 ],
   alphaCSR[ 124 ][ 249 ],
   alphaCSR[ 124 ][ 250 ],
   alphaCSR[ 124 ][ 251 ],
   alphaCSR[ 124 ][ 252 ],
   alphaCSR[ 124 ][ 253 ],
   alphaCSR[ 124 ][ 254 ],
   alphaCSR[ 124 ][ 255 ],
   alphaCSR[ 124 ][ 256 ],
   alphaCSR[ 124 ][ 257 ],
   alphaCSR[ 124 ][ 258 ],
   alphaCSR[ 124 ][ 259 ],
   alphaCSR[ 124 ][ 260 ],
   alphaCSR[ 124 ][ 261 ],
   alphaCSR[ 124 ][ 262 ],
   alphaCSR[ 124 ][ 263 ],
   alphaCSR[ 124 ][ 264 ],
   alphaCSR[ 124 ][ 265 ],
   alphaCSR[ 124 ][ 266 ],
   alphaCSR[ 124 ][ 267 ],
   alphaCSR[ 124 ][ 268 ],
   alphaCSR[ 124 ][ 269 ],
   alphaCSR[ 124 ][ 270 ],
   alphaCSR[ 124 ][ 271 ],
   alphaCSR[ 124 ][ 272 ],
   alphaCSR[ 124 ][ 273 ],
   alphaCSR[ 124 ][ 274 ],
   alphaCSR[ 124 ][ 275 ],
   alphaCSR[ 124 ][ 276 ],
   alphaCSR[ 124 ][ 277 ],
   alphaCSR[ 124 ][ 278 ],
   alphaCSR[ 124 ][ 279 ],
   alphaCSR[ 124 ][ 280 ],
   alphaCSR[ 124 ][ 281 ],
   alphaCSR[ 124 ][ 282 ],
   alphaCSR[ 124 ][ 283 ],
   alphaCSR[ 124 ][ 284 ],
   alphaCSR[ 124 ][ 285 ],
   alphaCSR[ 124 ][ 286 ],
   alphaCSR[ 124 ][ 287 ],
   alphaCSR[ 124 ][ 288 ],
   alphaCSR[ 124 ][ 289 ],
   alphaCSR[ 124 ][ 290 ],
   alphaCSR[ 124 ][ 291 ],
   alphaCSR[ 124 ][ 292 ],
   alphaCSR[ 124 ][ 293 ],
   alphaCSR[ 124 ][ 294 ],
   alphaCSR[ 124 ][ 295 ],
   alphaCSR[ 124 ][ 296 ],
   alphaCSR[ 124 ][ 297 ],
   alphaCSR[ 124 ][ 298 ],
   alphaCSR[ 124 ][ 299 ],
   alphaCSR[ 124 ][ 300 ],
   alphaCSR[ 124 ][ 301 ],
   alphaCSR[ 124 ][ 302 ],
   alphaCSR[ 124 ][ 303 ],
   alphaCSR[ 124 ][ 304 ],
   alphaCSR[ 124 ][ 305 ],
   alphaCSR[ 124 ][ 306 ],
   alphaCSR[ 124 ][ 307 ],
   alphaCSR[ 124 ][ 308 ],
   alphaCSR[ 124 ][ 309 ],
   alphaCSR[ 124 ][ 310 ],
   alphaCSR[ 124 ][ 311 ],
   alphaCSR[ 124 ][ 312 ],
   alphaCSR[ 124 ][ 313 ],
   alphaCSR[ 124 ][ 314 ],
   alphaCSR[ 124 ][ 315 ],
   alphaCSR[ 124 ][ 316 ],
   alphaCSR[ 124 ][ 317 ],
   alphaCSR[ 124 ][ 318 ],
   alphaCSR[ 124 ][ 319 ],
   alphaCSR[ 124 ][ 320 ],
   alphaCSR[ 124 ][ 321 ],
   alphaCSR[ 124 ][ 322 ],
   alphaCSR[ 124 ][ 323 ],
   alphaCSR[ 124 ][ 324 ],
   alphaCSR[ 124 ][ 325 ],
   alphaCSR[ 124 ][ 326 ],
   alphaCSR[ 124 ][ 327 ],
   alphaCSR[ 124 ][ 328 ],
   alphaCSR[ 124 ][ 329 ],
   alphaCSR[ 124 ][ 330 ],
   alphaCSR[ 124 ][ 331 ],
   alphaCSR[ 124 ][ 332 ],
   alphaCSR[ 124 ][ 333 ],
   alphaCSR[ 124 ][ 334 ],
   alphaCSR[ 124 ][ 335 ],
   alphaCSR[ 124 ][ 336 ],
   alphaCSR[ 124 ][ 337 ],
   alphaCSR[ 124 ][ 338 ],
   alphaCSR[ 124 ][ 339 ],
   alphaCSR[ 124 ][ 340 ],
   alphaCSR[ 124 ][ 341 ],
   alphaCSR[ 124 ][ 342 ],
   alphaCSR[ 124 ][ 343 ],
   alphaCSR[ 124 ][ 344 ],
   alphaCSR[ 124 ][ 345 ],
   alphaCSR[ 124 ][ 346 ],
   alphaCSR[ 124 ][ 347 ],
   alphaCSR[ 124 ][ 348 ],
   alphaCSR[ 124 ][ 349 ],
   alphaCSR[ 124 ][ 350 ],
   alphaCSR[ 124 ][ 351 ],
   alphaCSR[ 124 ][ 352 ],
   alphaCSR[ 124 ][ 353 ],
   alphaCSR[ 124 ][ 354 ],
   alphaCSR[ 124 ][ 355 ],
   alphaCSR[ 124 ][ 356 ],
   alphaCSR[ 124 ][ 357 ],
   alphaCSR[ 124 ][ 358 ],
   alphaCSR[ 124 ][ 359 ],
   alphaCSR[ 124 ][ 360 ],
   alphaCSR[ 124 ][ 361 ],
   alphaCSR[ 124 ][ 362 ],
   alphaCSR[ 124 ][ 363 ],
   alphaCSR[ 124 ][ 364 ],
   alphaCSR[ 124 ][ 365 ],
   alphaCSR[ 124 ][ 366 ],
   alphaCSR[ 124 ][ 367 ],
   alphaCSR[ 124 ][ 368 ],
   alphaCSR[ 124 ][ 369 ],
   alphaCSR[ 124 ][ 370 ],
   alphaCSR[ 124 ][ 371 ],
   alphaCSR[ 124 ][ 372 ],
   alphaCSR[ 124 ][ 373 ],
   alphaCSR[ 124 ][ 374 ],
   alphaCSR[ 124 ][ 375 ],
   alphaCSR[ 124 ][ 376 ],
   alphaCSR[ 124 ][ 377 ],
   alphaCSR[ 124 ][ 378 ],
   alphaCSR[ 124 ][ 379 ],
   alphaCSR[ 124 ][ 380 ],
   alphaCSR[ 124 ][ 381 ],
   alphaCSR[ 124 ][ 382 ],
   alphaCSR[ 124 ][ 383 ],
   alphaCSR[ 125 ][ 0 ],
   alphaCSR[ 125 ][ 1 ],
   alphaCSR[ 125 ][ 2 ],
   alphaCSR[ 125 ][ 3 ],
   alphaCSR[ 125 ][ 4 ],
   alphaCSR[ 125 ][ 5 ],
   alphaCSR[ 125 ][ 6 ],
   alphaCSR[ 125 ][ 7 ],
   alphaCSR[ 125 ][ 8 ],
   alphaCSR[ 125 ][ 9 ],
   alphaCSR[ 125 ][ 10 ],
   alphaCSR[ 125 ][ 11 ],
   alphaCSR[ 125 ][ 12 ],
   alphaCSR[ 125 ][ 13 ],
   alphaCSR[ 125 ][ 14 ],
   alphaCSR[ 125 ][ 15 ],
   alphaCSR[ 125 ][ 16 ],
   alphaCSR[ 125 ][ 17 ],
   alphaCSR[ 125 ][ 18 ],
   alphaCSR[ 125 ][ 19 ],
   alphaCSR[ 125 ][ 20 ],
   alphaCSR[ 125 ][ 21 ],
   alphaCSR[ 125 ][ 22 ],
   alphaCSR[ 125 ][ 23 ],
   alphaCSR[ 125 ][ 24 ],
   alphaCSR[ 125 ][ 25 ],
   alphaCSR[ 125 ][ 26 ],
   alphaCSR[ 125 ][ 27 ],
   alphaCSR[ 125 ][ 28 ],
   alphaCSR[ 125 ][ 29 ],
   alphaCSR[ 125 ][ 30 ],
   alphaCSR[ 125 ][ 31 ],
   alphaCSR[ 125 ][ 32 ],
   alphaCSR[ 125 ][ 33 ],
   alphaCSR[ 125 ][ 34 ],
   alphaCSR[ 125 ][ 35 ],
   alphaCSR[ 125 ][ 36 ],
   alphaCSR[ 125 ][ 37 ],
   alphaCSR[ 125 ][ 38 ],
   alphaCSR[ 125 ][ 39 ],
   alphaCSR[ 125 ][ 40 ],
   alphaCSR[ 125 ][ 41 ],
   alphaCSR[ 125 ][ 42 ],
   alphaCSR[ 125 ][ 43 ],
   alphaCSR[ 125 ][ 44 ],
   alphaCSR[ 125 ][ 45 ],
   alphaCSR[ 125 ][ 46 ],
   alphaCSR[ 125 ][ 47 ],
   alphaCSR[ 125 ][ 48 ],
   alphaCSR[ 125 ][ 49 ],
   alphaCSR[ 125 ][ 50 ],
   alphaCSR[ 125 ][ 51 ],
   alphaCSR[ 125 ][ 52 ],
   alphaCSR[ 125 ][ 53 ],
   alphaCSR[ 125 ][ 54 ],
   alphaCSR[ 125 ][ 55 ],
   alphaCSR[ 125 ][ 56 ],
   alphaCSR[ 125 ][ 57 ],
   alphaCSR[ 125 ][ 58 ],
   alphaCSR[ 125 ][ 59 ],
   alphaCSR[ 125 ][ 60 ],
   alphaCSR[ 125 ][ 61 ],
   alphaCSR[ 125 ][ 62 ],
   alphaCSR[ 125 ][ 63 ],
   alphaCSR[ 125 ][ 64 ],
   alphaCSR[ 125 ][ 65 ],
   alphaCSR[ 125 ][ 66 ],
   alphaCSR[ 125 ][ 67 ],
   alphaCSR[ 125 ][ 68 ],
   alphaCSR[ 125 ][ 69 ],
   alphaCSR[ 125 ][ 70 ],
   alphaCSR[ 125 ][ 71 ],
   alphaCSR[ 125 ][ 72 ],
   alphaCSR[ 125 ][ 73 ],
   alphaCSR[ 125 ][ 74 ],
   alphaCSR[ 125 ][ 75 ],
   alphaCSR[ 125 ][ 76 ],
   alphaCSR[ 125 ][ 77 ],
   alphaCSR[ 125 ][ 78 ],
   alphaCSR[ 125 ][ 79 ],
   alphaCSR[ 125 ][ 80 ],
   alphaCSR[ 125 ][ 81 ],
   alphaCSR[ 125 ][ 82 ],
   alphaCSR[ 125 ][ 83 ],
   alphaCSR[ 125 ][ 84 ],
   alphaCSR[ 125 ][ 85 ],
   alphaCSR[ 125 ][ 86 ],
   alphaCSR[ 125 ][ 87 ],
   alphaCSR[ 125 ][ 88 ],
   alphaCSR[ 125 ][ 89 ],
   alphaCSR[ 125 ][ 90 ],
   alphaCSR[ 125 ][ 91 ],
   alphaCSR[ 125 ][ 92 ],
   alphaCSR[ 125 ][ 93 ],
   alphaCSR[ 125 ][ 94 ],
   alphaCSR[ 125 ][ 95 ],
   alphaCSR[ 125 ][ 96 ],
   alphaCSR[ 125 ][ 97 ],
   alphaCSR[ 125 ][ 98 ],
   alphaCSR[ 125 ][ 99 ],
   alphaCSR[ 125 ][ 100 ],
   alphaCSR[ 125 ][ 101 ],
   alphaCSR[ 125 ][ 102 ],
   alphaCSR[ 125 ][ 103 ],
   alphaCSR[ 125 ][ 104 ],
   alphaCSR[ 125 ][ 105 ],
   alphaCSR[ 125 ][ 106 ],
   alphaCSR[ 125 ][ 107 ],
   alphaCSR[ 125 ][ 108 ],
   alphaCSR[ 125 ][ 109 ],
   alphaCSR[ 125 ][ 110 ],
   alphaCSR[ 125 ][ 111 ],
   alphaCSR[ 125 ][ 112 ],
   alphaCSR[ 125 ][ 113 ],
   alphaCSR[ 125 ][ 114 ],
   alphaCSR[ 125 ][ 115 ],
   alphaCSR[ 125 ][ 116 ],
   alphaCSR[ 125 ][ 117 ],
   alphaCSR[ 125 ][ 118 ],
   alphaCSR[ 125 ][ 119 ],
   alphaCSR[ 125 ][ 120 ],
   alphaCSR[ 125 ][ 121 ],
   alphaCSR[ 125 ][ 122 ],
   alphaCSR[ 125 ][ 123 ],
   alphaCSR[ 125 ][ 124 ],
   alphaCSR[ 125 ][ 125 ],
   alphaCSR[ 125 ][ 126 ],
   alphaCSR[ 125 ][ 127 ],
   alphaCSR[ 125 ][ 128 ],
   alphaCSR[ 125 ][ 129 ],
   alphaCSR[ 125 ][ 130 ],
   alphaCSR[ 125 ][ 131 ],
   alphaCSR[ 125 ][ 132 ],
   alphaCSR[ 125 ][ 133 ],
   alphaCSR[ 125 ][ 134 ],
   alphaCSR[ 125 ][ 135 ],
   alphaCSR[ 125 ][ 136 ],
   alphaCSR[ 125 ][ 137 ],
   alphaCSR[ 125 ][ 138 ],
   alphaCSR[ 125 ][ 139 ],
   alphaCSR[ 125 ][ 140 ],
   alphaCSR[ 125 ][ 141 ],
   alphaCSR[ 125 ][ 142 ],
   alphaCSR[ 125 ][ 143 ],
   alphaCSR[ 125 ][ 144 ],
   alphaCSR[ 125 ][ 145 ],
   alphaCSR[ 125 ][ 146 ],
   alphaCSR[ 125 ][ 147 ],
   alphaCSR[ 125 ][ 148 ],
   alphaCSR[ 125 ][ 149 ],
   alphaCSR[ 125 ][ 150 ],
   alphaCSR[ 125 ][ 151 ],
   alphaCSR[ 125 ][ 152 ],
   alphaCSR[ 125 ][ 153 ],
   alphaCSR[ 125 ][ 154 ],
   alphaCSR[ 125 ][ 155 ],
   alphaCSR[ 125 ][ 156 ],
   alphaCSR[ 125 ][ 157 ],
   alphaCSR[ 125 ][ 158 ],
   alphaCSR[ 125 ][ 159 ],
   alphaCSR[ 125 ][ 160 ],
   alphaCSR[ 125 ][ 161 ],
   alphaCSR[ 125 ][ 162 ],
   alphaCSR[ 125 ][ 163 ],
   alphaCSR[ 125 ][ 164 ],
   alphaCSR[ 125 ][ 165 ],
   alphaCSR[ 125 ][ 166 ],
   alphaCSR[ 125 ][ 167 ],
   alphaCSR[ 125 ][ 168 ],
   alphaCSR[ 125 ][ 169 ],
   alphaCSR[ 125 ][ 170 ],
   alphaCSR[ 125 ][ 171 ],
   alphaCSR[ 125 ][ 172 ],
   alphaCSR[ 125 ][ 173 ],
   alphaCSR[ 125 ][ 174 ],
   alphaCSR[ 125 ][ 175 ],
   alphaCSR[ 125 ][ 176 ],
   alphaCSR[ 125 ][ 177 ],
   alphaCSR[ 125 ][ 178 ],
   alphaCSR[ 125 ][ 179 ],
   alphaCSR[ 125 ][ 180 ],
   alphaCSR[ 125 ][ 181 ],
   alphaCSR[ 125 ][ 182 ],
   alphaCSR[ 125 ][ 183 ],
   alphaCSR[ 125 ][ 184 ],
   alphaCSR[ 125 ][ 185 ],
   alphaCSR[ 125 ][ 186 ],
   alphaCSR[ 125 ][ 187 ],
   alphaCSR[ 125 ][ 188 ],
   alphaCSR[ 125 ][ 189 ],
   alphaCSR[ 125 ][ 190 ],
   alphaCSR[ 125 ][ 191 ],
   alphaCSR[ 125 ][ 192 ],
   alphaCSR[ 125 ][ 193 ],
   alphaCSR[ 125 ][ 194 ],
   alphaCSR[ 125 ][ 195 ],
   alphaCSR[ 125 ][ 196 ],
   alphaCSR[ 125 ][ 197 ],
   alphaCSR[ 125 ][ 198 ],
   alphaCSR[ 125 ][ 199 ],
   alphaCSR[ 125 ][ 200 ],
   alphaCSR[ 125 ][ 201 ],
   alphaCSR[ 125 ][ 202 ],
   alphaCSR[ 125 ][ 203 ],
   alphaCSR[ 125 ][ 204 ],
   alphaCSR[ 125 ][ 205 ],
   alphaCSR[ 125 ][ 206 ],
   alphaCSR[ 125 ][ 207 ],
   alphaCSR[ 125 ][ 208 ],
   alphaCSR[ 125 ][ 209 ],
   alphaCSR[ 125 ][ 210 ],
   alphaCSR[ 125 ][ 211 ],
   alphaCSR[ 125 ][ 212 ],
   alphaCSR[ 125 ][ 213 ],
   alphaCSR[ 125 ][ 214 ],
   alphaCSR[ 125 ][ 215 ],
   alphaCSR[ 125 ][ 216 ],
   alphaCSR[ 125 ][ 217 ],
   alphaCSR[ 125 ][ 218 ],
   alphaCSR[ 125 ][ 219 ],
   alphaCSR[ 125 ][ 220 ],
   alphaCSR[ 125 ][ 221 ],
   alphaCSR[ 125 ][ 222 ],
   alphaCSR[ 125 ][ 223 ],
   alphaCSR[ 125 ][ 224 ],
   alphaCSR[ 125 ][ 225 ],
   alphaCSR[ 125 ][ 226 ],
   alphaCSR[ 125 ][ 227 ],
   alphaCSR[ 125 ][ 228 ],
   alphaCSR[ 125 ][ 229 ],
   alphaCSR[ 125 ][ 230 ],
   alphaCSR[ 125 ][ 231 ],
   alphaCSR[ 125 ][ 232 ],
   alphaCSR[ 125 ][ 233 ],
   alphaCSR[ 125 ][ 234 ],
   alphaCSR[ 125 ][ 235 ],
   alphaCSR[ 125 ][ 236 ],
   alphaCSR[ 125 ][ 237 ],
   alphaCSR[ 125 ][ 238 ],
   alphaCSR[ 125 ][ 239 ],
   alphaCSR[ 125 ][ 240 ],
   alphaCSR[ 125 ][ 241 ],
   alphaCSR[ 125 ][ 242 ],
   alphaCSR[ 125 ][ 243 ],
   alphaCSR[ 125 ][ 244 ],
   alphaCSR[ 125 ][ 245 ],
   alphaCSR[ 125 ][ 246 ],
   alphaCSR[ 125 ][ 247 ],
   alphaCSR[ 125 ][ 248 ],
   alphaCSR[ 125 ][ 249 ],
   alphaCSR[ 125 ][ 250 ],
   alphaCSR[ 125 ][ 251 ],
   alphaCSR[ 125 ][ 252 ],
   alphaCSR[ 125 ][ 253 ],
   alphaCSR[ 125 ][ 254 ],
   alphaCSR[ 125 ][ 255 ],
   alphaCSR[ 125 ][ 256 ],
   alphaCSR[ 125 ][ 257 ],
   alphaCSR[ 125 ][ 258 ],
   alphaCSR[ 125 ][ 259 ],
   alphaCSR[ 125 ][ 260 ],
   alphaCSR[ 125 ][ 261 ],
   alphaCSR[ 125 ][ 262 ],
   alphaCSR[ 125 ][ 263 ],
   alphaCSR[ 125 ][ 264 ],
   alphaCSR[ 125 ][ 265 ],
   alphaCSR[ 125 ][ 266 ],
   alphaCSR[ 125 ][ 267 ],
   alphaCSR[ 125 ][ 268 ],
   alphaCSR[ 125 ][ 269 ],
   alphaCSR[ 125 ][ 270 ],
   alphaCSR[ 125 ][ 271 ],
   alphaCSR[ 125 ][ 272 ],
   alphaCSR[ 125 ][ 273 ],
   alphaCSR[ 125 ][ 274 ],
   alphaCSR[ 125 ][ 275 ],
   alphaCSR[ 125 ][ 276 ],
   alphaCSR[ 125 ][ 277 ],
   alphaCSR[ 125 ][ 278 ],
   alphaCSR[ 125 ][ 279 ],
   alphaCSR[ 125 ][ 280 ],
   alphaCSR[ 125 ][ 281 ],
   alphaCSR[ 125 ][ 282 ],
   alphaCSR[ 125 ][ 283 ],
   alphaCSR[ 125 ][ 284 ],
   alphaCSR[ 125 ][ 285 ],
   alphaCSR[ 125 ][ 286 ],
   alphaCSR[ 125 ][ 287 ],
   alphaCSR[ 125 ][ 288 ],
   alphaCSR[ 125 ][ 289 ],
   alphaCSR[ 125 ][ 290 ],
   alphaCSR[ 125 ][ 291 ],
   alphaCSR[ 125 ][ 292 ],
   alphaCSR[ 125 ][ 293 ],
   alphaCSR[ 125 ][ 294 ],
   alphaCSR[ 125 ][ 295 ],
   alphaCSR[ 125 ][ 296 ],
   alphaCSR[ 125 ][ 297 ],
   alphaCSR[ 125 ][ 298 ],
   alphaCSR[ 125 ][ 299 ],
   alphaCSR[ 125 ][ 300 ],
   alphaCSR[ 125 ][ 301 ],
   alphaCSR[ 125 ][ 302 ],
   alphaCSR[ 125 ][ 303 ],
   alphaCSR[ 125 ][ 304 ],
   alphaCSR[ 125 ][ 305 ],
   alphaCSR[ 125 ][ 306 ],
   alphaCSR[ 125 ][ 307 ],
   alphaCSR[ 125 ][ 308 ],
   alphaCSR[ 125 ][ 309 ],
   alphaCSR[ 125 ][ 310 ],
   alphaCSR[ 125 ][ 311 ],
   alphaCSR[ 125 ][ 312 ],
   alphaCSR[ 125 ][ 313 ],
   alphaCSR[ 125 ][ 314 ],
   alphaCSR[ 125 ][ 315 ],
   alphaCSR[ 125 ][ 316 ],
   alphaCSR[ 125 ][ 317 ],
   alphaCSR[ 125 ][ 318 ],
   alphaCSR[ 125 ][ 319 ],
   alphaCSR[ 125 ][ 320 ],
   alphaCSR[ 125 ][ 321 ],
   alphaCSR[ 125 ][ 322 ],
   alphaCSR[ 125 ][ 323 ],
   alphaCSR[ 125 ][ 324 ],
   alphaCSR[ 125 ][ 325 ],
   alphaCSR[ 125 ][ 326 ],
   alphaCSR[ 125 ][ 327 ],
   alphaCSR[ 125 ][ 328 ],
   alphaCSR[ 125 ][ 329 ],
   alphaCSR[ 125 ][ 330 ],
   alphaCSR[ 125 ][ 331 ],
   alphaCSR[ 125 ][ 332 ],
   alphaCSR[ 125 ][ 333 ],
   alphaCSR[ 125 ][ 334 ],
   alphaCSR[ 125 ][ 335 ],
   alphaCSR[ 125 ][ 336 ],
   alphaCSR[ 125 ][ 337 ],
   alphaCSR[ 125 ][ 338 ],
   alphaCSR[ 125 ][ 339 ],
   alphaCSR[ 125 ][ 340 ],
   alphaCSR[ 125 ][ 341 ],
   alphaCSR[ 125 ][ 342 ],
   alphaCSR[ 125 ][ 343 ],
   alphaCSR[ 125 ][ 344 ],
   alphaCSR[ 125 ][ 345 ],
   alphaCSR[ 125 ][ 346 ],
   alphaCSR[ 125 ][ 347 ],
   alphaCSR[ 125 ][ 348 ],
   alphaCSR[ 125 ][ 349 ],
   alphaCSR[ 125 ][ 350 ],
   alphaCSR[ 125 ][ 351 ],
   alphaCSR[ 125 ][ 352 ],
   alphaCSR[ 125 ][ 353 ],
   alphaCSR[ 125 ][ 354 ],
   alphaCSR[ 125 ][ 355 ],
   alphaCSR[ 125 ][ 356 ],
   alphaCSR[ 125 ][ 357 ],
   alphaCSR[ 125 ][ 358 ],
   alphaCSR[ 125 ][ 359 ],
   alphaCSR[ 125 ][ 360 ],
   alphaCSR[ 125 ][ 361 ],
   alphaCSR[ 125 ][ 362 ],
   alphaCSR[ 125 ][ 363 ],
   alphaCSR[ 125 ][ 364 ],
   alphaCSR[ 125 ][ 365 ],
   alphaCSR[ 125 ][ 366 ],
   alphaCSR[ 125 ][ 367 ],
   alphaCSR[ 125 ][ 368 ],
   alphaCSR[ 125 ][ 369 ],
   alphaCSR[ 125 ][ 370 ],
   alphaCSR[ 125 ][ 371 ],
   alphaCSR[ 125 ][ 372 ],
   alphaCSR[ 125 ][ 373 ],
   alphaCSR[ 125 ][ 374 ],
   alphaCSR[ 125 ][ 375 ],
   alphaCSR[ 125 ][ 376 ],
   alphaCSR[ 125 ][ 377 ],
   alphaCSR[ 125 ][ 378 ],
   alphaCSR[ 125 ][ 379 ],
   alphaCSR[ 125 ][ 380 ],
   alphaCSR[ 125 ][ 381 ],
   alphaCSR[ 125 ][ 382 ],
   alphaCSR[ 125 ][ 383 ],
   alphaCSR[ 126 ][ 0 ],
   alphaCSR[ 126 ][ 1 ],
   alphaCSR[ 126 ][ 2 ],
   alphaCSR[ 126 ][ 3 ],
   alphaCSR[ 126 ][ 4 ],
   alphaCSR[ 126 ][ 5 ],
   alphaCSR[ 126 ][ 6 ],
   alphaCSR[ 126 ][ 7 ],
   alphaCSR[ 126 ][ 8 ],
   alphaCSR[ 126 ][ 9 ],
   alphaCSR[ 126 ][ 10 ],
   alphaCSR[ 126 ][ 11 ],
   alphaCSR[ 126 ][ 12 ],
   alphaCSR[ 126 ][ 13 ],
   alphaCSR[ 126 ][ 14 ],
   alphaCSR[ 126 ][ 15 ],
   alphaCSR[ 126 ][ 16 ],
   alphaCSR[ 126 ][ 17 ],
   alphaCSR[ 126 ][ 18 ],
   alphaCSR[ 126 ][ 19 ],
   alphaCSR[ 126 ][ 20 ],
   alphaCSR[ 126 ][ 21 ],
   alphaCSR[ 126 ][ 22 ],
   alphaCSR[ 126 ][ 23 ],
   alphaCSR[ 126 ][ 24 ],
   alphaCSR[ 126 ][ 25 ],
   alphaCSR[ 126 ][ 26 ],
   alphaCSR[ 126 ][ 27 ],
   alphaCSR[ 126 ][ 28 ],
   alphaCSR[ 126 ][ 29 ],
   alphaCSR[ 126 ][ 30 ],
   alphaCSR[ 126 ][ 31 ],
   alphaCSR[ 126 ][ 32 ],
   alphaCSR[ 126 ][ 33 ],
   alphaCSR[ 126 ][ 34 ],
   alphaCSR[ 126 ][ 35 ],
   alphaCSR[ 126 ][ 36 ],
   alphaCSR[ 126 ][ 37 ],
   alphaCSR[ 126 ][ 38 ],
   alphaCSR[ 126 ][ 39 ],
   alphaCSR[ 126 ][ 40 ],
   alphaCSR[ 126 ][ 41 ],
   alphaCSR[ 126 ][ 42 ],
   alphaCSR[ 126 ][ 43 ],
   alphaCSR[ 126 ][ 44 ],
   alphaCSR[ 126 ][ 45 ],
   alphaCSR[ 126 ][ 46 ],
   alphaCSR[ 126 ][ 47 ],
   alphaCSR[ 126 ][ 48 ],
   alphaCSR[ 126 ][ 49 ],
   alphaCSR[ 126 ][ 50 ],
   alphaCSR[ 126 ][ 51 ],
   alphaCSR[ 126 ][ 52 ],
   alphaCSR[ 126 ][ 53 ],
   alphaCSR[ 126 ][ 54 ],
   alphaCSR[ 126 ][ 55 ],
   alphaCSR[ 126 ][ 56 ],
   alphaCSR[ 126 ][ 57 ],
   alphaCSR[ 126 ][ 58 ],
   alphaCSR[ 126 ][ 59 ],
   alphaCSR[ 126 ][ 60 ],
   alphaCSR[ 126 ][ 61 ],
   alphaCSR[ 126 ][ 62 ],
   alphaCSR[ 126 ][ 63 ],
   alphaCSR[ 126 ][ 64 ],
   alphaCSR[ 126 ][ 65 ],
   alphaCSR[ 126 ][ 66 ],
   alphaCSR[ 126 ][ 67 ],
   alphaCSR[ 126 ][ 68 ],
   alphaCSR[ 126 ][ 69 ],
   alphaCSR[ 126 ][ 70 ],
   alphaCSR[ 126 ][ 71 ],
   alphaCSR[ 126 ][ 72 ],
   alphaCSR[ 126 ][ 73 ],
   alphaCSR[ 126 ][ 74 ],
   alphaCSR[ 126 ][ 75 ],
   alphaCSR[ 126 ][ 76 ],
   alphaCSR[ 126 ][ 77 ],
   alphaCSR[ 126 ][ 78 ],
   alphaCSR[ 126 ][ 79 ],
   alphaCSR[ 126 ][ 80 ],
   alphaCSR[ 126 ][ 81 ],
   alphaCSR[ 126 ][ 82 ],
   alphaCSR[ 126 ][ 83 ],
   alphaCSR[ 126 ][ 84 ],
   alphaCSR[ 126 ][ 85 ],
   alphaCSR[ 126 ][ 86 ],
   alphaCSR[ 126 ][ 87 ],
   alphaCSR[ 126 ][ 88 ],
   alphaCSR[ 126 ][ 89 ],
   alphaCSR[ 126 ][ 90 ],
   alphaCSR[ 126 ][ 91 ],
   alphaCSR[ 126 ][ 92 ],
   alphaCSR[ 126 ][ 93 ],
   alphaCSR[ 126 ][ 94 ],
   alphaCSR[ 126 ][ 95 ],
   alphaCSR[ 126 ][ 96 ],
   alphaCSR[ 126 ][ 97 ],
   alphaCSR[ 126 ][ 98 ],
   alphaCSR[ 126 ][ 99 ],
   alphaCSR[ 126 ][ 100 ],
   alphaCSR[ 126 ][ 101 ],
   alphaCSR[ 126 ][ 102 ],
   alphaCSR[ 126 ][ 103 ],
   alphaCSR[ 126 ][ 104 ],
   alphaCSR[ 126 ][ 105 ],
   alphaCSR[ 126 ][ 106 ],
   alphaCSR[ 126 ][ 107 ],
   alphaCSR[ 126 ][ 108 ],
   alphaCSR[ 126 ][ 109 ],
   alphaCSR[ 126 ][ 110 ],
   alphaCSR[ 126 ][ 111 ],
   alphaCSR[ 126 ][ 112 ],
   alphaCSR[ 126 ][ 113 ],
   alphaCSR[ 126 ][ 114 ],
   alphaCSR[ 126 ][ 115 ],
   alphaCSR[ 126 ][ 116 ],
   alphaCSR[ 126 ][ 117 ],
   alphaCSR[ 126 ][ 118 ],
   alphaCSR[ 126 ][ 119 ],
   alphaCSR[ 126 ][ 120 ],
   alphaCSR[ 126 ][ 121 ],
   alphaCSR[ 126 ][ 122 ],
   alphaCSR[ 126 ][ 123 ],
   alphaCSR[ 126 ][ 124 ],
   alphaCSR[ 126 ][ 125 ],
   alphaCSR[ 126 ][ 126 ],
   alphaCSR[ 126 ][ 127 ],
   alphaCSR[ 126 ][ 128 ],
   alphaCSR[ 126 ][ 129 ],
   alphaCSR[ 126 ][ 130 ],
   alphaCSR[ 126 ][ 131 ],
   alphaCSR[ 126 ][ 132 ],
   alphaCSR[ 126 ][ 133 ],
   alphaCSR[ 126 ][ 134 ],
   alphaCSR[ 126 ][ 135 ],
   alphaCSR[ 126 ][ 136 ],
   alphaCSR[ 126 ][ 137 ],
   alphaCSR[ 126 ][ 138 ],
   alphaCSR[ 126 ][ 139 ],
   alphaCSR[ 126 ][ 140 ],
   alphaCSR[ 126 ][ 141 ],
   alphaCSR[ 126 ][ 142 ],
   alphaCSR[ 126 ][ 143 ],
   alphaCSR[ 126 ][ 144 ],
   alphaCSR[ 126 ][ 145 ],
   alphaCSR[ 126 ][ 146 ],
   alphaCSR[ 126 ][ 147 ],
   alphaCSR[ 126 ][ 148 ],
   alphaCSR[ 126 ][ 149 ],
   alphaCSR[ 126 ][ 150 ],
   alphaCSR[ 126 ][ 151 ],
   alphaCSR[ 126 ][ 152 ],
   alphaCSR[ 126 ][ 153 ],
   alphaCSR[ 126 ][ 154 ],
   alphaCSR[ 126 ][ 155 ],
   alphaCSR[ 126 ][ 156 ],
   alphaCSR[ 126 ][ 157 ],
   alphaCSR[ 126 ][ 158 ],
   alphaCSR[ 126 ][ 159 ],
   alphaCSR[ 126 ][ 160 ],
   alphaCSR[ 126 ][ 161 ],
   alphaCSR[ 126 ][ 162 ],
   alphaCSR[ 126 ][ 163 ],
   alphaCSR[ 126 ][ 164 ],
   alphaCSR[ 126 ][ 165 ],
   alphaCSR[ 126 ][ 166 ],
   alphaCSR[ 126 ][ 167 ],
   alphaCSR[ 126 ][ 168 ],
   alphaCSR[ 126 ][ 169 ],
   alphaCSR[ 126 ][ 170 ],
   alphaCSR[ 126 ][ 171 ],
   alphaCSR[ 126 ][ 172 ],
   alphaCSR[ 126 ][ 173 ],
   alphaCSR[ 126 ][ 174 ],
   alphaCSR[ 126 ][ 175 ],
   alphaCSR[ 126 ][ 176 ],
   alphaCSR[ 126 ][ 177 ],
   alphaCSR[ 126 ][ 178 ],
   alphaCSR[ 126 ][ 179 ],
   alphaCSR[ 126 ][ 180 ],
   alphaCSR[ 126 ][ 181 ],
   alphaCSR[ 126 ][ 182 ],
   alphaCSR[ 126 ][ 183 ],
   alphaCSR[ 126 ][ 184 ],
   alphaCSR[ 126 ][ 185 ],
   alphaCSR[ 126 ][ 186 ],
   alphaCSR[ 126 ][ 187 ],
   alphaCSR[ 126 ][ 188 ],
   alphaCSR[ 126 ][ 189 ],
   alphaCSR[ 126 ][ 190 ],
   alphaCSR[ 126 ][ 191 ],
   alphaCSR[ 126 ][ 192 ],
   alphaCSR[ 126 ][ 193 ],
   alphaCSR[ 126 ][ 194 ],
   alphaCSR[ 126 ][ 195 ],
   alphaCSR[ 126 ][ 196 ],
   alphaCSR[ 126 ][ 197 ],
   alphaCSR[ 126 ][ 198 ],
   alphaCSR[ 126 ][ 199 ],
   alphaCSR[ 126 ][ 200 ],
   alphaCSR[ 126 ][ 201 ],
   alphaCSR[ 126 ][ 202 ],
   alphaCSR[ 126 ][ 203 ],
   alphaCSR[ 126 ][ 204 ],
   alphaCSR[ 126 ][ 205 ],
   alphaCSR[ 126 ][ 206 ],
   alphaCSR[ 126 ][ 207 ],
   alphaCSR[ 126 ][ 208 ],
   alphaCSR[ 126 ][ 209 ],
   alphaCSR[ 126 ][ 210 ],
   alphaCSR[ 126 ][ 211 ],
   alphaCSR[ 126 ][ 212 ],
   alphaCSR[ 126 ][ 213 ],
   alphaCSR[ 126 ][ 214 ],
   alphaCSR[ 126 ][ 215 ],
   alphaCSR[ 126 ][ 216 ],
   alphaCSR[ 126 ][ 217 ],
   alphaCSR[ 126 ][ 218 ],
   alphaCSR[ 126 ][ 219 ],
   alphaCSR[ 126 ][ 220 ],
   alphaCSR[ 126 ][ 221 ],
   alphaCSR[ 126 ][ 222 ],
   alphaCSR[ 126 ][ 223 ],
   alphaCSR[ 126 ][ 224 ],
   alphaCSR[ 126 ][ 225 ],
   alphaCSR[ 126 ][ 226 ],
   alphaCSR[ 126 ][ 227 ],
   alphaCSR[ 126 ][ 228 ],
   alphaCSR[ 126 ][ 229 ],
   alphaCSR[ 126 ][ 230 ],
   alphaCSR[ 126 ][ 231 ],
   alphaCSR[ 126 ][ 232 ],
   alphaCSR[ 126 ][ 233 ],
   alphaCSR[ 126 ][ 234 ],
   alphaCSR[ 126 ][ 235 ],
   alphaCSR[ 126 ][ 236 ],
   alphaCSR[ 126 ][ 237 ],
   alphaCSR[ 126 ][ 238 ],
   alphaCSR[ 126 ][ 239 ],
   alphaCSR[ 126 ][ 240 ],
   alphaCSR[ 126 ][ 241 ],
   alphaCSR[ 126 ][ 242 ],
   alphaCSR[ 126 ][ 243 ],
   alphaCSR[ 126 ][ 244 ],
   alphaCSR[ 126 ][ 245 ],
   alphaCSR[ 126 ][ 246 ],
   alphaCSR[ 126 ][ 247 ],
   alphaCSR[ 126 ][ 248 ],
   alphaCSR[ 126 ][ 249 ],
   alphaCSR[ 126 ][ 250 ],
   alphaCSR[ 126 ][ 251 ],
   alphaCSR[ 126 ][ 252 ],
   alphaCSR[ 126 ][ 253 ],
   alphaCSR[ 126 ][ 254 ],
   alphaCSR[ 126 ][ 255 ],
   alphaCSR[ 126 ][ 256 ],
   alphaCSR[ 126 ][ 257 ],
   alphaCSR[ 126 ][ 258 ],
   alphaCSR[ 126 ][ 259 ],
   alphaCSR[ 126 ][ 260 ],
   alphaCSR[ 126 ][ 261 ],
   alphaCSR[ 126 ][ 262 ],
   alphaCSR[ 126 ][ 263 ],
   alphaCSR[ 126 ][ 264 ],
   alphaCSR[ 126 ][ 265 ],
   alphaCSR[ 126 ][ 266 ],
   alphaCSR[ 126 ][ 267 ],
   alphaCSR[ 126 ][ 268 ],
   alphaCSR[ 126 ][ 269 ],
   alphaCSR[ 126 ][ 270 ],
   alphaCSR[ 126 ][ 271 ],
   alphaCSR[ 126 ][ 272 ],
   alphaCSR[ 126 ][ 273 ],
   alphaCSR[ 126 ][ 274 ],
   alphaCSR[ 126 ][ 275 ],
   alphaCSR[ 126 ][ 276 ],
   alphaCSR[ 126 ][ 277 ],
   alphaCSR[ 126 ][ 278 ],
   alphaCSR[ 126 ][ 279 ],
   alphaCSR[ 126 ][ 280 ],
   alphaCSR[ 126 ][ 281 ],
   alphaCSR[ 126 ][ 282 ],
   alphaCSR[ 126 ][ 283 ],
   alphaCSR[ 126 ][ 284 ],
   alphaCSR[ 126 ][ 285 ],
   alphaCSR[ 126 ][ 286 ],
   alphaCSR[ 126 ][ 287 ],
   alphaCSR[ 126 ][ 288 ],
   alphaCSR[ 126 ][ 289 ],
   alphaCSR[ 126 ][ 290 ],
   alphaCSR[ 126 ][ 291 ],
   alphaCSR[ 126 ][ 292 ],
   alphaCSR[ 126 ][ 293 ],
   alphaCSR[ 126 ][ 294 ],
   alphaCSR[ 126 ][ 295 ],
   alphaCSR[ 126 ][ 296 ],
   alphaCSR[ 126 ][ 297 ],
   alphaCSR[ 126 ][ 298 ],
   alphaCSR[ 126 ][ 299 ],
   alphaCSR[ 126 ][ 300 ],
   alphaCSR[ 126 ][ 301 ],
   alphaCSR[ 126 ][ 302 ],
   alphaCSR[ 126 ][ 303 ],
   alphaCSR[ 126 ][ 304 ],
   alphaCSR[ 126 ][ 305 ],
   alphaCSR[ 126 ][ 306 ],
   alphaCSR[ 126 ][ 307 ],
   alphaCSR[ 126 ][ 308 ],
   alphaCSR[ 126 ][ 309 ],
   alphaCSR[ 126 ][ 310 ],
   alphaCSR[ 126 ][ 311 ],
   alphaCSR[ 126 ][ 312 ],
   alphaCSR[ 126 ][ 313 ],
   alphaCSR[ 126 ][ 314 ],
   alphaCSR[ 126 ][ 315 ],
   alphaCSR[ 126 ][ 316 ],
   alphaCSR[ 126 ][ 317 ],
   alphaCSR[ 126 ][ 318 ],
   alphaCSR[ 126 ][ 319 ],
   alphaCSR[ 126 ][ 320 ],
   alphaCSR[ 126 ][ 321 ],
   alphaCSR[ 126 ][ 322 ],
   alphaCSR[ 126 ][ 323 ],
   alphaCSR[ 126 ][ 324 ],
   alphaCSR[ 126 ][ 325 ],
   alphaCSR[ 126 ][ 326 ],
   alphaCSR[ 126 ][ 327 ],
   alphaCSR[ 126 ][ 328 ],
   alphaCSR[ 126 ][ 329 ],
   alphaCSR[ 126 ][ 330 ],
   alphaCSR[ 126 ][ 331 ],
   alphaCSR[ 126 ][ 332 ],
   alphaCSR[ 126 ][ 333 ],
   alphaCSR[ 126 ][ 334 ],
   alphaCSR[ 126 ][ 335 ],
   alphaCSR[ 126 ][ 336 ],
   alphaCSR[ 126 ][ 337 ],
   alphaCSR[ 126 ][ 338 ],
   alphaCSR[ 126 ][ 339 ],
   alphaCSR[ 126 ][ 340 ],
   alphaCSR[ 126 ][ 341 ],
   alphaCSR[ 126 ][ 342 ],
   alphaCSR[ 126 ][ 343 ],
   alphaCSR[ 126 ][ 344 ],
   alphaCSR[ 126 ][ 345 ],
   alphaCSR[ 126 ][ 346 ],
   alphaCSR[ 126 ][ 347 ],
   alphaCSR[ 126 ][ 348 ],
   alphaCSR[ 126 ][ 349 ],
   alphaCSR[ 126 ][ 350 ],
   alphaCSR[ 126 ][ 351 ],
   alphaCSR[ 126 ][ 352 ],
   alphaCSR[ 126 ][ 353 ],
   alphaCSR[ 126 ][ 354 ],
   alphaCSR[ 126 ][ 355 ],
   alphaCSR[ 126 ][ 356 ],
   alphaCSR[ 126 ][ 357 ],
   alphaCSR[ 126 ][ 358 ],
   alphaCSR[ 126 ][ 359 ],
   alphaCSR[ 126 ][ 360 ],
   alphaCSR[ 126 ][ 361 ],
   alphaCSR[ 126 ][ 362 ],
   alphaCSR[ 126 ][ 363 ],
   alphaCSR[ 126 ][ 364 ],
   alphaCSR[ 126 ][ 365 ],
   alphaCSR[ 126 ][ 366 ],
   alphaCSR[ 126 ][ 367 ],
   alphaCSR[ 126 ][ 368 ],
   alphaCSR[ 126 ][ 369 ],
   alphaCSR[ 126 ][ 370 ],
   alphaCSR[ 126 ][ 371 ],
   alphaCSR[ 126 ][ 372 ],
   alphaCSR[ 126 ][ 373 ],
   alphaCSR[ 126 ][ 374 ],
   alphaCSR[ 126 ][ 375 ],
   alphaCSR[ 126 ][ 376 ],
   alphaCSR[ 126 ][ 377 ],
   alphaCSR[ 126 ][ 378 ],
   alphaCSR[ 126 ][ 379 ],
   alphaCSR[ 126 ][ 380 ],
   alphaCSR[ 126 ][ 381 ],
   alphaCSR[ 126 ][ 382 ],
   alphaCSR[ 126 ][ 383 ],
   alphaCSR[ 127 ][ 0 ],
   alphaCSR[ 127 ][ 1 ],
   alphaCSR[ 127 ][ 2 ],
   alphaCSR[ 127 ][ 3 ],
   alphaCSR[ 127 ][ 4 ],
   alphaCSR[ 127 ][ 5 ],
   alphaCSR[ 127 ][ 6 ],
   alphaCSR[ 127 ][ 7 ],
   alphaCSR[ 127 ][ 8 ],
   alphaCSR[ 127 ][ 9 ],
   alphaCSR[ 127 ][ 10 ],
   alphaCSR[ 127 ][ 11 ],
   alphaCSR[ 127 ][ 12 ],
   alphaCSR[ 127 ][ 13 ],
   alphaCSR[ 127 ][ 14 ],
   alphaCSR[ 127 ][ 15 ],
   alphaCSR[ 127 ][ 16 ],
   alphaCSR[ 127 ][ 17 ],
   alphaCSR[ 127 ][ 18 ],
   alphaCSR[ 127 ][ 19 ],
   alphaCSR[ 127 ][ 20 ],
   alphaCSR[ 127 ][ 21 ],
   alphaCSR[ 127 ][ 22 ],
   alphaCSR[ 127 ][ 23 ],
   alphaCSR[ 127 ][ 24 ],
   alphaCSR[ 127 ][ 25 ],
   alphaCSR[ 127 ][ 26 ],
   alphaCSR[ 127 ][ 27 ],
   alphaCSR[ 127 ][ 28 ],
   alphaCSR[ 127 ][ 29 ],
   alphaCSR[ 127 ][ 30 ],
   alphaCSR[ 127 ][ 31 ],
   alphaCSR[ 127 ][ 32 ],
   alphaCSR[ 127 ][ 33 ],
   alphaCSR[ 127 ][ 34 ],
   alphaCSR[ 127 ][ 35 ],
   alphaCSR[ 127 ][ 36 ],
   alphaCSR[ 127 ][ 37 ],
   alphaCSR[ 127 ][ 38 ],
   alphaCSR[ 127 ][ 39 ],
   alphaCSR[ 127 ][ 40 ],
   alphaCSR[ 127 ][ 41 ],
   alphaCSR[ 127 ][ 42 ],
   alphaCSR[ 127 ][ 43 ],
   alphaCSR[ 127 ][ 44 ],
   alphaCSR[ 127 ][ 45 ],
   alphaCSR[ 127 ][ 46 ],
   alphaCSR[ 127 ][ 47 ],
   alphaCSR[ 127 ][ 48 ],
   alphaCSR[ 127 ][ 49 ],
   alphaCSR[ 127 ][ 50 ],
   alphaCSR[ 127 ][ 51 ],
   alphaCSR[ 127 ][ 52 ],
   alphaCSR[ 127 ][ 53 ],
   alphaCSR[ 127 ][ 54 ],
   alphaCSR[ 127 ][ 55 ],
   alphaCSR[ 127 ][ 56 ],
   alphaCSR[ 127 ][ 57 ],
   alphaCSR[ 127 ][ 58 ],
   alphaCSR[ 127 ][ 59 ],
   alphaCSR[ 127 ][ 60 ],
   alphaCSR[ 127 ][ 61 ],
   alphaCSR[ 127 ][ 62 ],
   alphaCSR[ 127 ][ 63 ],
   alphaCSR[ 127 ][ 64 ],
   alphaCSR[ 127 ][ 65 ],
   alphaCSR[ 127 ][ 66 ],
   alphaCSR[ 127 ][ 67 ],
   alphaCSR[ 127 ][ 68 ],
   alphaCSR[ 127 ][ 69 ],
   alphaCSR[ 127 ][ 70 ],
   alphaCSR[ 127 ][ 71 ],
   alphaCSR[ 127 ][ 72 ],
   alphaCSR[ 127 ][ 73 ],
   alphaCSR[ 127 ][ 74 ],
   alphaCSR[ 127 ][ 75 ],
   alphaCSR[ 127 ][ 76 ],
   alphaCSR[ 127 ][ 77 ],
   alphaCSR[ 127 ][ 78 ],
   alphaCSR[ 127 ][ 79 ],
   alphaCSR[ 127 ][ 80 ],
   alphaCSR[ 127 ][ 81 ],
   alphaCSR[ 127 ][ 82 ],
   alphaCSR[ 127 ][ 83 ],
   alphaCSR[ 127 ][ 84 ],
   alphaCSR[ 127 ][ 85 ],
   alphaCSR[ 127 ][ 86 ],
   alphaCSR[ 127 ][ 87 ],
   alphaCSR[ 127 ][ 88 ],
   alphaCSR[ 127 ][ 89 ],
   alphaCSR[ 127 ][ 90 ],
   alphaCSR[ 127 ][ 91 ],
   alphaCSR[ 127 ][ 92 ],
   alphaCSR[ 127 ][ 93 ],
   alphaCSR[ 127 ][ 94 ],
   alphaCSR[ 127 ][ 95 ],
   alphaCSR[ 127 ][ 96 ],
   alphaCSR[ 127 ][ 97 ],
   alphaCSR[ 127 ][ 98 ],
   alphaCSR[ 127 ][ 99 ],
   alphaCSR[ 127 ][ 100 ],
   alphaCSR[ 127 ][ 101 ],
   alphaCSR[ 127 ][ 102 ],
   alphaCSR[ 127 ][ 103 ],
   alphaCSR[ 127 ][ 104 ],
   alphaCSR[ 127 ][ 105 ],
   alphaCSR[ 127 ][ 106 ],
   alphaCSR[ 127 ][ 107 ],
   alphaCSR[ 127 ][ 108 ],
   alphaCSR[ 127 ][ 109 ],
   alphaCSR[ 127 ][ 110 ],
   alphaCSR[ 127 ][ 111 ],
   alphaCSR[ 127 ][ 112 ],
   alphaCSR[ 127 ][ 113 ],
   alphaCSR[ 127 ][ 114 ],
   alphaCSR[ 127 ][ 115 ],
   alphaCSR[ 127 ][ 116 ],
   alphaCSR[ 127 ][ 117 ],
   alphaCSR[ 127 ][ 118 ],
   alphaCSR[ 127 ][ 119 ],
   alphaCSR[ 127 ][ 120 ],
   alphaCSR[ 127 ][ 121 ],
   alphaCSR[ 127 ][ 122 ],
   alphaCSR[ 127 ][ 123 ],
   alphaCSR[ 127 ][ 124 ],
   alphaCSR[ 127 ][ 125 ],
   alphaCSR[ 127 ][ 126 ],
   alphaCSR[ 127 ][ 127 ],
   alphaCSR[ 127 ][ 128 ],
   alphaCSR[ 127 ][ 129 ],
   alphaCSR[ 127 ][ 130 ],
   alphaCSR[ 127 ][ 131 ],
   alphaCSR[ 127 ][ 132 ],
   alphaCSR[ 127 ][ 133 ],
   alphaCSR[ 127 ][ 134 ],
   alphaCSR[ 127 ][ 135 ],
   alphaCSR[ 127 ][ 136 ],
   alphaCSR[ 127 ][ 137 ],
   alphaCSR[ 127 ][ 138 ],
   alphaCSR[ 127 ][ 139 ],
   alphaCSR[ 127 ][ 140 ],
   alphaCSR[ 127 ][ 141 ],
   alphaCSR[ 127 ][ 142 ],
   alphaCSR[ 127 ][ 143 ],
   alphaCSR[ 127 ][ 144 ],
   alphaCSR[ 127 ][ 145 ],
   alphaCSR[ 127 ][ 146 ],
   alphaCSR[ 127 ][ 147 ],
   alphaCSR[ 127 ][ 148 ],
   alphaCSR[ 127 ][ 149 ],
   alphaCSR[ 127 ][ 150 ],
   alphaCSR[ 127 ][ 151 ],
   alphaCSR[ 127 ][ 152 ],
   alphaCSR[ 127 ][ 153 ],
   alphaCSR[ 127 ][ 154 ],
   alphaCSR[ 127 ][ 155 ],
   alphaCSR[ 127 ][ 156 ],
   alphaCSR[ 127 ][ 157 ],
   alphaCSR[ 127 ][ 158 ],
   alphaCSR[ 127 ][ 159 ],
   alphaCSR[ 127 ][ 160 ],
   alphaCSR[ 127 ][ 161 ],
   alphaCSR[ 127 ][ 162 ],
   alphaCSR[ 127 ][ 163 ],
   alphaCSR[ 127 ][ 164 ],
   alphaCSR[ 127 ][ 165 ],
   alphaCSR[ 127 ][ 166 ],
   alphaCSR[ 127 ][ 167 ],
   alphaCSR[ 127 ][ 168 ],
   alphaCSR[ 127 ][ 169 ],
   alphaCSR[ 127 ][ 170 ],
   alphaCSR[ 127 ][ 171 ],
   alphaCSR[ 127 ][ 172 ],
   alphaCSR[ 127 ][ 173 ],
   alphaCSR[ 127 ][ 174 ],
   alphaCSR[ 127 ][ 175 ],
   alphaCSR[ 127 ][ 176 ],
   alphaCSR[ 127 ][ 177 ],
   alphaCSR[ 127 ][ 178 ],
   alphaCSR[ 127 ][ 179 ],
   alphaCSR[ 127 ][ 180 ],
   alphaCSR[ 127 ][ 181 ],
   alphaCSR[ 127 ][ 182 ],
   alphaCSR[ 127 ][ 183 ],
   alphaCSR[ 127 ][ 184 ],
   alphaCSR[ 127 ][ 185 ],
   alphaCSR[ 127 ][ 186 ],
   alphaCSR[ 127 ][ 187 ],
   alphaCSR[ 127 ][ 188 ],
   alphaCSR[ 127 ][ 189 ],
   alphaCSR[ 127 ][ 190 ],
   alphaCSR[ 127 ][ 191 ],
   alphaCSR[ 127 ][ 192 ],
   alphaCSR[ 127 ][ 193 ],
   alphaCSR[ 127 ][ 194 ],
   alphaCSR[ 127 ][ 195 ],
   alphaCSR[ 127 ][ 196 ],
   alphaCSR[ 127 ][ 197 ],
   alphaCSR[ 127 ][ 198 ],
   alphaCSR[ 127 ][ 199 ],
   alphaCSR[ 127 ][ 200 ],
   alphaCSR[ 127 ][ 201 ],
   alphaCSR[ 127 ][ 202 ],
   alphaCSR[ 127 ][ 203 ],
   alphaCSR[ 127 ][ 204 ],
   alphaCSR[ 127 ][ 205 ],
   alphaCSR[ 127 ][ 206 ],
   alphaCSR[ 127 ][ 207 ],
   alphaCSR[ 127 ][ 208 ],
   alphaCSR[ 127 ][ 209 ],
   alphaCSR[ 127 ][ 210 ],
   alphaCSR[ 127 ][ 211 ],
   alphaCSR[ 127 ][ 212 ],
   alphaCSR[ 127 ][ 213 ],
   alphaCSR[ 127 ][ 214 ],
   alphaCSR[ 127 ][ 215 ],
   alphaCSR[ 127 ][ 216 ],
   alphaCSR[ 127 ][ 217 ],
   alphaCSR[ 127 ][ 218 ],
   alphaCSR[ 127 ][ 219 ],
   alphaCSR[ 127 ][ 220 ],
   alphaCSR[ 127 ][ 221 ],
   alphaCSR[ 127 ][ 222 ],
   alphaCSR[ 127 ][ 223 ],
   alphaCSR[ 127 ][ 224 ],
   alphaCSR[ 127 ][ 225 ],
   alphaCSR[ 127 ][ 226 ],
   alphaCSR[ 127 ][ 227 ],
   alphaCSR[ 127 ][ 228 ],
   alphaCSR[ 127 ][ 229 ],
   alphaCSR[ 127 ][ 230 ],
   alphaCSR[ 127 ][ 231 ],
   alphaCSR[ 127 ][ 232 ],
   alphaCSR[ 127 ][ 233 ],
   alphaCSR[ 127 ][ 234 ],
   alphaCSR[ 127 ][ 235 ],
   alphaCSR[ 127 ][ 236 ],
   alphaCSR[ 127 ][ 237 ],
   alphaCSR[ 127 ][ 238 ],
   alphaCSR[ 127 ][ 239 ],
   alphaCSR[ 127 ][ 240 ],
   alphaCSR[ 127 ][ 241 ],
   alphaCSR[ 127 ][ 242 ],
   alphaCSR[ 127 ][ 243 ],
   alphaCSR[ 127 ][ 244 ],
   alphaCSR[ 127 ][ 245 ],
   alphaCSR[ 127 ][ 246 ],
   alphaCSR[ 127 ][ 247 ],
   alphaCSR[ 127 ][ 248 ],
   alphaCSR[ 127 ][ 249 ],
   alphaCSR[ 127 ][ 250 ],
   alphaCSR[ 127 ][ 251 ],
   alphaCSR[ 127 ][ 252 ],
   alphaCSR[ 127 ][ 253 ],
   alphaCSR[ 127 ][ 254 ],
   alphaCSR[ 127 ][ 255 ],
   alphaCSR[ 127 ][ 256 ],
   alphaCSR[ 127 ][ 257 ],
   alphaCSR[ 127 ][ 258 ],
   alphaCSR[ 127 ][ 259 ],
   alphaCSR[ 127 ][ 260 ],
   alphaCSR[ 127 ][ 261 ],
   alphaCSR[ 127 ][ 262 ],
   alphaCSR[ 127 ][ 263 ],
   alphaCSR[ 127 ][ 264 ],
   alphaCSR[ 127 ][ 265 ],
   alphaCSR[ 127 ][ 266 ],
   alphaCSR[ 127 ][ 267 ],
   alphaCSR[ 127 ][ 268 ],
   alphaCSR[ 127 ][ 269 ],
   alphaCSR[ 127 ][ 270 ],
   alphaCSR[ 127 ][ 271 ],
   alphaCSR[ 127 ][ 272 ],
   alphaCSR[ 127 ][ 273 ],
   alphaCSR[ 127 ][ 274 ],
   alphaCSR[ 127 ][ 275 ],
   alphaCSR[ 127 ][ 276 ],
   alphaCSR[ 127 ][ 277 ],
   alphaCSR[ 127 ][ 278 ],
   alphaCSR[ 127 ][ 279 ],
   alphaCSR[ 127 ][ 280 ],
   alphaCSR[ 127 ][ 281 ],
   alphaCSR[ 127 ][ 282 ],
   alphaCSR[ 127 ][ 283 ],
   alphaCSR[ 127 ][ 284 ],
   alphaCSR[ 127 ][ 285 ],
   alphaCSR[ 127 ][ 286 ],
   alphaCSR[ 127 ][ 287 ],
   alphaCSR[ 127 ][ 288 ],
   alphaCSR[ 127 ][ 289 ],
   alphaCSR[ 127 ][ 290 ],
   alphaCSR[ 127 ][ 291 ],
   alphaCSR[ 127 ][ 292 ],
   alphaCSR[ 127 ][ 293 ],
   alphaCSR[ 127 ][ 294 ],
   alphaCSR[ 127 ][ 295 ],
   alphaCSR[ 127 ][ 296 ],
   alphaCSR[ 127 ][ 297 ],
   alphaCSR[ 127 ][ 298 ],
   alphaCSR[ 127 ][ 299 ],
   alphaCSR[ 127 ][ 300 ],
   alphaCSR[ 127 ][ 301 ],
   alphaCSR[ 127 ][ 302 ],
   alphaCSR[ 127 ][ 303 ],
   alphaCSR[ 127 ][ 304 ],
   alphaCSR[ 127 ][ 305 ],
   alphaCSR[ 127 ][ 306 ],
   alphaCSR[ 127 ][ 307 ],
   alphaCSR[ 127 ][ 308 ],
   alphaCSR[ 127 ][ 309 ],
   alphaCSR[ 127 ][ 310 ],
   alphaCSR[ 127 ][ 311 ],
   alphaCSR[ 127 ][ 312 ],
   alphaCSR[ 127 ][ 313 ],
   alphaCSR[ 127 ][ 314 ],
   alphaCSR[ 127 ][ 315 ],
   alphaCSR[ 127 ][ 316 ],
   alphaCSR[ 127 ][ 317 ],
   alphaCSR[ 127 ][ 318 ],
   alphaCSR[ 127 ][ 319 ],
   alphaCSR[ 127 ][ 320 ],
   alphaCSR[ 127 ][ 321 ],
   alphaCSR[ 127 ][ 322 ],
   alphaCSR[ 127 ][ 323 ],
   alphaCSR[ 127 ][ 324 ],
   alphaCSR[ 127 ][ 325 ],
   alphaCSR[ 127 ][ 326 ],
   alphaCSR[ 127 ][ 327 ],
   alphaCSR[ 127 ][ 328 ],
   alphaCSR[ 127 ][ 329 ],
   alphaCSR[ 127 ][ 330 ],
   alphaCSR[ 127 ][ 331 ],
   alphaCSR[ 127 ][ 332 ],
   alphaCSR[ 127 ][ 333 ],
   alphaCSR[ 127 ][ 334 ],
   alphaCSR[ 127 ][ 335 ],
   alphaCSR[ 127 ][ 336 ],
   alphaCSR[ 127 ][ 337 ],
   alphaCSR[ 127 ][ 338 ],
   alphaCSR[ 127 ][ 339 ],
   alphaCSR[ 127 ][ 340 ],
   alphaCSR[ 127 ][ 341 ],
   alphaCSR[ 127 ][ 342 ],
   alphaCSR[ 127 ][ 343 ],
   alphaCSR[ 127 ][ 344 ],
   alphaCSR[ 127 ][ 345 ],
   alphaCSR[ 127 ][ 346 ],
   alphaCSR[ 127 ][ 347 ],
   alphaCSR[ 127 ][ 348 ],
   alphaCSR[ 127 ][ 349 ],
   alphaCSR[ 127 ][ 350 ],
   alphaCSR[ 127 ][ 351 ],
   alphaCSR[ 127 ][ 352 ],
   alphaCSR[ 127 ][ 353 ],
   alphaCSR[ 127 ][ 354 ],
   alphaCSR[ 127 ][ 355 ],
   alphaCSR[ 127 ][ 356 ],
   alphaCSR[ 127 ][ 357 ],
   alphaCSR[ 127 ][ 358 ],
   alphaCSR[ 127 ][ 359 ],
   alphaCSR[ 127 ][ 360 ],
   alphaCSR[ 127 ][ 361 ],
   alphaCSR[ 127 ][ 362 ],
   alphaCSR[ 127 ][ 363 ],
   alphaCSR[ 127 ][ 364 ],
   alphaCSR[ 127 ][ 365 ],
   alphaCSR[ 127 ][ 366 ],
   alphaCSR[ 127 ][ 367 ],
   alphaCSR[ 127 ][ 368 ],
   alphaCSR[ 127 ][ 369 ],
   alphaCSR[ 127 ][ 370 ],
   alphaCSR[ 127 ][ 371 ],
   alphaCSR[ 127 ][ 372 ],
   alphaCSR[ 127 ][ 373 ],
   alphaCSR[ 127 ][ 374 ],
   alphaCSR[ 127 ][ 375 ],
   alphaCSR[ 127 ][ 376 ],
   alphaCSR[ 127 ][ 377 ],
   alphaCSR[ 127 ][ 378 ],
   alphaCSR[ 127 ][ 379 ],
   alphaCSR[ 127 ][ 380 ],
   alphaCSR[ 127 ][ 381 ],
   alphaCSR[ 127 ][ 382 ],
   alphaCSR[ 127 ][ 383 ],
   alphaCSR[ 128 ][ 0 ],
   alphaCSR[ 128 ][ 1 ],
   alphaCSR[ 128 ][ 2 ],
   alphaCSR[ 128 ][ 3 ],
   alphaCSR[ 128 ][ 4 ],
   alphaCSR[ 128 ][ 5 ],
   alphaCSR[ 128 ][ 6 ],
   alphaCSR[ 128 ][ 7 ],
   alphaCSR[ 128 ][ 8 ],
   alphaCSR[ 128 ][ 9 ],
   alphaCSR[ 128 ][ 10 ],
   alphaCSR[ 128 ][ 11 ],
   alphaCSR[ 128 ][ 12 ],
   alphaCSR[ 128 ][ 13 ],
   alphaCSR[ 128 ][ 14 ],
   alphaCSR[ 128 ][ 15 ],
   alphaCSR[ 128 ][ 16 ],
   alphaCSR[ 128 ][ 17 ],
   alphaCSR[ 128 ][ 18 ],
   alphaCSR[ 128 ][ 19 ],
   alphaCSR[ 128 ][ 20 ],
   alphaCSR[ 128 ][ 21 ],
   alphaCSR[ 128 ][ 22 ],
   alphaCSR[ 128 ][ 23 ],
   alphaCSR[ 128 ][ 24 ],
   alphaCSR[ 128 ][ 25 ],
   alphaCSR[ 128 ][ 26 ],
   alphaCSR[ 128 ][ 27 ],
   alphaCSR[ 128 ][ 28 ],
   alphaCSR[ 128 ][ 29 ],
   alphaCSR[ 128 ][ 30 ],
   alphaCSR[ 128 ][ 31 ],
   alphaCSR[ 128 ][ 32 ],
   alphaCSR[ 128 ][ 33 ],
   alphaCSR[ 128 ][ 34 ],
   alphaCSR[ 128 ][ 35 ],
   alphaCSR[ 128 ][ 36 ],
   alphaCSR[ 128 ][ 37 ],
   alphaCSR[ 128 ][ 38 ],
   alphaCSR[ 128 ][ 39 ],
   alphaCSR[ 128 ][ 40 ],
   alphaCSR[ 128 ][ 41 ],
   alphaCSR[ 128 ][ 42 ],
   alphaCSR[ 128 ][ 43 ],
   alphaCSR[ 128 ][ 44 ],
   alphaCSR[ 128 ][ 45 ],
   alphaCSR[ 128 ][ 46 ],
   alphaCSR[ 128 ][ 47 ],
   alphaCSR[ 128 ][ 48 ],
   alphaCSR[ 128 ][ 49 ],
   alphaCSR[ 128 ][ 50 ],
   alphaCSR[ 128 ][ 51 ],
   alphaCSR[ 128 ][ 52 ],
   alphaCSR[ 128 ][ 53 ],
   alphaCSR[ 128 ][ 54 ],
   alphaCSR[ 128 ][ 55 ],
   alphaCSR[ 128 ][ 56 ],
   alphaCSR[ 128 ][ 57 ],
   alphaCSR[ 128 ][ 58 ],
   alphaCSR[ 128 ][ 59 ],
   alphaCSR[ 128 ][ 60 ],
   alphaCSR[ 128 ][ 61 ],
   alphaCSR[ 128 ][ 62 ],
   alphaCSR[ 128 ][ 63 ],
   alphaCSR[ 128 ][ 64 ],
   alphaCSR[ 128 ][ 65 ],
   alphaCSR[ 128 ][ 66 ],
   alphaCSR[ 128 ][ 67 ],
   alphaCSR[ 128 ][ 68 ],
   alphaCSR[ 128 ][ 69 ],
   alphaCSR[ 128 ][ 70 ],
   alphaCSR[ 128 ][ 71 ],
   alphaCSR[ 128 ][ 72 ],
   alphaCSR[ 128 ][ 73 ],
   alphaCSR[ 128 ][ 74 ],
   alphaCSR[ 128 ][ 75 ],
   alphaCSR[ 128 ][ 76 ],
   alphaCSR[ 128 ][ 77 ],
   alphaCSR[ 128 ][ 78 ],
   alphaCSR[ 128 ][ 79 ],
   alphaCSR[ 128 ][ 80 ],
   alphaCSR[ 128 ][ 81 ],
   alphaCSR[ 128 ][ 82 ],
   alphaCSR[ 128 ][ 83 ],
   alphaCSR[ 128 ][ 84 ],
   alphaCSR[ 128 ][ 85 ],
   alphaCSR[ 128 ][ 86 ],
   alphaCSR[ 128 ][ 87 ],
   alphaCSR[ 128 ][ 88 ],
   alphaCSR[ 128 ][ 89 ],
   alphaCSR[ 128 ][ 90 ],
   alphaCSR[ 128 ][ 91 ],
   alphaCSR[ 128 ][ 92 ],
   alphaCSR[ 128 ][ 93 ],
   alphaCSR[ 128 ][ 94 ],
   alphaCSR[ 128 ][ 95 ],
   alphaCSR[ 128 ][ 96 ],
   alphaCSR[ 128 ][ 97 ],
   alphaCSR[ 128 ][ 98 ],
   alphaCSR[ 128 ][ 99 ],
   alphaCSR[ 128 ][ 100 ],
   alphaCSR[ 128 ][ 101 ],
   alphaCSR[ 128 ][ 102 ],
   alphaCSR[ 128 ][ 103 ],
   alphaCSR[ 128 ][ 104 ],
   alphaCSR[ 128 ][ 105 ],
   alphaCSR[ 128 ][ 106 ],
   alphaCSR[ 128 ][ 107 ],
   alphaCSR[ 128 ][ 108 ],
   alphaCSR[ 128 ][ 109 ],
   alphaCSR[ 128 ][ 110 ],
   alphaCSR[ 128 ][ 111 ],
   alphaCSR[ 128 ][ 112 ],
   alphaCSR[ 128 ][ 113 ],
   alphaCSR[ 128 ][ 114 ],
   alphaCSR[ 128 ][ 115 ],
   alphaCSR[ 128 ][ 116 ],
   alphaCSR[ 128 ][ 117 ],
   alphaCSR[ 128 ][ 118 ],
   alphaCSR[ 128 ][ 119 ],
   alphaCSR[ 128 ][ 120 ],
   alphaCSR[ 128 ][ 121 ],
   alphaCSR[ 128 ][ 122 ],
   alphaCSR[ 128 ][ 123 ],
   alphaCSR[ 128 ][ 124 ],
   alphaCSR[ 128 ][ 125 ],
   alphaCSR[ 128 ][ 126 ],
   alphaCSR[ 128 ][ 127 ],
   alphaCSR[ 128 ][ 128 ],
   alphaCSR[ 128 ][ 129 ],
   alphaCSR[ 128 ][ 130 ],
   alphaCSR[ 128 ][ 131 ],
   alphaCSR[ 128 ][ 132 ],
   alphaCSR[ 128 ][ 133 ],
   alphaCSR[ 128 ][ 134 ],
   alphaCSR[ 128 ][ 135 ],
   alphaCSR[ 128 ][ 136 ],
   alphaCSR[ 128 ][ 137 ],
   alphaCSR[ 128 ][ 138 ],
   alphaCSR[ 128 ][ 139 ],
   alphaCSR[ 128 ][ 140 ],
   alphaCSR[ 128 ][ 141 ],
   alphaCSR[ 128 ][ 142 ],
   alphaCSR[ 128 ][ 143 ],
   alphaCSR[ 128 ][ 144 ],
   alphaCSR[ 128 ][ 145 ],
   alphaCSR[ 128 ][ 146 ],
   alphaCSR[ 128 ][ 147 ],
   alphaCSR[ 128 ][ 148 ],
   alphaCSR[ 128 ][ 149 ],
   alphaCSR[ 128 ][ 150 ],
   alphaCSR[ 128 ][ 151 ],
   alphaCSR[ 128 ][ 152 ],
   alphaCSR[ 128 ][ 153 ],
   alphaCSR[ 128 ][ 154 ],
   alphaCSR[ 128 ][ 155 ],
   alphaCSR[ 128 ][ 156 ],
   alphaCSR[ 128 ][ 157 ],
   alphaCSR[ 128 ][ 158 ],
   alphaCSR[ 128 ][ 159 ],
   alphaCSR[ 128 ][ 160 ],
   alphaCSR[ 128 ][ 161 ],
   alphaCSR[ 128 ][ 162 ],
   alphaCSR[ 128 ][ 163 ],
   alphaCSR[ 128 ][ 164 ],
   alphaCSR[ 128 ][ 165 ],
   alphaCSR[ 128 ][ 166 ],
   alphaCSR[ 128 ][ 167 ],
   alphaCSR[ 128 ][ 168 ],
   alphaCSR[ 128 ][ 169 ],
   alphaCSR[ 128 ][ 170 ],
   alphaCSR[ 128 ][ 171 ],
   alphaCSR[ 128 ][ 172 ],
   alphaCSR[ 128 ][ 173 ],
   alphaCSR[ 128 ][ 174 ],
   alphaCSR[ 128 ][ 175 ],
   alphaCSR[ 128 ][ 176 ],
   alphaCSR[ 128 ][ 177 ],
   alphaCSR[ 128 ][ 178 ],
   alphaCSR[ 128 ][ 179 ],
   alphaCSR[ 128 ][ 180 ],
   alphaCSR[ 128 ][ 181 ],
   alphaCSR[ 128 ][ 182 ],
   alphaCSR[ 128 ][ 183 ],
   alphaCSR[ 128 ][ 184 ],
   alphaCSR[ 128 ][ 185 ],
   alphaCSR[ 128 ][ 186 ],
   alphaCSR[ 128 ][ 187 ],
   alphaCSR[ 128 ][ 188 ],
   alphaCSR[ 128 ][ 189 ],
   alphaCSR[ 128 ][ 190 ],
   alphaCSR[ 128 ][ 191 ],
   alphaCSR[ 128 ][ 192 ],
   alphaCSR[ 128 ][ 193 ],
   alphaCSR[ 128 ][ 194 ],
   alphaCSR[ 128 ][ 195 ],
   alphaCSR[ 128 ][ 196 ],
   alphaCSR[ 128 ][ 197 ],
   alphaCSR[ 128 ][ 198 ],
   alphaCSR[ 128 ][ 199 ],
   alphaCSR[ 128 ][ 200 ],
   alphaCSR[ 128 ][ 201 ],
   alphaCSR[ 128 ][ 202 ],
   alphaCSR[ 128 ][ 203 ],
   alphaCSR[ 128 ][ 204 ],
   alphaCSR[ 128 ][ 205 ],
   alphaCSR[ 128 ][ 206 ],
   alphaCSR[ 128 ][ 207 ],
   alphaCSR[ 128 ][ 208 ],
   alphaCSR[ 128 ][ 209 ],
   alphaCSR[ 128 ][ 210 ],
   alphaCSR[ 128 ][ 211 ],
   alphaCSR[ 128 ][ 212 ],
   alphaCSR[ 128 ][ 213 ],
   alphaCSR[ 128 ][ 214 ],
   alphaCSR[ 128 ][ 215 ],
   alphaCSR[ 128 ][ 216 ],
   alphaCSR[ 128 ][ 217 ],
   alphaCSR[ 128 ][ 218 ],
   alphaCSR[ 128 ][ 219 ],
   alphaCSR[ 128 ][ 220 ],
   alphaCSR[ 128 ][ 221 ],
   alphaCSR[ 128 ][ 222 ],
   alphaCSR[ 128 ][ 223 ],
   alphaCSR[ 128 ][ 224 ],
   alphaCSR[ 128 ][ 225 ],
   alphaCSR[ 128 ][ 226 ],
   alphaCSR[ 128 ][ 227 ],
   alphaCSR[ 128 ][ 228 ],
   alphaCSR[ 128 ][ 229 ],
   alphaCSR[ 128 ][ 230 ],
   alphaCSR[ 128 ][ 231 ],
   alphaCSR[ 128 ][ 232 ],
   alphaCSR[ 128 ][ 233 ],
   alphaCSR[ 128 ][ 234 ],
   alphaCSR[ 128 ][ 235 ],
   alphaCSR[ 128 ][ 236 ],
   alphaCSR[ 128 ][ 237 ],
   alphaCSR[ 128 ][ 238 ],
   alphaCSR[ 128 ][ 239 ],
   alphaCSR[ 128 ][ 240 ],
   alphaCSR[ 128 ][ 241 ],
   alphaCSR[ 128 ][ 242 ],
   alphaCSR[ 128 ][ 243 ],
   alphaCSR[ 128 ][ 244 ],
   alphaCSR[ 128 ][ 245 ],
   alphaCSR[ 128 ][ 246 ],
   alphaCSR[ 128 ][ 247 ],
   alphaCSR[ 128 ][ 248 ],
   alphaCSR[ 128 ][ 249 ],
   alphaCSR[ 128 ][ 250 ],
   alphaCSR[ 128 ][ 251 ],
   alphaCSR[ 128 ][ 252 ],
   alphaCSR[ 128 ][ 253 ],
   alphaCSR[ 128 ][ 254 ],
   alphaCSR[ 128 ][ 255 ],
   alphaCSR[ 128 ][ 256 ],
   alphaCSR[ 128 ][ 257 ],
   alphaCSR[ 128 ][ 258 ],
   alphaCSR[ 128 ][ 259 ],
   alphaCSR[ 128 ][ 260 ],
   alphaCSR[ 128 ][ 261 ],
   alphaCSR[ 128 ][ 262 ],
   alphaCSR[ 128 ][ 263 ],
   alphaCSR[ 128 ][ 264 ],
   alphaCSR[ 128 ][ 265 ],
   alphaCSR[ 128 ][ 266 ],
   alphaCSR[ 128 ][ 267 ],
   alphaCSR[ 128 ][ 268 ],
   alphaCSR[ 128 ][ 269 ],
   alphaCSR[ 128 ][ 270 ],
   alphaCSR[ 128 ][ 271 ],
   alphaCSR[ 128 ][ 272 ],
   alphaCSR[ 128 ][ 273 ],
   alphaCSR[ 128 ][ 274 ],
   alphaCSR[ 128 ][ 275 ],
   alphaCSR[ 128 ][ 276 ],
   alphaCSR[ 128 ][ 277 ],
   alphaCSR[ 128 ][ 278 ],
   alphaCSR[ 128 ][ 279 ],
   alphaCSR[ 128 ][ 280 ],
   alphaCSR[ 128 ][ 281 ],
   alphaCSR[ 128 ][ 282 ],
   alphaCSR[ 128 ][ 283 ],
   alphaCSR[ 128 ][ 284 ],
   alphaCSR[ 128 ][ 285 ],
   alphaCSR[ 128 ][ 286 ],
   alphaCSR[ 128 ][ 287 ],
   alphaCSR[ 128 ][ 288 ],
   alphaCSR[ 128 ][ 289 ],
   alphaCSR[ 128 ][ 290 ],
   alphaCSR[ 128 ][ 291 ],
   alphaCSR[ 128 ][ 292 ],
   alphaCSR[ 128 ][ 293 ],
   alphaCSR[ 128 ][ 294 ],
   alphaCSR[ 128 ][ 295 ],
   alphaCSR[ 128 ][ 296 ],
   alphaCSR[ 128 ][ 297 ],
   alphaCSR[ 128 ][ 298 ],
   alphaCSR[ 128 ][ 299 ],
   alphaCSR[ 128 ][ 300 ],
   alphaCSR[ 128 ][ 301 ],
   alphaCSR[ 128 ][ 302 ],
   alphaCSR[ 128 ][ 303 ],
   alphaCSR[ 128 ][ 304 ],
   alphaCSR[ 128 ][ 305 ],
   alphaCSR[ 128 ][ 306 ],
   alphaCSR[ 128 ][ 307 ],
   alphaCSR[ 128 ][ 308 ],
   alphaCSR[ 128 ][ 309 ],
   alphaCSR[ 128 ][ 310 ],
   alphaCSR[ 128 ][ 311 ],
   alphaCSR[ 128 ][ 312 ],
   alphaCSR[ 128 ][ 313 ],
   alphaCSR[ 128 ][ 314 ],
   alphaCSR[ 128 ][ 315 ],
   alphaCSR[ 128 ][ 316 ],
   alphaCSR[ 128 ][ 317 ],
   alphaCSR[ 128 ][ 318 ],
   alphaCSR[ 128 ][ 319 ],
   alphaCSR[ 128 ][ 320 ],
   alphaCSR[ 128 ][ 321 ],
   alphaCSR[ 128 ][ 322 ],
   alphaCSR[ 128 ][ 323 ],
   alphaCSR[ 128 ][ 324 ],
   alphaCSR[ 128 ][ 325 ],
   alphaCSR[ 128 ][ 326 ],
   alphaCSR[ 128 ][ 327 ],
   alphaCSR[ 128 ][ 328 ],
   alphaCSR[ 128 ][ 329 ],
   alphaCSR[ 128 ][ 330 ],
   alphaCSR[ 128 ][ 331 ],
   alphaCSR[ 128 ][ 332 ],
   alphaCSR[ 128 ][ 333 ],
   alphaCSR[ 128 ][ 334 ],
   alphaCSR[ 128 ][ 335 ],
   alphaCSR[ 128 ][ 336 ],
   alphaCSR[ 128 ][ 337 ],
   alphaCSR[ 128 ][ 338 ],
   alphaCSR[ 128 ][ 339 ],
   alphaCSR[ 128 ][ 340 ],
   alphaCSR[ 128 ][ 341 ],
   alphaCSR[ 128 ][ 342 ],
   alphaCSR[ 128 ][ 343 ],
   alphaCSR[ 128 ][ 344 ],
   alphaCSR[ 128 ][ 345 ],
   alphaCSR[ 128 ][ 346 ],
   alphaCSR[ 128 ][ 347 ],
   alphaCSR[ 128 ][ 348 ],
   alphaCSR[ 128 ][ 349 ],
   alphaCSR[ 128 ][ 350 ],
   alphaCSR[ 128 ][ 351 ],
   alphaCSR[ 128 ][ 352 ],
   alphaCSR[ 128 ][ 353 ],
   alphaCSR[ 128 ][ 354 ],
   alphaCSR[ 128 ][ 355 ],
   alphaCSR[ 128 ][ 356 ],
   alphaCSR[ 128 ][ 357 ],
   alphaCSR[ 128 ][ 358 ],
   alphaCSR[ 128 ][ 359 ],
   alphaCSR[ 128 ][ 360 ],
   alphaCSR[ 128 ][ 361 ],
   alphaCSR[ 128 ][ 362 ],
   alphaCSR[ 128 ][ 363 ],
   alphaCSR[ 128 ][ 364 ],
   alphaCSR[ 128 ][ 365 ],
   alphaCSR[ 128 ][ 366 ],
   alphaCSR[ 128 ][ 367 ],
   alphaCSR[ 128 ][ 368 ],
   alphaCSR[ 128 ][ 369 ],
   alphaCSR[ 128 ][ 370 ],
   alphaCSR[ 128 ][ 371 ],
   alphaCSR[ 128 ][ 372 ],
   alphaCSR[ 128 ][ 373 ],
   alphaCSR[ 128 ][ 374 ],
   alphaCSR[ 128 ][ 375 ],
   alphaCSR[ 128 ][ 376 ],
   alphaCSR[ 128 ][ 377 ],
   alphaCSR[ 128 ][ 378 ],
   alphaCSR[ 128 ][ 379 ],
   alphaCSR[ 128 ][ 380 ],
   alphaCSR[ 128 ][ 381 ],
   alphaCSR[ 128 ][ 382 ],
   alphaCSR[ 128 ][ 383 ],
   alphaCSR[ 129 ][ 0 ],
   alphaCSR[ 129 ][ 1 ],
   alphaCSR[ 129 ][ 2 ],
   alphaCSR[ 129 ][ 3 ],
   alphaCSR[ 129 ][ 4 ],
   alphaCSR[ 129 ][ 5 ],
   alphaCSR[ 129 ][ 6 ],
   alphaCSR[ 129 ][ 7 ],
   alphaCSR[ 129 ][ 8 ],
   alphaCSR[ 129 ][ 9 ],
   alphaCSR[ 129 ][ 10 ],
   alphaCSR[ 129 ][ 11 ],
   alphaCSR[ 129 ][ 12 ],
   alphaCSR[ 129 ][ 13 ],
   alphaCSR[ 129 ][ 14 ],
   alphaCSR[ 129 ][ 15 ],
   alphaCSR[ 129 ][ 16 ],
   alphaCSR[ 129 ][ 17 ],
   alphaCSR[ 129 ][ 18 ],
   alphaCSR[ 129 ][ 19 ],
   alphaCSR[ 129 ][ 20 ],
   alphaCSR[ 129 ][ 21 ],
   alphaCSR[ 129 ][ 22 ],
   alphaCSR[ 129 ][ 23 ],
   alphaCSR[ 129 ][ 24 ],
   alphaCSR[ 129 ][ 25 ],
   alphaCSR[ 129 ][ 26 ],
   alphaCSR[ 129 ][ 27 ],
   alphaCSR[ 129 ][ 28 ],
   alphaCSR[ 129 ][ 29 ],
   alphaCSR[ 129 ][ 30 ],
   alphaCSR[ 129 ][ 31 ],
   alphaCSR[ 129 ][ 32 ],
   alphaCSR[ 129 ][ 33 ],
   alphaCSR[ 129 ][ 34 ],
   alphaCSR[ 129 ][ 35 ],
   alphaCSR[ 129 ][ 36 ],
   alphaCSR[ 129 ][ 37 ],
   alphaCSR[ 129 ][ 38 ],
   alphaCSR[ 129 ][ 39 ],
   alphaCSR[ 129 ][ 40 ],
   alphaCSR[ 129 ][ 41 ],
   alphaCSR[ 129 ][ 42 ],
   alphaCSR[ 129 ][ 43 ],
   alphaCSR[ 129 ][ 44 ],
   alphaCSR[ 129 ][ 45 ],
   alphaCSR[ 129 ][ 46 ],
   alphaCSR[ 129 ][ 47 ],
   alphaCSR[ 129 ][ 48 ],
   alphaCSR[ 129 ][ 49 ],
   alphaCSR[ 129 ][ 50 ],
   alphaCSR[ 129 ][ 51 ],
   alphaCSR[ 129 ][ 52 ],
   alphaCSR[ 129 ][ 53 ],
   alphaCSR[ 129 ][ 54 ],
   alphaCSR[ 129 ][ 55 ],
   alphaCSR[ 129 ][ 56 ],
   alphaCSR[ 129 ][ 57 ],
   alphaCSR[ 129 ][ 58 ],
   alphaCSR[ 129 ][ 59 ],
   alphaCSR[ 129 ][ 60 ],
   alphaCSR[ 129 ][ 61 ],
   alphaCSR[ 129 ][ 62 ],
   alphaCSR[ 129 ][ 63 ],
   alphaCSR[ 129 ][ 64 ],
   alphaCSR[ 129 ][ 65 ],
   alphaCSR[ 129 ][ 66 ],
   alphaCSR[ 129 ][ 67 ],
   alphaCSR[ 129 ][ 68 ],
   alphaCSR[ 129 ][ 69 ],
   alphaCSR[ 129 ][ 70 ],
   alphaCSR[ 129 ][ 71 ],
   alphaCSR[ 129 ][ 72 ],
   alphaCSR[ 129 ][ 73 ],
   alphaCSR[ 129 ][ 74 ],
   alphaCSR[ 129 ][ 75 ],
   alphaCSR[ 129 ][ 76 ],
   alphaCSR[ 129 ][ 77 ],
   alphaCSR[ 129 ][ 78 ],
   alphaCSR[ 129 ][ 79 ],
   alphaCSR[ 129 ][ 80 ],
   alphaCSR[ 129 ][ 81 ],
   alphaCSR[ 129 ][ 82 ],
   alphaCSR[ 129 ][ 83 ],
   alphaCSR[ 129 ][ 84 ],
   alphaCSR[ 129 ][ 85 ],
   alphaCSR[ 129 ][ 86 ],
   alphaCSR[ 129 ][ 87 ],
   alphaCSR[ 129 ][ 88 ],
   alphaCSR[ 129 ][ 89 ],
   alphaCSR[ 129 ][ 90 ],
   alphaCSR[ 129 ][ 91 ],
   alphaCSR[ 129 ][ 92 ],
   alphaCSR[ 129 ][ 93 ],
   alphaCSR[ 129 ][ 94 ],
   alphaCSR[ 129 ][ 95 ],
   alphaCSR[ 129 ][ 96 ],
   alphaCSR[ 129 ][ 97 ],
   alphaCSR[ 129 ][ 98 ],
   alphaCSR[ 129 ][ 99 ],
   alphaCSR[ 129 ][ 100 ],
   alphaCSR[ 129 ][ 101 ],
   alphaCSR[ 129 ][ 102 ],
   alphaCSR[ 129 ][ 103 ],
   alphaCSR[ 129 ][ 104 ],
   alphaCSR[ 129 ][ 105 ],
   alphaCSR[ 129 ][ 106 ],
   alphaCSR[ 129 ][ 107 ],
   alphaCSR[ 129 ][ 108 ],
   alphaCSR[ 129 ][ 109 ],
   alphaCSR[ 129 ][ 110 ],
   alphaCSR[ 129 ][ 111 ],
   alphaCSR[ 129 ][ 112 ],
   alphaCSR[ 129 ][ 113 ],
   alphaCSR[ 129 ][ 114 ],
   alphaCSR[ 129 ][ 115 ],
   alphaCSR[ 129 ][ 116 ],
   alphaCSR[ 129 ][ 117 ],
   alphaCSR[ 129 ][ 118 ],
   alphaCSR[ 129 ][ 119 ],
   alphaCSR[ 129 ][ 120 ],
   alphaCSR[ 129 ][ 121 ],
   alphaCSR[ 129 ][ 122 ],
   alphaCSR[ 129 ][ 123 ],
   alphaCSR[ 129 ][ 124 ],
   alphaCSR[ 129 ][ 125 ],
   alphaCSR[ 129 ][ 126 ],
   alphaCSR[ 129 ][ 127 ],
   alphaCSR[ 129 ][ 128 ],
   alphaCSR[ 129 ][ 129 ],
   alphaCSR[ 129 ][ 130 ],
   alphaCSR[ 129 ][ 131 ],
   alphaCSR[ 129 ][ 132 ],
   alphaCSR[ 129 ][ 133 ],
   alphaCSR[ 129 ][ 134 ],
   alphaCSR[ 129 ][ 135 ],
   alphaCSR[ 129 ][ 136 ],
   alphaCSR[ 129 ][ 137 ],
   alphaCSR[ 129 ][ 138 ],
   alphaCSR[ 129 ][ 139 ],
   alphaCSR[ 129 ][ 140 ],
   alphaCSR[ 129 ][ 141 ],
   alphaCSR[ 129 ][ 142 ],
   alphaCSR[ 129 ][ 143 ],
   alphaCSR[ 129 ][ 144 ],
   alphaCSR[ 129 ][ 145 ],
   alphaCSR[ 129 ][ 146 ],
   alphaCSR[ 129 ][ 147 ],
   alphaCSR[ 129 ][ 148 ],
   alphaCSR[ 129 ][ 149 ],
   alphaCSR[ 129 ][ 150 ],
   alphaCSR[ 129 ][ 151 ],
   alphaCSR[ 129 ][ 152 ],
   alphaCSR[ 129 ][ 153 ],
   alphaCSR[ 129 ][ 154 ],
   alphaCSR[ 129 ][ 155 ],
   alphaCSR[ 129 ][ 156 ],
   alphaCSR[ 129 ][ 157 ],
   alphaCSR[ 129 ][ 158 ],
   alphaCSR[ 129 ][ 159 ],
   alphaCSR[ 129 ][ 160 ],
   alphaCSR[ 129 ][ 161 ],
   alphaCSR[ 129 ][ 162 ],
   alphaCSR[ 129 ][ 163 ],
   alphaCSR[ 129 ][ 164 ],
   alphaCSR[ 129 ][ 165 ],
   alphaCSR[ 129 ][ 166 ],
   alphaCSR[ 129 ][ 167 ],
   alphaCSR[ 129 ][ 168 ],
   alphaCSR[ 129 ][ 169 ],
   alphaCSR[ 129 ][ 170 ],
   alphaCSR[ 129 ][ 171 ],
   alphaCSR[ 129 ][ 172 ],
   alphaCSR[ 129 ][ 173 ],
   alphaCSR[ 129 ][ 174 ],
   alphaCSR[ 129 ][ 175 ],
   alphaCSR[ 129 ][ 176 ],
   alphaCSR[ 129 ][ 177 ],
   alphaCSR[ 129 ][ 178 ],
   alphaCSR[ 129 ][ 179 ],
   alphaCSR[ 129 ][ 180 ],
   alphaCSR[ 129 ][ 181 ],
   alphaCSR[ 129 ][ 182 ],
   alphaCSR[ 129 ][ 183 ],
   alphaCSR[ 129 ][ 184 ],
   alphaCSR[ 129 ][ 185 ],
   alphaCSR[ 129 ][ 186 ],
   alphaCSR[ 129 ][ 187 ],
   alphaCSR[ 129 ][ 188 ],
   alphaCSR[ 129 ][ 189 ],
   alphaCSR[ 129 ][ 190 ],
   alphaCSR[ 129 ][ 191 ],
   alphaCSR[ 129 ][ 192 ],
   alphaCSR[ 129 ][ 193 ],
   alphaCSR[ 129 ][ 194 ],
   alphaCSR[ 129 ][ 195 ],
   alphaCSR[ 129 ][ 196 ],
   alphaCSR[ 129 ][ 197 ],
   alphaCSR[ 129 ][ 198 ],
   alphaCSR[ 129 ][ 199 ],
   alphaCSR[ 129 ][ 200 ],
   alphaCSR[ 129 ][ 201 ],
   alphaCSR[ 129 ][ 202 ],
   alphaCSR[ 129 ][ 203 ],
   alphaCSR[ 129 ][ 204 ],
   alphaCSR[ 129 ][ 205 ],
   alphaCSR[ 129 ][ 206 ],
   alphaCSR[ 129 ][ 207 ],
   alphaCSR[ 129 ][ 208 ],
   alphaCSR[ 129 ][ 209 ],
   alphaCSR[ 129 ][ 210 ],
   alphaCSR[ 129 ][ 211 ],
   alphaCSR[ 129 ][ 212 ],
   alphaCSR[ 129 ][ 213 ],
   alphaCSR[ 129 ][ 214 ],
   alphaCSR[ 129 ][ 215 ],
   alphaCSR[ 129 ][ 216 ],
   alphaCSR[ 129 ][ 217 ],
   alphaCSR[ 129 ][ 218 ],
   alphaCSR[ 129 ][ 219 ],
   alphaCSR[ 129 ][ 220 ],
   alphaCSR[ 129 ][ 221 ],
   alphaCSR[ 129 ][ 222 ],
   alphaCSR[ 129 ][ 223 ],
   alphaCSR[ 129 ][ 224 ],
   alphaCSR[ 129 ][ 225 ],
   alphaCSR[ 129 ][ 226 ],
   alphaCSR[ 129 ][ 227 ],
   alphaCSR[ 129 ][ 228 ],
   alphaCSR[ 129 ][ 229 ],
   alphaCSR[ 129 ][ 230 ],
   alphaCSR[ 129 ][ 231 ],
   alphaCSR[ 129 ][ 232 ],
   alphaCSR[ 129 ][ 233 ],
   alphaCSR[ 129 ][ 234 ],
   alphaCSR[ 129 ][ 235 ],
   alphaCSR[ 129 ][ 236 ],
   alphaCSR[ 129 ][ 237 ],
   alphaCSR[ 129 ][ 238 ],
   alphaCSR[ 129 ][ 239 ],
   alphaCSR[ 129 ][ 240 ],
   alphaCSR[ 129 ][ 241 ],
   alphaCSR[ 129 ][ 242 ],
   alphaCSR[ 129 ][ 243 ],
   alphaCSR[ 129 ][ 244 ],
   alphaCSR[ 129 ][ 245 ],
   alphaCSR[ 129 ][ 246 ],
   alphaCSR[ 129 ][ 247 ],
   alphaCSR[ 129 ][ 248 ],
   alphaCSR[ 129 ][ 249 ],
   alphaCSR[ 129 ][ 250 ],
   alphaCSR[ 129 ][ 251 ],
   alphaCSR[ 129 ][ 252 ],
   alphaCSR[ 129 ][ 253 ],
   alphaCSR[ 129 ][ 254 ],
   alphaCSR[ 129 ][ 255 ],
   alphaCSR[ 129 ][ 256 ],
   alphaCSR[ 129 ][ 257 ],
   alphaCSR[ 129 ][ 258 ],
   alphaCSR[ 129 ][ 259 ],
   alphaCSR[ 129 ][ 260 ],
   alphaCSR[ 129 ][ 261 ],
   alphaCSR[ 129 ][ 262 ],
   alphaCSR[ 129 ][ 263 ],
   alphaCSR[ 129 ][ 264 ],
   alphaCSR[ 129 ][ 265 ],
   alphaCSR[ 129 ][ 266 ],
   alphaCSR[ 129 ][ 267 ],
   alphaCSR[ 129 ][ 268 ],
   alphaCSR[ 129 ][ 269 ],
   alphaCSR[ 129 ][ 270 ],
   alphaCSR[ 129 ][ 271 ],
   alphaCSR[ 129 ][ 272 ],
   alphaCSR[ 129 ][ 273 ],
   alphaCSR[ 129 ][ 274 ],
   alphaCSR[ 129 ][ 275 ],
   alphaCSR[ 129 ][ 276 ],
   alphaCSR[ 129 ][ 277 ],
   alphaCSR[ 129 ][ 278 ],
   alphaCSR[ 129 ][ 279 ],
   alphaCSR[ 129 ][ 280 ],
   alphaCSR[ 129 ][ 281 ],
   alphaCSR[ 129 ][ 282 ],
   alphaCSR[ 129 ][ 283 ],
   alphaCSR[ 129 ][ 284 ],
   alphaCSR[ 129 ][ 285 ],
   alphaCSR[ 129 ][ 286 ],
   alphaCSR[ 129 ][ 287 ],
   alphaCSR[ 129 ][ 288 ],
   alphaCSR[ 129 ][ 289 ],
   alphaCSR[ 129 ][ 290 ],
   alphaCSR[ 129 ][ 291 ],
   alphaCSR[ 129 ][ 292 ],
   alphaCSR[ 129 ][ 293 ],
   alphaCSR[ 129 ][ 294 ],
   alphaCSR[ 129 ][ 295 ],
   alphaCSR[ 129 ][ 296 ],
   alphaCSR[ 129 ][ 297 ],
   alphaCSR[ 129 ][ 298 ],
   alphaCSR[ 129 ][ 299 ],
   alphaCSR[ 129 ][ 300 ],
   alphaCSR[ 129 ][ 301 ],
   alphaCSR[ 129 ][ 302 ],
   alphaCSR[ 129 ][ 303 ],
   alphaCSR[ 129 ][ 304 ],
   alphaCSR[ 129 ][ 305 ],
   alphaCSR[ 129 ][ 306 ],
   alphaCSR[ 129 ][ 307 ],
   alphaCSR[ 129 ][ 308 ],
   alphaCSR[ 129 ][ 309 ],
   alphaCSR[ 129 ][ 310 ],
   alphaCSR[ 129 ][ 311 ],
   alphaCSR[ 129 ][ 312 ],
   alphaCSR[ 129 ][ 313 ],
   alphaCSR[ 129 ][ 314 ],
   alphaCSR[ 129 ][ 315 ],
   alphaCSR[ 129 ][ 316 ],
   alphaCSR[ 129 ][ 317 ],
   alphaCSR[ 129 ][ 318 ],
   alphaCSR[ 129 ][ 319 ],
   alphaCSR[ 129 ][ 320 ],
   alphaCSR[ 129 ][ 321 ],
   alphaCSR[ 129 ][ 322 ],
   alphaCSR[ 129 ][ 323 ],
   alphaCSR[ 129 ][ 324 ],
   alphaCSR[ 129 ][ 325 ],
   alphaCSR[ 129 ][ 326 ],
   alphaCSR[ 129 ][ 327 ],
   alphaCSR[ 129 ][ 328 ],
   alphaCSR[ 129 ][ 329 ],
   alphaCSR[ 129 ][ 330 ],
   alphaCSR[ 129 ][ 331 ],
   alphaCSR[ 129 ][ 332 ],
   alphaCSR[ 129 ][ 333 ],
   alphaCSR[ 129 ][ 334 ],
   alphaCSR[ 129 ][ 335 ],
   alphaCSR[ 129 ][ 336 ],
   alphaCSR[ 129 ][ 337 ],
   alphaCSR[ 129 ][ 338 ],
   alphaCSR[ 129 ][ 339 ],
   alphaCSR[ 129 ][ 340 ],
   alphaCSR[ 129 ][ 341 ],
   alphaCSR[ 129 ][ 342 ],
   alphaCSR[ 129 ][ 343 ],
   alphaCSR[ 129 ][ 344 ],
   alphaCSR[ 129 ][ 345 ],
   alphaCSR[ 129 ][ 346 ],
   alphaCSR[ 129 ][ 347 ],
   alphaCSR[ 129 ][ 348 ],
   alphaCSR[ 129 ][ 349 ],
   alphaCSR[ 129 ][ 350 ],
   alphaCSR[ 129 ][ 351 ],
   alphaCSR[ 129 ][ 352 ],
   alphaCSR[ 129 ][ 353 ],
   alphaCSR[ 129 ][ 354 ],
   alphaCSR[ 129 ][ 355 ],
   alphaCSR[ 129 ][ 356 ],
   alphaCSR[ 129 ][ 357 ],
   alphaCSR[ 129 ][ 358 ],
   alphaCSR[ 129 ][ 359 ],
   alphaCSR[ 129 ][ 360 ],
   alphaCSR[ 129 ][ 361 ],
   alphaCSR[ 129 ][ 362 ],
   alphaCSR[ 129 ][ 363 ],
   alphaCSR[ 129 ][ 364 ],
   alphaCSR[ 129 ][ 365 ],
   alphaCSR[ 129 ][ 366 ],
   alphaCSR[ 129 ][ 367 ],
   alphaCSR[ 129 ][ 368 ],
   alphaCSR[ 129 ][ 369 ],
   alphaCSR[ 129 ][ 370 ],
   alphaCSR[ 129 ][ 371 ],
   alphaCSR[ 129 ][ 372 ],
   alphaCSR[ 129 ][ 373 ],
   alphaCSR[ 129 ][ 374 ],
   alphaCSR[ 129 ][ 375 ],
   alphaCSR[ 129 ][ 376 ],
   alphaCSR[ 129 ][ 377 ],
   alphaCSR[ 129 ][ 378 ],
   alphaCSR[ 129 ][ 379 ],
   alphaCSR[ 129 ][ 380 ],
   alphaCSR[ 129 ][ 381 ],
   alphaCSR[ 129 ][ 382 ],
   alphaCSR[ 129 ][ 383 ],
   alphaCSR[ 130 ][ 0 ],
   alphaCSR[ 130 ][ 1 ],
   alphaCSR[ 130 ][ 2 ],
   alphaCSR[ 130 ][ 3 ],
   alphaCSR[ 130 ][ 4 ],
   alphaCSR[ 130 ][ 5 ],
   alphaCSR[ 130 ][ 6 ],
   alphaCSR[ 130 ][ 7 ],
   alphaCSR[ 130 ][ 8 ],
   alphaCSR[ 130 ][ 9 ],
   alphaCSR[ 130 ][ 10 ],
   alphaCSR[ 130 ][ 11 ],
   alphaCSR[ 130 ][ 12 ],
   alphaCSR[ 130 ][ 13 ],
   alphaCSR[ 130 ][ 14 ],
   alphaCSR[ 130 ][ 15 ],
   alphaCSR[ 130 ][ 16 ],
   alphaCSR[ 130 ][ 17 ],
   alphaCSR[ 130 ][ 18 ],
   alphaCSR[ 130 ][ 19 ],
   alphaCSR[ 130 ][ 20 ],
   alphaCSR[ 130 ][ 21 ],
   alphaCSR[ 130 ][ 22 ],
   alphaCSR[ 130 ][ 23 ],
   alphaCSR[ 130 ][ 24 ],
   alphaCSR[ 130 ][ 25 ],
   alphaCSR[ 130 ][ 26 ],
   alphaCSR[ 130 ][ 27 ],
   alphaCSR[ 130 ][ 28 ],
   alphaCSR[ 130 ][ 29 ],
   alphaCSR[ 130 ][ 30 ],
   alphaCSR[ 130 ][ 31 ],
   alphaCSR[ 130 ][ 32 ],
   alphaCSR[ 130 ][ 33 ],
   alphaCSR[ 130 ][ 34 ],
   alphaCSR[ 130 ][ 35 ],
   alphaCSR[ 130 ][ 36 ],
   alphaCSR[ 130 ][ 37 ],
   alphaCSR[ 130 ][ 38 ],
   alphaCSR[ 130 ][ 39 ],
   alphaCSR[ 130 ][ 40 ],
   alphaCSR[ 130 ][ 41 ],
   alphaCSR[ 130 ][ 42 ],
   alphaCSR[ 130 ][ 43 ],
   alphaCSR[ 130 ][ 44 ],
   alphaCSR[ 130 ][ 45 ],
   alphaCSR[ 130 ][ 46 ],
   alphaCSR[ 130 ][ 47 ],
   alphaCSR[ 130 ][ 48 ],
   alphaCSR[ 130 ][ 49 ],
   alphaCSR[ 130 ][ 50 ],
   alphaCSR[ 130 ][ 51 ],
   alphaCSR[ 130 ][ 52 ],
   alphaCSR[ 130 ][ 53 ],
   alphaCSR[ 130 ][ 54 ],
   alphaCSR[ 130 ][ 55 ],
   alphaCSR[ 130 ][ 56 ],
   alphaCSR[ 130 ][ 57 ],
   alphaCSR[ 130 ][ 58 ],
   alphaCSR[ 130 ][ 59 ],
   alphaCSR[ 130 ][ 60 ],
   alphaCSR[ 130 ][ 61 ],
   alphaCSR[ 130 ][ 62 ],
   alphaCSR[ 130 ][ 63 ],
   alphaCSR[ 130 ][ 64 ],
   alphaCSR[ 130 ][ 65 ],
   alphaCSR[ 130 ][ 66 ],
   alphaCSR[ 130 ][ 67 ],
   alphaCSR[ 130 ][ 68 ],
   alphaCSR[ 130 ][ 69 ],
   alphaCSR[ 130 ][ 70 ],
   alphaCSR[ 130 ][ 71 ],
   alphaCSR[ 130 ][ 72 ],
   alphaCSR[ 130 ][ 73 ],
   alphaCSR[ 130 ][ 74 ],
   alphaCSR[ 130 ][ 75 ],
   alphaCSR[ 130 ][ 76 ],
   alphaCSR[ 130 ][ 77 ],
   alphaCSR[ 130 ][ 78 ],
   alphaCSR[ 130 ][ 79 ],
   alphaCSR[ 130 ][ 80 ],
   alphaCSR[ 130 ][ 81 ],
   alphaCSR[ 130 ][ 82 ],
   alphaCSR[ 130 ][ 83 ],
   alphaCSR[ 130 ][ 84 ],
   alphaCSR[ 130 ][ 85 ],
   alphaCSR[ 130 ][ 86 ],
   alphaCSR[ 130 ][ 87 ],
   alphaCSR[ 130 ][ 88 ],
   alphaCSR[ 130 ][ 89 ],
   alphaCSR[ 130 ][ 90 ],
   alphaCSR[ 130 ][ 91 ],
   alphaCSR[ 130 ][ 92 ],
   alphaCSR[ 130 ][ 93 ],
   alphaCSR[ 130 ][ 94 ],
   alphaCSR[ 130 ][ 95 ],
   alphaCSR[ 130 ][ 96 ],
   alphaCSR[ 130 ][ 97 ],
   alphaCSR[ 130 ][ 98 ],
   alphaCSR[ 130 ][ 99 ],
   alphaCSR[ 130 ][ 100 ],
   alphaCSR[ 130 ][ 101 ],
   alphaCSR[ 130 ][ 102 ],
   alphaCSR[ 130 ][ 103 ],
   alphaCSR[ 130 ][ 104 ],
   alphaCSR[ 130 ][ 105 ],
   alphaCSR[ 130 ][ 106 ],
   alphaCSR[ 130 ][ 107 ],
   alphaCSR[ 130 ][ 108 ],
   alphaCSR[ 130 ][ 109 ],
   alphaCSR[ 130 ][ 110 ],
   alphaCSR[ 130 ][ 111 ],
   alphaCSR[ 130 ][ 112 ],
   alphaCSR[ 130 ][ 113 ],
   alphaCSR[ 130 ][ 114 ],
   alphaCSR[ 130 ][ 115 ],
   alphaCSR[ 130 ][ 116 ],
   alphaCSR[ 130 ][ 117 ],
   alphaCSR[ 130 ][ 118 ],
   alphaCSR[ 130 ][ 119 ],
   alphaCSR[ 130 ][ 120 ],
   alphaCSR[ 130 ][ 121 ],
   alphaCSR[ 130 ][ 122 ],
   alphaCSR[ 130 ][ 123 ],
   alphaCSR[ 130 ][ 124 ],
   alphaCSR[ 130 ][ 125 ],
   alphaCSR[ 130 ][ 126 ],
   alphaCSR[ 130 ][ 127 ],
   alphaCSR[ 130 ][ 128 ],
   alphaCSR[ 130 ][ 129 ],
   alphaCSR[ 130 ][ 130 ],
   alphaCSR[ 130 ][ 131 ],
   alphaCSR[ 130 ][ 132 ],
   alphaCSR[ 130 ][ 133 ],
   alphaCSR[ 130 ][ 134 ],
   alphaCSR[ 130 ][ 135 ],
   alphaCSR[ 130 ][ 136 ],
   alphaCSR[ 130 ][ 137 ],
   alphaCSR[ 130 ][ 138 ],
   alphaCSR[ 130 ][ 139 ],
   alphaCSR[ 130 ][ 140 ],
   alphaCSR[ 130 ][ 141 ],
   alphaCSR[ 130 ][ 142 ],
   alphaCSR[ 130 ][ 143 ],
   alphaCSR[ 130 ][ 144 ],
   alphaCSR[ 130 ][ 145 ],
   alphaCSR[ 130 ][ 146 ],
   alphaCSR[ 130 ][ 147 ],
   alphaCSR[ 130 ][ 148 ],
   alphaCSR[ 130 ][ 149 ],
   alphaCSR[ 130 ][ 150 ],
   alphaCSR[ 130 ][ 151 ],
   alphaCSR[ 130 ][ 152 ],
   alphaCSR[ 130 ][ 153 ],
   alphaCSR[ 130 ][ 154 ],
   alphaCSR[ 130 ][ 155 ],
   alphaCSR[ 130 ][ 156 ],
   alphaCSR[ 130 ][ 157 ],
   alphaCSR[ 130 ][ 158 ],
   alphaCSR[ 130 ][ 159 ],
   alphaCSR[ 130 ][ 160 ],
   alphaCSR[ 130 ][ 161 ],
   alphaCSR[ 130 ][ 162 ],
   alphaCSR[ 130 ][ 163 ],
   alphaCSR[ 130 ][ 164 ],
   alphaCSR[ 130 ][ 165 ],
   alphaCSR[ 130 ][ 166 ],
   alphaCSR[ 130 ][ 167 ],
   alphaCSR[ 130 ][ 168 ],
   alphaCSR[ 130 ][ 169 ],
   alphaCSR[ 130 ][ 170 ],
   alphaCSR[ 130 ][ 171 ],
   alphaCSR[ 130 ][ 172 ],
   alphaCSR[ 130 ][ 173 ],
   alphaCSR[ 130 ][ 174 ],
   alphaCSR[ 130 ][ 175 ],
   alphaCSR[ 130 ][ 176 ],
   alphaCSR[ 130 ][ 177 ],
   alphaCSR[ 130 ][ 178 ],
   alphaCSR[ 130 ][ 179 ],
   alphaCSR[ 130 ][ 180 ],
   alphaCSR[ 130 ][ 181 ],
   alphaCSR[ 130 ][ 182 ],
   alphaCSR[ 130 ][ 183 ],
   alphaCSR[ 130 ][ 184 ],
   alphaCSR[ 130 ][ 185 ],
   alphaCSR[ 130 ][ 186 ],
   alphaCSR[ 130 ][ 187 ],
   alphaCSR[ 130 ][ 188 ],
   alphaCSR[ 130 ][ 189 ],
   alphaCSR[ 130 ][ 190 ],
   alphaCSR[ 130 ][ 191 ],
   alphaCSR[ 130 ][ 192 ],
   alphaCSR[ 130 ][ 193 ],
   alphaCSR[ 130 ][ 194 ],
   alphaCSR[ 130 ][ 195 ],
   alphaCSR[ 130 ][ 196 ],
   alphaCSR[ 130 ][ 197 ],
   alphaCSR[ 130 ][ 198 ],
   alphaCSR[ 130 ][ 199 ],
   alphaCSR[ 130 ][ 200 ],
   alphaCSR[ 130 ][ 201 ],
   alphaCSR[ 130 ][ 202 ],
   alphaCSR[ 130 ][ 203 ],
   alphaCSR[ 130 ][ 204 ],
   alphaCSR[ 130 ][ 205 ],
   alphaCSR[ 130 ][ 206 ],
   alphaCSR[ 130 ][ 207 ],
   alphaCSR[ 130 ][ 208 ],
   alphaCSR[ 130 ][ 209 ],
   alphaCSR[ 130 ][ 210 ],
   alphaCSR[ 130 ][ 211 ],
   alphaCSR[ 130 ][ 212 ],
   alphaCSR[ 130 ][ 213 ],
   alphaCSR[ 130 ][ 214 ],
   alphaCSR[ 130 ][ 215 ],
   alphaCSR[ 130 ][ 216 ],
   alphaCSR[ 130 ][ 217 ],
   alphaCSR[ 130 ][ 218 ],
   alphaCSR[ 130 ][ 219 ],
   alphaCSR[ 130 ][ 220 ],
   alphaCSR[ 130 ][ 221 ],
   alphaCSR[ 130 ][ 222 ],
   alphaCSR[ 130 ][ 223 ],
   alphaCSR[ 130 ][ 224 ],
   alphaCSR[ 130 ][ 225 ],
   alphaCSR[ 130 ][ 226 ],
   alphaCSR[ 130 ][ 227 ],
   alphaCSR[ 130 ][ 228 ],
   alphaCSR[ 130 ][ 229 ],
   alphaCSR[ 130 ][ 230 ],
   alphaCSR[ 130 ][ 231 ],
   alphaCSR[ 130 ][ 232 ],
   alphaCSR[ 130 ][ 233 ],
   alphaCSR[ 130 ][ 234 ],
   alphaCSR[ 130 ][ 235 ],
   alphaCSR[ 130 ][ 236 ],
   alphaCSR[ 130 ][ 237 ],
   alphaCSR[ 130 ][ 238 ],
   alphaCSR[ 130 ][ 239 ],
   alphaCSR[ 130 ][ 240 ],
   alphaCSR[ 130 ][ 241 ],
   alphaCSR[ 130 ][ 242 ],
   alphaCSR[ 130 ][ 243 ],
   alphaCSR[ 130 ][ 244 ],
   alphaCSR[ 130 ][ 245 ],
   alphaCSR[ 130 ][ 246 ],
   alphaCSR[ 130 ][ 247 ],
   alphaCSR[ 130 ][ 248 ],
   alphaCSR[ 130 ][ 249 ],
   alphaCSR[ 130 ][ 250 ],
   alphaCSR[ 130 ][ 251 ],
   alphaCSR[ 130 ][ 252 ],
   alphaCSR[ 130 ][ 253 ],
   alphaCSR[ 130 ][ 254 ],
   alphaCSR[ 130 ][ 255 ],
   alphaCSR[ 130 ][ 256 ],
   alphaCSR[ 130 ][ 257 ],
   alphaCSR[ 130 ][ 258 ],
   alphaCSR[ 130 ][ 259 ],
   alphaCSR[ 130 ][ 260 ],
   alphaCSR[ 130 ][ 261 ],
   alphaCSR[ 130 ][ 262 ],
   alphaCSR[ 130 ][ 263 ],
   alphaCSR[ 130 ][ 264 ],
   alphaCSR[ 130 ][ 265 ],
   alphaCSR[ 130 ][ 266 ],
   alphaCSR[ 130 ][ 267 ],
   alphaCSR[ 130 ][ 268 ],
   alphaCSR[ 130 ][ 269 ],
   alphaCSR[ 130 ][ 270 ],
   alphaCSR[ 130 ][ 271 ],
   alphaCSR[ 130 ][ 272 ],
   alphaCSR[ 130 ][ 273 ],
   alphaCSR[ 130 ][ 274 ],
   alphaCSR[ 130 ][ 275 ],
   alphaCSR[ 130 ][ 276 ],
   alphaCSR[ 130 ][ 277 ],
   alphaCSR[ 130 ][ 278 ],
   alphaCSR[ 130 ][ 279 ],
   alphaCSR[ 130 ][ 280 ],
   alphaCSR[ 130 ][ 281 ],
   alphaCSR[ 130 ][ 282 ],
   alphaCSR[ 130 ][ 283 ],
   alphaCSR[ 130 ][ 284 ],
   alphaCSR[ 130 ][ 285 ],
   alphaCSR[ 130 ][ 286 ],
   alphaCSR[ 130 ][ 287 ],
   alphaCSR[ 130 ][ 288 ],
   alphaCSR[ 130 ][ 289 ],
   alphaCSR[ 130 ][ 290 ],
   alphaCSR[ 130 ][ 291 ],
   alphaCSR[ 130 ][ 292 ],
   alphaCSR[ 130 ][ 293 ],
   alphaCSR[ 130 ][ 294 ],
   alphaCSR[ 130 ][ 295 ],
   alphaCSR[ 130 ][ 296 ],
   alphaCSR[ 130 ][ 297 ],
   alphaCSR[ 130 ][ 298 ],
   alphaCSR[ 130 ][ 299 ],
   alphaCSR[ 130 ][ 300 ],
   alphaCSR[ 130 ][ 301 ],
   alphaCSR[ 130 ][ 302 ],
   alphaCSR[ 130 ][ 303 ],
   alphaCSR[ 130 ][ 304 ],
   alphaCSR[ 130 ][ 305 ],
   alphaCSR[ 130 ][ 306 ],
   alphaCSR[ 130 ][ 307 ],
   alphaCSR[ 130 ][ 308 ],
   alphaCSR[ 130 ][ 309 ],
   alphaCSR[ 130 ][ 310 ],
   alphaCSR[ 130 ][ 311 ],
   alphaCSR[ 130 ][ 312 ],
   alphaCSR[ 130 ][ 313 ],
   alphaCSR[ 130 ][ 314 ],
   alphaCSR[ 130 ][ 315 ],
   alphaCSR[ 130 ][ 316 ],
   alphaCSR[ 130 ][ 317 ],
   alphaCSR[ 130 ][ 318 ],
   alphaCSR[ 130 ][ 319 ],
   alphaCSR[ 130 ][ 320 ],
   alphaCSR[ 130 ][ 321 ],
   alphaCSR[ 130 ][ 322 ],
   alphaCSR[ 130 ][ 323 ],
   alphaCSR[ 130 ][ 324 ],
   alphaCSR[ 130 ][ 325 ],
   alphaCSR[ 130 ][ 326 ],
   alphaCSR[ 130 ][ 327 ],
   alphaCSR[ 130 ][ 328 ],
   alphaCSR[ 130 ][ 329 ],
   alphaCSR[ 130 ][ 330 ],
   alphaCSR[ 130 ][ 331 ],
   alphaCSR[ 130 ][ 332 ],
   alphaCSR[ 130 ][ 333 ],
   alphaCSR[ 130 ][ 334 ],
   alphaCSR[ 130 ][ 335 ],
   alphaCSR[ 130 ][ 336 ],
   alphaCSR[ 130 ][ 337 ],
   alphaCSR[ 130 ][ 338 ],
   alphaCSR[ 130 ][ 339 ],
   alphaCSR[ 130 ][ 340 ],
   alphaCSR[ 130 ][ 341 ],
   alphaCSR[ 130 ][ 342 ],
   alphaCSR[ 130 ][ 343 ],
   alphaCSR[ 130 ][ 344 ],
   alphaCSR[ 130 ][ 345 ],
   alphaCSR[ 130 ][ 346 ],
   alphaCSR[ 130 ][ 347 ],
   alphaCSR[ 130 ][ 348 ],
   alphaCSR[ 130 ][ 349 ],
   alphaCSR[ 130 ][ 350 ],
   alphaCSR[ 130 ][ 351 ],
   alphaCSR[ 130 ][ 352 ],
   alphaCSR[ 130 ][ 353 ],
   alphaCSR[ 130 ][ 354 ],
   alphaCSR[ 130 ][ 355 ],
   alphaCSR[ 130 ][ 356 ],
   alphaCSR[ 130 ][ 357 ],
   alphaCSR[ 130 ][ 358 ],
   alphaCSR[ 130 ][ 359 ],
   alphaCSR[ 130 ][ 360 ],
   alphaCSR[ 130 ][ 361 ],
   alphaCSR[ 130 ][ 362 ],
   alphaCSR[ 130 ][ 363 ],
   alphaCSR[ 130 ][ 364 ],
   alphaCSR[ 130 ][ 365 ],
   alphaCSR[ 130 ][ 366 ],
   alphaCSR[ 130 ][ 367 ],
   alphaCSR[ 130 ][ 368 ],
   alphaCSR[ 130 ][ 369 ],
   alphaCSR[ 130 ][ 370 ],
   alphaCSR[ 130 ][ 371 ],
   alphaCSR[ 130 ][ 372 ],
   alphaCSR[ 130 ][ 373 ],
   alphaCSR[ 130 ][ 374 ],
   alphaCSR[ 130 ][ 375 ],
   alphaCSR[ 130 ][ 376 ],
   alphaCSR[ 130 ][ 377 ],
   alphaCSR[ 130 ][ 378 ],
   alphaCSR[ 130 ][ 379 ],
   alphaCSR[ 130 ][ 380 ],
   alphaCSR[ 130 ][ 381 ],
   alphaCSR[ 130 ][ 382 ],
   alphaCSR[ 130 ][ 383 ],
   alphaCSR[ 131 ][ 0 ],
   alphaCSR[ 131 ][ 1 ],
   alphaCSR[ 131 ][ 2 ],
   alphaCSR[ 131 ][ 3 ],
   alphaCSR[ 131 ][ 4 ],
   alphaCSR[ 131 ][ 5 ],
   alphaCSR[ 131 ][ 6 ],
   alphaCSR[ 131 ][ 7 ],
   alphaCSR[ 131 ][ 8 ],
   alphaCSR[ 131 ][ 9 ],
   alphaCSR[ 131 ][ 10 ],
   alphaCSR[ 131 ][ 11 ],
   alphaCSR[ 131 ][ 12 ],
   alphaCSR[ 131 ][ 13 ],
   alphaCSR[ 131 ][ 14 ],
   alphaCSR[ 131 ][ 15 ],
   alphaCSR[ 131 ][ 16 ],
   alphaCSR[ 131 ][ 17 ],
   alphaCSR[ 131 ][ 18 ],
   alphaCSR[ 131 ][ 19 ],
   alphaCSR[ 131 ][ 20 ],
   alphaCSR[ 131 ][ 21 ],
   alphaCSR[ 131 ][ 22 ],
   alphaCSR[ 131 ][ 23 ],
   alphaCSR[ 131 ][ 24 ],
   alphaCSR[ 131 ][ 25 ],
   alphaCSR[ 131 ][ 26 ],
   alphaCSR[ 131 ][ 27 ],
   alphaCSR[ 131 ][ 28 ],
   alphaCSR[ 131 ][ 29 ],
   alphaCSR[ 131 ][ 30 ],
   alphaCSR[ 131 ][ 31 ],
   alphaCSR[ 131 ][ 32 ],
   alphaCSR[ 131 ][ 33 ],
   alphaCSR[ 131 ][ 34 ],
   alphaCSR[ 131 ][ 35 ],
   alphaCSR[ 131 ][ 36 ],
   alphaCSR[ 131 ][ 37 ],
   alphaCSR[ 131 ][ 38 ],
   alphaCSR[ 131 ][ 39 ],
   alphaCSR[ 131 ][ 40 ],
   alphaCSR[ 131 ][ 41 ],
   alphaCSR[ 131 ][ 42 ],
   alphaCSR[ 131 ][ 43 ],
   alphaCSR[ 131 ][ 44 ],
   alphaCSR[ 131 ][ 45 ],
   alphaCSR[ 131 ][ 46 ],
   alphaCSR[ 131 ][ 47 ],
   alphaCSR[ 131 ][ 48 ],
   alphaCSR[ 131 ][ 49 ],
   alphaCSR[ 131 ][ 50 ],
   alphaCSR[ 131 ][ 51 ],
   alphaCSR[ 131 ][ 52 ],
   alphaCSR[ 131 ][ 53 ],
   alphaCSR[ 131 ][ 54 ],
   alphaCSR[ 131 ][ 55 ],
   alphaCSR[ 131 ][ 56 ],
   alphaCSR[ 131 ][ 57 ],
   alphaCSR[ 131 ][ 58 ],
   alphaCSR[ 131 ][ 59 ],
   alphaCSR[ 131 ][ 60 ],
   alphaCSR[ 131 ][ 61 ],
   alphaCSR[ 131 ][ 62 ],
   alphaCSR[ 131 ][ 63 ],
   alphaCSR[ 131 ][ 64 ],
   alphaCSR[ 131 ][ 65 ],
   alphaCSR[ 131 ][ 66 ],
   alphaCSR[ 131 ][ 67 ],
   alphaCSR[ 131 ][ 68 ],
   alphaCSR[ 131 ][ 69 ],
   alphaCSR[ 131 ][ 70 ],
   alphaCSR[ 131 ][ 71 ],
   alphaCSR[ 131 ][ 72 ],
   alphaCSR[ 131 ][ 73 ],
   alphaCSR[ 131 ][ 74 ],
   alphaCSR[ 131 ][ 75 ],
   alphaCSR[ 131 ][ 76 ],
   alphaCSR[ 131 ][ 77 ],
   alphaCSR[ 131 ][ 78 ],
   alphaCSR[ 131 ][ 79 ],
   alphaCSR[ 131 ][ 80 ],
   alphaCSR[ 131 ][ 81 ],
   alphaCSR[ 131 ][ 82 ],
   alphaCSR[ 131 ][ 83 ],
   alphaCSR[ 131 ][ 84 ],
   alphaCSR[ 131 ][ 85 ],
   alphaCSR[ 131 ][ 86 ],
   alphaCSR[ 131 ][ 87 ],
   alphaCSR[ 131 ][ 88 ],
   alphaCSR[ 131 ][ 89 ],
   alphaCSR[ 131 ][ 90 ],
   alphaCSR[ 131 ][ 91 ],
   alphaCSR[ 131 ][ 92 ],
   alphaCSR[ 131 ][ 93 ],
   alphaCSR[ 131 ][ 94 ],
   alphaCSR[ 131 ][ 95 ],
   alphaCSR[ 131 ][ 96 ],
   alphaCSR[ 131 ][ 97 ],
   alphaCSR[ 131 ][ 98 ],
   alphaCSR[ 131 ][ 99 ],
   alphaCSR[ 131 ][ 100 ],
   alphaCSR[ 131 ][ 101 ],
   alphaCSR[ 131 ][ 102 ],
   alphaCSR[ 131 ][ 103 ],
   alphaCSR[ 131 ][ 104 ],
   alphaCSR[ 131 ][ 105 ],
   alphaCSR[ 131 ][ 106 ],
   alphaCSR[ 131 ][ 107 ],
   alphaCSR[ 131 ][ 108 ],
   alphaCSR[ 131 ][ 109 ],
   alphaCSR[ 131 ][ 110 ],
   alphaCSR[ 131 ][ 111 ],
   alphaCSR[ 131 ][ 112 ],
   alphaCSR[ 131 ][ 113 ],
   alphaCSR[ 131 ][ 114 ],
   alphaCSR[ 131 ][ 115 ],
   alphaCSR[ 131 ][ 116 ],
   alphaCSR[ 131 ][ 117 ],
   alphaCSR[ 131 ][ 118 ],
   alphaCSR[ 131 ][ 119 ],
   alphaCSR[ 131 ][ 120 ],
   alphaCSR[ 131 ][ 121 ],
   alphaCSR[ 131 ][ 122 ],
   alphaCSR[ 131 ][ 123 ],
   alphaCSR[ 131 ][ 124 ],
   alphaCSR[ 131 ][ 125 ],
   alphaCSR[ 131 ][ 126 ],
   alphaCSR[ 131 ][ 127 ],
   alphaCSR[ 131 ][ 128 ],
   alphaCSR[ 131 ][ 129 ],
   alphaCSR[ 131 ][ 130 ],
   alphaCSR[ 131 ][ 131 ],
   alphaCSR[ 131 ][ 132 ],
   alphaCSR[ 131 ][ 133 ],
   alphaCSR[ 131 ][ 134 ],
   alphaCSR[ 131 ][ 135 ],
   alphaCSR[ 131 ][ 136 ],
   alphaCSR[ 131 ][ 137 ],
   alphaCSR[ 131 ][ 138 ],
   alphaCSR[ 131 ][ 139 ],
   alphaCSR[ 131 ][ 140 ],
   alphaCSR[ 131 ][ 141 ],
   alphaCSR[ 131 ][ 142 ],
   alphaCSR[ 131 ][ 143 ],
   alphaCSR[ 131 ][ 144 ],
   alphaCSR[ 131 ][ 145 ],
   alphaCSR[ 131 ][ 146 ],
   alphaCSR[ 131 ][ 147 ],
   alphaCSR[ 131 ][ 148 ],
   alphaCSR[ 131 ][ 149 ],
   alphaCSR[ 131 ][ 150 ],
   alphaCSR[ 131 ][ 151 ],
   alphaCSR[ 131 ][ 152 ],
   alphaCSR[ 131 ][ 153 ],
   alphaCSR[ 131 ][ 154 ],
   alphaCSR[ 131 ][ 155 ],
   alphaCSR[ 131 ][ 156 ],
   alphaCSR[ 131 ][ 157 ],
   alphaCSR[ 131 ][ 158 ],
   alphaCSR[ 131 ][ 159 ],
   alphaCSR[ 131 ][ 160 ],
   alphaCSR[ 131 ][ 161 ],
   alphaCSR[ 131 ][ 162 ],
   alphaCSR[ 131 ][ 163 ],
   alphaCSR[ 131 ][ 164 ],
   alphaCSR[ 131 ][ 165 ],
   alphaCSR[ 131 ][ 166 ],
   alphaCSR[ 131 ][ 167 ],
   alphaCSR[ 131 ][ 168 ],
   alphaCSR[ 131 ][ 169 ],
   alphaCSR[ 131 ][ 170 ],
   alphaCSR[ 131 ][ 171 ],
   alphaCSR[ 131 ][ 172 ],
   alphaCSR[ 131 ][ 173 ],
   alphaCSR[ 131 ][ 174 ],
   alphaCSR[ 131 ][ 175 ],
   alphaCSR[ 131 ][ 176 ],
   alphaCSR[ 131 ][ 177 ],
   alphaCSR[ 131 ][ 178 ],
   alphaCSR[ 131 ][ 179 ],
   alphaCSR[ 131 ][ 180 ],
   alphaCSR[ 131 ][ 181 ],
   alphaCSR[ 131 ][ 182 ],
   alphaCSR[ 131 ][ 183 ],
   alphaCSR[ 131 ][ 184 ],
   alphaCSR[ 131 ][ 185 ],
   alphaCSR[ 131 ][ 186 ],
   alphaCSR[ 131 ][ 187 ],
   alphaCSR[ 131 ][ 188 ],
   alphaCSR[ 131 ][ 189 ],
   alphaCSR[ 131 ][ 190 ],
   alphaCSR[ 131 ][ 191 ],
   alphaCSR[ 131 ][ 192 ],
   alphaCSR[ 131 ][ 193 ],
   alphaCSR[ 131 ][ 194 ],
   alphaCSR[ 131 ][ 195 ],
   alphaCSR[ 131 ][ 196 ],
   alphaCSR[ 131 ][ 197 ],
   alphaCSR[ 131 ][ 198 ],
   alphaCSR[ 131 ][ 199 ],
   alphaCSR[ 131 ][ 200 ],
   alphaCSR[ 131 ][ 201 ],
   alphaCSR[ 131 ][ 202 ],
   alphaCSR[ 131 ][ 203 ],
   alphaCSR[ 131 ][ 204 ],
   alphaCSR[ 131 ][ 205 ],
   alphaCSR[ 131 ][ 206 ],
   alphaCSR[ 131 ][ 207 ],
   alphaCSR[ 131 ][ 208 ],
   alphaCSR[ 131 ][ 209 ],
   alphaCSR[ 131 ][ 210 ],
   alphaCSR[ 131 ][ 211 ],
   alphaCSR[ 131 ][ 212 ],
   alphaCSR[ 131 ][ 213 ],
   alphaCSR[ 131 ][ 214 ],
   alphaCSR[ 131 ][ 215 ],
   alphaCSR[ 131 ][ 216 ],
   alphaCSR[ 131 ][ 217 ],
   alphaCSR[ 131 ][ 218 ],
   alphaCSR[ 131 ][ 219 ],
   alphaCSR[ 131 ][ 220 ],
   alphaCSR[ 131 ][ 221 ],
   alphaCSR[ 131 ][ 222 ],
   alphaCSR[ 131 ][ 223 ],
   alphaCSR[ 131 ][ 224 ],
   alphaCSR[ 131 ][ 225 ],
   alphaCSR[ 131 ][ 226 ],
   alphaCSR[ 131 ][ 227 ],
   alphaCSR[ 131 ][ 228 ],
   alphaCSR[ 131 ][ 229 ],
   alphaCSR[ 131 ][ 230 ],
   alphaCSR[ 131 ][ 231 ],
   alphaCSR[ 131 ][ 232 ],
   alphaCSR[ 131 ][ 233 ],
   alphaCSR[ 131 ][ 234 ],
   alphaCSR[ 131 ][ 235 ],
   alphaCSR[ 131 ][ 236 ],
   alphaCSR[ 131 ][ 237 ],
   alphaCSR[ 131 ][ 238 ],
   alphaCSR[ 131 ][ 239 ],
   alphaCSR[ 131 ][ 240 ],
   alphaCSR[ 131 ][ 241 ],
   alphaCSR[ 131 ][ 242 ],
   alphaCSR[ 131 ][ 243 ],
   alphaCSR[ 131 ][ 244 ],
   alphaCSR[ 131 ][ 245 ],
   alphaCSR[ 131 ][ 246 ],
   alphaCSR[ 131 ][ 247 ],
   alphaCSR[ 131 ][ 248 ],
   alphaCSR[ 131 ][ 249 ],
   alphaCSR[ 131 ][ 250 ],
   alphaCSR[ 131 ][ 251 ],
   alphaCSR[ 131 ][ 252 ],
   alphaCSR[ 131 ][ 253 ],
   alphaCSR[ 131 ][ 254 ],
   alphaCSR[ 131 ][ 255 ],
   alphaCSR[ 131 ][ 256 ],
   alphaCSR[ 131 ][ 257 ],
   alphaCSR[ 131 ][ 258 ],
   alphaCSR[ 131 ][ 259 ],
   alphaCSR[ 131 ][ 260 ],
   alphaCSR[ 131 ][ 261 ],
   alphaCSR[ 131 ][ 262 ],
   alphaCSR[ 131 ][ 263 ],
   alphaCSR[ 131 ][ 264 ],
   alphaCSR[ 131 ][ 265 ],
   alphaCSR[ 131 ][ 266 ],
   alphaCSR[ 131 ][ 267 ],
   alphaCSR[ 131 ][ 268 ],
   alphaCSR[ 131 ][ 269 ],
   alphaCSR[ 131 ][ 270 ],
   alphaCSR[ 131 ][ 271 ],
   alphaCSR[ 131 ][ 272 ],
   alphaCSR[ 131 ][ 273 ],
   alphaCSR[ 131 ][ 274 ],
   alphaCSR[ 131 ][ 275 ],
   alphaCSR[ 131 ][ 276 ],
   alphaCSR[ 131 ][ 277 ],
   alphaCSR[ 131 ][ 278 ],
   alphaCSR[ 131 ][ 279 ],
   alphaCSR[ 131 ][ 280 ],
   alphaCSR[ 131 ][ 281 ],
   alphaCSR[ 131 ][ 282 ],
   alphaCSR[ 131 ][ 283 ],
   alphaCSR[ 131 ][ 284 ],
   alphaCSR[ 131 ][ 285 ],
   alphaCSR[ 131 ][ 286 ],
   alphaCSR[ 131 ][ 287 ],
   alphaCSR[ 131 ][ 288 ],
   alphaCSR[ 131 ][ 289 ],
   alphaCSR[ 131 ][ 290 ],
   alphaCSR[ 131 ][ 291 ],
   alphaCSR[ 131 ][ 292 ],
   alphaCSR[ 131 ][ 293 ],
   alphaCSR[ 131 ][ 294 ],
   alphaCSR[ 131 ][ 295 ],
   alphaCSR[ 131 ][ 296 ],
   alphaCSR[ 131 ][ 297 ],
   alphaCSR[ 131 ][ 298 ],
   alphaCSR[ 131 ][ 299 ],
   alphaCSR[ 131 ][ 300 ],
   alphaCSR[ 131 ][ 301 ],
   alphaCSR[ 131 ][ 302 ],
   alphaCSR[ 131 ][ 303 ],
   alphaCSR[ 131 ][ 304 ],
   alphaCSR[ 131 ][ 305 ],
   alphaCSR[ 131 ][ 306 ],
   alphaCSR[ 131 ][ 307 ],
   alphaCSR[ 131 ][ 308 ],
   alphaCSR[ 131 ][ 309 ],
   alphaCSR[ 131 ][ 310 ],
   alphaCSR[ 131 ][ 311 ],
   alphaCSR[ 131 ][ 312 ],
   alphaCSR[ 131 ][ 313 ],
   alphaCSR[ 131 ][ 314 ],
   alphaCSR[ 131 ][ 315 ],
   alphaCSR[ 131 ][ 316 ],
   alphaCSR[ 131 ][ 317 ],
   alphaCSR[ 131 ][ 318 ],
   alphaCSR[ 131 ][ 319 ],
   alphaCSR[ 131 ][ 320 ],
   alphaCSR[ 131 ][ 321 ],
   alphaCSR[ 131 ][ 322 ],
   alphaCSR[ 131 ][ 323 ],
   alphaCSR[ 131 ][ 324 ],
   alphaCSR[ 131 ][ 325 ],
   alphaCSR[ 131 ][ 326 ],
   alphaCSR[ 131 ][ 327 ],
   alphaCSR[ 131 ][ 328 ],
   alphaCSR[ 131 ][ 329 ],
   alphaCSR[ 131 ][ 330 ],
   alphaCSR[ 131 ][ 331 ],
   alphaCSR[ 131 ][ 332 ],
   alphaCSR[ 131 ][ 333 ],
   alphaCSR[ 131 ][ 334 ],
   alphaCSR[ 131 ][ 335 ],
   alphaCSR[ 131 ][ 336 ],
   alphaCSR[ 131 ][ 337 ],
   alphaCSR[ 131 ][ 338 ],
   alphaCSR[ 131 ][ 339 ],
   alphaCSR[ 131 ][ 340 ],
   alphaCSR[ 131 ][ 341 ],
   alphaCSR[ 131 ][ 342 ],
   alphaCSR[ 131 ][ 343 ],
   alphaCSR[ 131 ][ 344 ],
   alphaCSR[ 131 ][ 345 ],
   alphaCSR[ 131 ][ 346 ],
   alphaCSR[ 131 ][ 347 ],
   alphaCSR[ 131 ][ 348 ],
   alphaCSR[ 131 ][ 349 ],
   alphaCSR[ 131 ][ 350 ],
   alphaCSR[ 131 ][ 351 ],
   alphaCSR[ 131 ][ 352 ],
   alphaCSR[ 131 ][ 353 ],
   alphaCSR[ 131 ][ 354 ],
   alphaCSR[ 131 ][ 355 ],
   alphaCSR[ 131 ][ 356 ],
   alphaCSR[ 131 ][ 357 ],
   alphaCSR[ 131 ][ 358 ],
   alphaCSR[ 131 ][ 359 ],
   alphaCSR[ 131 ][ 360 ],
   alphaCSR[ 131 ][ 361 ],
   alphaCSR[ 131 ][ 362 ],
   alphaCSR[ 131 ][ 363 ],
   alphaCSR[ 131 ][ 364 ],
   alphaCSR[ 131 ][ 365 ],
   alphaCSR[ 131 ][ 366 ],
   alphaCSR[ 131 ][ 367 ],
   alphaCSR[ 131 ][ 368 ],
   alphaCSR[ 131 ][ 369 ],
   alphaCSR[ 131 ][ 370 ],
   alphaCSR[ 131 ][ 371 ],
   alphaCSR[ 131 ][ 372 ],
   alphaCSR[ 131 ][ 373 ],
   alphaCSR[ 131 ][ 374 ],
   alphaCSR[ 131 ][ 375 ],
   alphaCSR[ 131 ][ 376 ],
   alphaCSR[ 131 ][ 377 ],
   alphaCSR[ 131 ][ 378 ],
   alphaCSR[ 131 ][ 379 ],
   alphaCSR[ 131 ][ 380 ],
   alphaCSR[ 131 ][ 381 ],
   alphaCSR[ 131 ][ 382 ],
   alphaCSR[ 131 ][ 383 ],
   alphaCSR[ 132 ][ 0 ],
   alphaCSR[ 132 ][ 1 ],
   alphaCSR[ 132 ][ 2 ],
   alphaCSR[ 132 ][ 3 ],
   alphaCSR[ 132 ][ 4 ],
   alphaCSR[ 132 ][ 5 ],
   alphaCSR[ 132 ][ 6 ],
   alphaCSR[ 132 ][ 7 ],
   alphaCSR[ 132 ][ 8 ],
   alphaCSR[ 132 ][ 9 ],
   alphaCSR[ 132 ][ 10 ],
   alphaCSR[ 132 ][ 11 ],
   alphaCSR[ 132 ][ 12 ],
   alphaCSR[ 132 ][ 13 ],
   alphaCSR[ 132 ][ 14 ],
   alphaCSR[ 132 ][ 15 ],
   alphaCSR[ 132 ][ 16 ],
   alphaCSR[ 132 ][ 17 ],
   alphaCSR[ 132 ][ 18 ],
   alphaCSR[ 132 ][ 19 ],
   alphaCSR[ 132 ][ 20 ],
   alphaCSR[ 132 ][ 21 ],
   alphaCSR[ 132 ][ 22 ],
   alphaCSR[ 132 ][ 23 ],
   alphaCSR[ 132 ][ 24 ],
   alphaCSR[ 132 ][ 25 ],
   alphaCSR[ 132 ][ 26 ],
   alphaCSR[ 132 ][ 27 ],
   alphaCSR[ 132 ][ 28 ],
   alphaCSR[ 132 ][ 29 ],
   alphaCSR[ 132 ][ 30 ],
   alphaCSR[ 132 ][ 31 ],
   alphaCSR[ 132 ][ 32 ],
   alphaCSR[ 132 ][ 33 ],
   alphaCSR[ 132 ][ 34 ],
   alphaCSR[ 132 ][ 35 ],
   alphaCSR[ 132 ][ 36 ],
   alphaCSR[ 132 ][ 37 ],
   alphaCSR[ 132 ][ 38 ],
   alphaCSR[ 132 ][ 39 ],
   alphaCSR[ 132 ][ 40 ],
   alphaCSR[ 132 ][ 41 ],
   alphaCSR[ 132 ][ 42 ],
   alphaCSR[ 132 ][ 43 ],
   alphaCSR[ 132 ][ 44 ],
   alphaCSR[ 132 ][ 45 ],
   alphaCSR[ 132 ][ 46 ],
   alphaCSR[ 132 ][ 47 ],
   alphaCSR[ 132 ][ 48 ],
   alphaCSR[ 132 ][ 49 ],
   alphaCSR[ 132 ][ 50 ],
   alphaCSR[ 132 ][ 51 ],
   alphaCSR[ 132 ][ 52 ],
   alphaCSR[ 132 ][ 53 ],
   alphaCSR[ 132 ][ 54 ],
   alphaCSR[ 132 ][ 55 ],
   alphaCSR[ 132 ][ 56 ],
   alphaCSR[ 132 ][ 57 ],
   alphaCSR[ 132 ][ 58 ],
   alphaCSR[ 132 ][ 59 ],
   alphaCSR[ 132 ][ 60 ],
   alphaCSR[ 132 ][ 61 ],
   alphaCSR[ 132 ][ 62 ],
   alphaCSR[ 132 ][ 63 ],
   alphaCSR[ 132 ][ 64 ],
   alphaCSR[ 132 ][ 65 ],
   alphaCSR[ 132 ][ 66 ],
   alphaCSR[ 132 ][ 67 ],
   alphaCSR[ 132 ][ 68 ],
   alphaCSR[ 132 ][ 69 ],
   alphaCSR[ 132 ][ 70 ],
   alphaCSR[ 132 ][ 71 ],
   alphaCSR[ 132 ][ 72 ],
   alphaCSR[ 132 ][ 73 ],
   alphaCSR[ 132 ][ 74 ],
   alphaCSR[ 132 ][ 75 ],
   alphaCSR[ 132 ][ 76 ],
   alphaCSR[ 132 ][ 77 ],
   alphaCSR[ 132 ][ 78 ],
   alphaCSR[ 132 ][ 79 ],
   alphaCSR[ 132 ][ 80 ],
   alphaCSR[ 132 ][ 81 ],
   alphaCSR[ 132 ][ 82 ],
   alphaCSR[ 132 ][ 83 ],
   alphaCSR[ 132 ][ 84 ],
   alphaCSR[ 132 ][ 85 ],
   alphaCSR[ 132 ][ 86 ],
   alphaCSR[ 132 ][ 87 ],
   alphaCSR[ 132 ][ 88 ],
   alphaCSR[ 132 ][ 89 ],
   alphaCSR[ 132 ][ 90 ],
   alphaCSR[ 132 ][ 91 ],
   alphaCSR[ 132 ][ 92 ],
   alphaCSR[ 132 ][ 93 ],
   alphaCSR[ 132 ][ 94 ],
   alphaCSR[ 132 ][ 95 ],
   alphaCSR[ 132 ][ 96 ],
   alphaCSR[ 132 ][ 97 ],
   alphaCSR[ 132 ][ 98 ],
   alphaCSR[ 132 ][ 99 ],
   alphaCSR[ 132 ][ 100 ],
   alphaCSR[ 132 ][ 101 ],
   alphaCSR[ 132 ][ 102 ],
   alphaCSR[ 132 ][ 103 ],
   alphaCSR[ 132 ][ 104 ],
   alphaCSR[ 132 ][ 105 ],
   alphaCSR[ 132 ][ 106 ],
   alphaCSR[ 132 ][ 107 ],
   alphaCSR[ 132 ][ 108 ],
   alphaCSR[ 132 ][ 109 ],
   alphaCSR[ 132 ][ 110 ],
   alphaCSR[ 132 ][ 111 ],
   alphaCSR[ 132 ][ 112 ],
   alphaCSR[ 132 ][ 113 ],
   alphaCSR[ 132 ][ 114 ],
   alphaCSR[ 132 ][ 115 ],
   alphaCSR[ 132 ][ 116 ],
   alphaCSR[ 132 ][ 117 ],
   alphaCSR[ 132 ][ 118 ],
   alphaCSR[ 132 ][ 119 ],
   alphaCSR[ 132 ][ 120 ],
   alphaCSR[ 132 ][ 121 ],
   alphaCSR[ 132 ][ 122 ],
   alphaCSR[ 132 ][ 123 ],
   alphaCSR[ 132 ][ 124 ],
   alphaCSR[ 132 ][ 125 ],
   alphaCSR[ 132 ][ 126 ],
   alphaCSR[ 132 ][ 127 ],
   alphaCSR[ 132 ][ 128 ],
   alphaCSR[ 132 ][ 129 ],
   alphaCSR[ 132 ][ 130 ],
   alphaCSR[ 132 ][ 131 ],
   alphaCSR[ 132 ][ 132 ],
   alphaCSR[ 132 ][ 133 ],
   alphaCSR[ 132 ][ 134 ],
   alphaCSR[ 132 ][ 135 ],
   alphaCSR[ 132 ][ 136 ],
   alphaCSR[ 132 ][ 137 ],
   alphaCSR[ 132 ][ 138 ],
   alphaCSR[ 132 ][ 139 ],
   alphaCSR[ 132 ][ 140 ],
   alphaCSR[ 132 ][ 141 ],
   alphaCSR[ 132 ][ 142 ],
   alphaCSR[ 132 ][ 143 ],
   alphaCSR[ 132 ][ 144 ],
   alphaCSR[ 132 ][ 145 ],
   alphaCSR[ 132 ][ 146 ],
   alphaCSR[ 132 ][ 147 ],
   alphaCSR[ 132 ][ 148 ],
   alphaCSR[ 132 ][ 149 ],
   alphaCSR[ 132 ][ 150 ],
   alphaCSR[ 132 ][ 151 ],
   alphaCSR[ 132 ][ 152 ],
   alphaCSR[ 132 ][ 153 ],
   alphaCSR[ 132 ][ 154 ],
   alphaCSR[ 132 ][ 155 ],
   alphaCSR[ 132 ][ 156 ],
   alphaCSR[ 132 ][ 157 ],
   alphaCSR[ 132 ][ 158 ],
   alphaCSR[ 132 ][ 159 ],
   alphaCSR[ 132 ][ 160 ],
   alphaCSR[ 132 ][ 161 ],
   alphaCSR[ 132 ][ 162 ],
   alphaCSR[ 132 ][ 163 ],
   alphaCSR[ 132 ][ 164 ],
   alphaCSR[ 132 ][ 165 ],
   alphaCSR[ 132 ][ 166 ],
   alphaCSR[ 132 ][ 167 ],
   alphaCSR[ 132 ][ 168 ],
   alphaCSR[ 132 ][ 169 ],
   alphaCSR[ 132 ][ 170 ],
   alphaCSR[ 132 ][ 171 ],
   alphaCSR[ 132 ][ 172 ],
   alphaCSR[ 132 ][ 173 ],
   alphaCSR[ 132 ][ 174 ],
   alphaCSR[ 132 ][ 175 ],
   alphaCSR[ 132 ][ 176 ],
   alphaCSR[ 132 ][ 177 ],
   alphaCSR[ 132 ][ 178 ],
   alphaCSR[ 132 ][ 179 ],
   alphaCSR[ 132 ][ 180 ],
   alphaCSR[ 132 ][ 181 ],
   alphaCSR[ 132 ][ 182 ],
   alphaCSR[ 132 ][ 183 ],
   alphaCSR[ 132 ][ 184 ],
   alphaCSR[ 132 ][ 185 ],
   alphaCSR[ 132 ][ 186 ],
   alphaCSR[ 132 ][ 187 ],
   alphaCSR[ 132 ][ 188 ],
   alphaCSR[ 132 ][ 189 ],
   alphaCSR[ 132 ][ 190 ],
   alphaCSR[ 132 ][ 191 ],
   alphaCSR[ 132 ][ 192 ],
   alphaCSR[ 132 ][ 193 ],
   alphaCSR[ 132 ][ 194 ],
   alphaCSR[ 132 ][ 195 ],
   alphaCSR[ 132 ][ 196 ],
   alphaCSR[ 132 ][ 197 ],
   alphaCSR[ 132 ][ 198 ],
   alphaCSR[ 132 ][ 199 ],
   alphaCSR[ 132 ][ 200 ],
   alphaCSR[ 132 ][ 201 ],
   alphaCSR[ 132 ][ 202 ],
   alphaCSR[ 132 ][ 203 ],
   alphaCSR[ 132 ][ 204 ],
   alphaCSR[ 132 ][ 205 ],
   alphaCSR[ 132 ][ 206 ],
   alphaCSR[ 132 ][ 207 ],
   alphaCSR[ 132 ][ 208 ],
   alphaCSR[ 132 ][ 209 ],
   alphaCSR[ 132 ][ 210 ],
   alphaCSR[ 132 ][ 211 ],
   alphaCSR[ 132 ][ 212 ],
   alphaCSR[ 132 ][ 213 ],
   alphaCSR[ 132 ][ 214 ],
   alphaCSR[ 132 ][ 215 ],
   alphaCSR[ 132 ][ 216 ],
   alphaCSR[ 132 ][ 217 ],
   alphaCSR[ 132 ][ 218 ],
   alphaCSR[ 132 ][ 219 ],
   alphaCSR[ 132 ][ 220 ],
   alphaCSR[ 132 ][ 221 ],
   alphaCSR[ 132 ][ 222 ],
   alphaCSR[ 132 ][ 223 ],
   alphaCSR[ 132 ][ 224 ],
   alphaCSR[ 132 ][ 225 ],
   alphaCSR[ 132 ][ 226 ],
   alphaCSR[ 132 ][ 227 ],
   alphaCSR[ 132 ][ 228 ],
   alphaCSR[ 132 ][ 229 ],
   alphaCSR[ 132 ][ 230 ],
   alphaCSR[ 132 ][ 231 ],
   alphaCSR[ 132 ][ 232 ],
   alphaCSR[ 132 ][ 233 ],
   alphaCSR[ 132 ][ 234 ],
   alphaCSR[ 132 ][ 235 ],
   alphaCSR[ 132 ][ 236 ],
   alphaCSR[ 132 ][ 237 ],
   alphaCSR[ 132 ][ 238 ],
   alphaCSR[ 132 ][ 239 ],
   alphaCSR[ 132 ][ 240 ],
   alphaCSR[ 132 ][ 241 ],
   alphaCSR[ 132 ][ 242 ],
   alphaCSR[ 132 ][ 243 ],
   alphaCSR[ 132 ][ 244 ],
   alphaCSR[ 132 ][ 245 ],
   alphaCSR[ 132 ][ 246 ],
   alphaCSR[ 132 ][ 247 ],
   alphaCSR[ 132 ][ 248 ],
   alphaCSR[ 132 ][ 249 ],
   alphaCSR[ 132 ][ 250 ],
   alphaCSR[ 132 ][ 251 ],
   alphaCSR[ 132 ][ 252 ],
   alphaCSR[ 132 ][ 253 ],
   alphaCSR[ 132 ][ 254 ],
   alphaCSR[ 132 ][ 255 ],
   alphaCSR[ 132 ][ 256 ],
   alphaCSR[ 132 ][ 257 ],
   alphaCSR[ 132 ][ 258 ],
   alphaCSR[ 132 ][ 259 ],
   alphaCSR[ 132 ][ 260 ],
   alphaCSR[ 132 ][ 261 ],
   alphaCSR[ 132 ][ 262 ],
   alphaCSR[ 132 ][ 263 ],
   alphaCSR[ 132 ][ 264 ],
   alphaCSR[ 132 ][ 265 ],
   alphaCSR[ 132 ][ 266 ],
   alphaCSR[ 132 ][ 267 ],
   alphaCSR[ 132 ][ 268 ],
   alphaCSR[ 132 ][ 269 ],
   alphaCSR[ 132 ][ 270 ],
   alphaCSR[ 132 ][ 271 ],
   alphaCSR[ 132 ][ 272 ],
   alphaCSR[ 132 ][ 273 ],
   alphaCSR[ 132 ][ 274 ],
   alphaCSR[ 132 ][ 275 ],
   alphaCSR[ 132 ][ 276 ],
   alphaCSR[ 132 ][ 277 ],
   alphaCSR[ 132 ][ 278 ],
   alphaCSR[ 132 ][ 279 ],
   alphaCSR[ 132 ][ 280 ],
   alphaCSR[ 132 ][ 281 ],
   alphaCSR[ 132 ][ 282 ],
   alphaCSR[ 132 ][ 283 ],
   alphaCSR[ 132 ][ 284 ],
   alphaCSR[ 132 ][ 285 ],
   alphaCSR[ 132 ][ 286 ],
   alphaCSR[ 132 ][ 287 ],
   alphaCSR[ 132 ][ 288 ],
   alphaCSR[ 132 ][ 289 ],
   alphaCSR[ 132 ][ 290 ],
   alphaCSR[ 132 ][ 291 ],
   alphaCSR[ 132 ][ 292 ],
   alphaCSR[ 132 ][ 293 ],
   alphaCSR[ 132 ][ 294 ],
   alphaCSR[ 132 ][ 295 ],
   alphaCSR[ 132 ][ 296 ],
   alphaCSR[ 132 ][ 297 ],
   alphaCSR[ 132 ][ 298 ],
   alphaCSR[ 132 ][ 299 ],
   alphaCSR[ 132 ][ 300 ],
   alphaCSR[ 132 ][ 301 ],
   alphaCSR[ 132 ][ 302 ],
   alphaCSR[ 132 ][ 303 ],
   alphaCSR[ 132 ][ 304 ],
   alphaCSR[ 132 ][ 305 ],
   alphaCSR[ 132 ][ 306 ],
   alphaCSR[ 132 ][ 307 ],
   alphaCSR[ 132 ][ 308 ],
   alphaCSR[ 132 ][ 309 ],
   alphaCSR[ 132 ][ 310 ],
   alphaCSR[ 132 ][ 311 ],
   alphaCSR[ 132 ][ 312 ],
   alphaCSR[ 132 ][ 313 ],
   alphaCSR[ 132 ][ 314 ],
   alphaCSR[ 132 ][ 315 ],
   alphaCSR[ 132 ][ 316 ],
   alphaCSR[ 132 ][ 317 ],
   alphaCSR[ 132 ][ 318 ],
   alphaCSR[ 132 ][ 319 ],
   alphaCSR[ 132 ][ 320 ],
   alphaCSR[ 132 ][ 321 ],
   alphaCSR[ 132 ][ 322 ],
   alphaCSR[ 132 ][ 323 ],
   alphaCSR[ 132 ][ 324 ],
   alphaCSR[ 132 ][ 325 ],
   alphaCSR[ 132 ][ 326 ],
   alphaCSR[ 132 ][ 327 ],
   alphaCSR[ 132 ][ 328 ],
   alphaCSR[ 132 ][ 329 ],
   alphaCSR[ 132 ][ 330 ],
   alphaCSR[ 132 ][ 331 ],
   alphaCSR[ 132 ][ 332 ],
   alphaCSR[ 132 ][ 333 ],
   alphaCSR[ 132 ][ 334 ],
   alphaCSR[ 132 ][ 335 ],
   alphaCSR[ 132 ][ 336 ],
   alphaCSR[ 132 ][ 337 ],
   alphaCSR[ 132 ][ 338 ],
   alphaCSR[ 132 ][ 339 ],
   alphaCSR[ 132 ][ 340 ],
   alphaCSR[ 132 ][ 341 ],
   alphaCSR[ 132 ][ 342 ],
   alphaCSR[ 132 ][ 343 ],
   alphaCSR[ 132 ][ 344 ],
   alphaCSR[ 132 ][ 345 ],
   alphaCSR[ 132 ][ 346 ],
   alphaCSR[ 132 ][ 347 ],
   alphaCSR[ 132 ][ 348 ],
   alphaCSR[ 132 ][ 349 ],
   alphaCSR[ 132 ][ 350 ],
   alphaCSR[ 132 ][ 351 ],
   alphaCSR[ 132 ][ 352 ],
   alphaCSR[ 132 ][ 353 ],
   alphaCSR[ 132 ][ 354 ],
   alphaCSR[ 132 ][ 355 ],
   alphaCSR[ 132 ][ 356 ],
   alphaCSR[ 132 ][ 357 ],
   alphaCSR[ 132 ][ 358 ],
   alphaCSR[ 132 ][ 359 ],
   alphaCSR[ 132 ][ 360 ],
   alphaCSR[ 132 ][ 361 ],
   alphaCSR[ 132 ][ 362 ],
   alphaCSR[ 132 ][ 363 ],
   alphaCSR[ 132 ][ 364 ],
   alphaCSR[ 132 ][ 365 ],
   alphaCSR[ 132 ][ 366 ],
   alphaCSR[ 132 ][ 367 ],
   alphaCSR[ 132 ][ 368 ],
   alphaCSR[ 132 ][ 369 ],
   alphaCSR[ 132 ][ 370 ],
   alphaCSR[ 132 ][ 371 ],
   alphaCSR[ 132 ][ 372 ],
   alphaCSR[ 132 ][ 373 ],
   alphaCSR[ 132 ][ 374 ],
   alphaCSR[ 132 ][ 375 ],
   alphaCSR[ 132 ][ 376 ],
   alphaCSR[ 132 ][ 377 ],
   alphaCSR[ 132 ][ 378 ],
   alphaCSR[ 132 ][ 379 ],
   alphaCSR[ 132 ][ 380 ],
   alphaCSR[ 132 ][ 381 ],
   alphaCSR[ 132 ][ 382 ],
   alphaCSR[ 132 ][ 383 ],
   alphaCSR[ 133 ][ 0 ],
   alphaCSR[ 133 ][ 1 ],
   alphaCSR[ 133 ][ 2 ],
   alphaCSR[ 133 ][ 3 ],
   alphaCSR[ 133 ][ 4 ],
   alphaCSR[ 133 ][ 5 ],
   alphaCSR[ 133 ][ 6 ],
   alphaCSR[ 133 ][ 7 ],
   alphaCSR[ 133 ][ 8 ],
   alphaCSR[ 133 ][ 9 ],
   alphaCSR[ 133 ][ 10 ],
   alphaCSR[ 133 ][ 11 ],
   alphaCSR[ 133 ][ 12 ],
   alphaCSR[ 133 ][ 13 ],
   alphaCSR[ 133 ][ 14 ],
   alphaCSR[ 133 ][ 15 ],
   alphaCSR[ 133 ][ 16 ],
   alphaCSR[ 133 ][ 17 ],
   alphaCSR[ 133 ][ 18 ],
   alphaCSR[ 133 ][ 19 ],
   alphaCSR[ 133 ][ 20 ],
   alphaCSR[ 133 ][ 21 ],
   alphaCSR[ 133 ][ 22 ],
   alphaCSR[ 133 ][ 23 ],
   alphaCSR[ 133 ][ 24 ],
   alphaCSR[ 133 ][ 25 ],
   alphaCSR[ 133 ][ 26 ],
   alphaCSR[ 133 ][ 27 ],
   alphaCSR[ 133 ][ 28 ],
   alphaCSR[ 133 ][ 29 ],
   alphaCSR[ 133 ][ 30 ],
   alphaCSR[ 133 ][ 31 ],
   alphaCSR[ 133 ][ 32 ],
   alphaCSR[ 133 ][ 33 ],
   alphaCSR[ 133 ][ 34 ],
   alphaCSR[ 133 ][ 35 ],
   alphaCSR[ 133 ][ 36 ],
   alphaCSR[ 133 ][ 37 ],
   alphaCSR[ 133 ][ 38 ],
   alphaCSR[ 133 ][ 39 ],
   alphaCSR[ 133 ][ 40 ],
   alphaCSR[ 133 ][ 41 ],
   alphaCSR[ 133 ][ 42 ],
   alphaCSR[ 133 ][ 43 ],
   alphaCSR[ 133 ][ 44 ],
   alphaCSR[ 133 ][ 45 ],
   alphaCSR[ 133 ][ 46 ],
   alphaCSR[ 133 ][ 47 ],
   alphaCSR[ 133 ][ 48 ],
   alphaCSR[ 133 ][ 49 ],
   alphaCSR[ 133 ][ 50 ],
   alphaCSR[ 133 ][ 51 ],
   alphaCSR[ 133 ][ 52 ],
   alphaCSR[ 133 ][ 53 ],
   alphaCSR[ 133 ][ 54 ],
   alphaCSR[ 133 ][ 55 ],
   alphaCSR[ 133 ][ 56 ],
   alphaCSR[ 133 ][ 57 ],
   alphaCSR[ 133 ][ 58 ],
   alphaCSR[ 133 ][ 59 ],
   alphaCSR[ 133 ][ 60 ],
   alphaCSR[ 133 ][ 61 ],
   alphaCSR[ 133 ][ 62 ],
   alphaCSR[ 133 ][ 63 ],
   alphaCSR[ 133 ][ 64 ],
   alphaCSR[ 133 ][ 65 ],
   alphaCSR[ 133 ][ 66 ],
   alphaCSR[ 133 ][ 67 ],
   alphaCSR[ 133 ][ 68 ],
   alphaCSR[ 133 ][ 69 ],
   alphaCSR[ 133 ][ 70 ],
   alphaCSR[ 133 ][ 71 ],
   alphaCSR[ 133 ][ 72 ],
   alphaCSR[ 133 ][ 73 ],
   alphaCSR[ 133 ][ 74 ],
   alphaCSR[ 133 ][ 75 ],
   alphaCSR[ 133 ][ 76 ],
   alphaCSR[ 133 ][ 77 ],
   alphaCSR[ 133 ][ 78 ],
   alphaCSR[ 133 ][ 79 ],
   alphaCSR[ 133 ][ 80 ],
   alphaCSR[ 133 ][ 81 ],
   alphaCSR[ 133 ][ 82 ],
   alphaCSR[ 133 ][ 83 ],
   alphaCSR[ 133 ][ 84 ],
   alphaCSR[ 133 ][ 85 ],
   alphaCSR[ 133 ][ 86 ],
   alphaCSR[ 133 ][ 87 ],
   alphaCSR[ 133 ][ 88 ],
   alphaCSR[ 133 ][ 89 ],
   alphaCSR[ 133 ][ 90 ],
   alphaCSR[ 133 ][ 91 ],
   alphaCSR[ 133 ][ 92 ],
   alphaCSR[ 133 ][ 93 ],
   alphaCSR[ 133 ][ 94 ],
   alphaCSR[ 133 ][ 95 ],
   alphaCSR[ 133 ][ 96 ],
   alphaCSR[ 133 ][ 97 ],
   alphaCSR[ 133 ][ 98 ],
   alphaCSR[ 133 ][ 99 ],
   alphaCSR[ 133 ][ 100 ],
   alphaCSR[ 133 ][ 101 ],
   alphaCSR[ 133 ][ 102 ],
   alphaCSR[ 133 ][ 103 ],
   alphaCSR[ 133 ][ 104 ],
   alphaCSR[ 133 ][ 105 ],
   alphaCSR[ 133 ][ 106 ],
   alphaCSR[ 133 ][ 107 ],
   alphaCSR[ 133 ][ 108 ],
   alphaCSR[ 133 ][ 109 ],
   alphaCSR[ 133 ][ 110 ],
   alphaCSR[ 133 ][ 111 ],
   alphaCSR[ 133 ][ 112 ],
   alphaCSR[ 133 ][ 113 ],
   alphaCSR[ 133 ][ 114 ],
   alphaCSR[ 133 ][ 115 ],
   alphaCSR[ 133 ][ 116 ],
   alphaCSR[ 133 ][ 117 ],
   alphaCSR[ 133 ][ 118 ],
   alphaCSR[ 133 ][ 119 ],
   alphaCSR[ 133 ][ 120 ],
   alphaCSR[ 133 ][ 121 ],
   alphaCSR[ 133 ][ 122 ],
   alphaCSR[ 133 ][ 123 ],
   alphaCSR[ 133 ][ 124 ],
   alphaCSR[ 133 ][ 125 ],
   alphaCSR[ 133 ][ 126 ],
   alphaCSR[ 133 ][ 127 ],
   alphaCSR[ 133 ][ 128 ],
   alphaCSR[ 133 ][ 129 ],
   alphaCSR[ 133 ][ 130 ],
   alphaCSR[ 133 ][ 131 ],
   alphaCSR[ 133 ][ 132 ],
   alphaCSR[ 133 ][ 133 ],
   alphaCSR[ 133 ][ 134 ],
   alphaCSR[ 133 ][ 135 ],
   alphaCSR[ 133 ][ 136 ],
   alphaCSR[ 133 ][ 137 ],
   alphaCSR[ 133 ][ 138 ],
   alphaCSR[ 133 ][ 139 ],
   alphaCSR[ 133 ][ 140 ],
   alphaCSR[ 133 ][ 141 ],
   alphaCSR[ 133 ][ 142 ],
   alphaCSR[ 133 ][ 143 ],
   alphaCSR[ 133 ][ 144 ],
   alphaCSR[ 133 ][ 145 ],
   alphaCSR[ 133 ][ 146 ],
   alphaCSR[ 133 ][ 147 ],
   alphaCSR[ 133 ][ 148 ],
   alphaCSR[ 133 ][ 149 ],
   alphaCSR[ 133 ][ 150 ],
   alphaCSR[ 133 ][ 151 ],
   alphaCSR[ 133 ][ 152 ],
   alphaCSR[ 133 ][ 153 ],
   alphaCSR[ 133 ][ 154 ],
   alphaCSR[ 133 ][ 155 ],
   alphaCSR[ 133 ][ 156 ],
   alphaCSR[ 133 ][ 157 ],
   alphaCSR[ 133 ][ 158 ],
   alphaCSR[ 133 ][ 159 ],
   alphaCSR[ 133 ][ 160 ],
   alphaCSR[ 133 ][ 161 ],
   alphaCSR[ 133 ][ 162 ],
   alphaCSR[ 133 ][ 163 ],
   alphaCSR[ 133 ][ 164 ],
   alphaCSR[ 133 ][ 165 ],
   alphaCSR[ 133 ][ 166 ],
   alphaCSR[ 133 ][ 167 ],
   alphaCSR[ 133 ][ 168 ],
   alphaCSR[ 133 ][ 169 ],
   alphaCSR[ 133 ][ 170 ],
   alphaCSR[ 133 ][ 171 ],
   alphaCSR[ 133 ][ 172 ],
   alphaCSR[ 133 ][ 173 ],
   alphaCSR[ 133 ][ 174 ],
   alphaCSR[ 133 ][ 175 ],
   alphaCSR[ 133 ][ 176 ],
   alphaCSR[ 133 ][ 177 ],
   alphaCSR[ 133 ][ 178 ],
   alphaCSR[ 133 ][ 179 ],
   alphaCSR[ 133 ][ 180 ],
   alphaCSR[ 133 ][ 181 ],
   alphaCSR[ 133 ][ 182 ],
   alphaCSR[ 133 ][ 183 ],
   alphaCSR[ 133 ][ 184 ],
   alphaCSR[ 133 ][ 185 ],
   alphaCSR[ 133 ][ 186 ],
   alphaCSR[ 133 ][ 187 ],
   alphaCSR[ 133 ][ 188 ],
   alphaCSR[ 133 ][ 189 ],
   alphaCSR[ 133 ][ 190 ],
   alphaCSR[ 133 ][ 191 ],
   alphaCSR[ 133 ][ 192 ],
   alphaCSR[ 133 ][ 193 ],
   alphaCSR[ 133 ][ 194 ],
   alphaCSR[ 133 ][ 195 ],
   alphaCSR[ 133 ][ 196 ],
   alphaCSR[ 133 ][ 197 ],
   alphaCSR[ 133 ][ 198 ],
   alphaCSR[ 133 ][ 199 ],
   alphaCSR[ 133 ][ 200 ],
   alphaCSR[ 133 ][ 201 ],
   alphaCSR[ 133 ][ 202 ],
   alphaCSR[ 133 ][ 203 ],
   alphaCSR[ 133 ][ 204 ],
   alphaCSR[ 133 ][ 205 ],
   alphaCSR[ 133 ][ 206 ],
   alphaCSR[ 133 ][ 207 ],
   alphaCSR[ 133 ][ 208 ],
   alphaCSR[ 133 ][ 209 ],
   alphaCSR[ 133 ][ 210 ],
   alphaCSR[ 133 ][ 211 ],
   alphaCSR[ 133 ][ 212 ],
   alphaCSR[ 133 ][ 213 ],
   alphaCSR[ 133 ][ 214 ],
   alphaCSR[ 133 ][ 215 ],
   alphaCSR[ 133 ][ 216 ],
   alphaCSR[ 133 ][ 217 ],
   alphaCSR[ 133 ][ 218 ],
   alphaCSR[ 133 ][ 219 ],
   alphaCSR[ 133 ][ 220 ],
   alphaCSR[ 133 ][ 221 ],
   alphaCSR[ 133 ][ 222 ],
   alphaCSR[ 133 ][ 223 ],
   alphaCSR[ 133 ][ 224 ],
   alphaCSR[ 133 ][ 225 ],
   alphaCSR[ 133 ][ 226 ],
   alphaCSR[ 133 ][ 227 ],
   alphaCSR[ 133 ][ 228 ],
   alphaCSR[ 133 ][ 229 ],
   alphaCSR[ 133 ][ 230 ],
   alphaCSR[ 133 ][ 231 ],
   alphaCSR[ 133 ][ 232 ],
   alphaCSR[ 133 ][ 233 ],
   alphaCSR[ 133 ][ 234 ],
   alphaCSR[ 133 ][ 235 ],
   alphaCSR[ 133 ][ 236 ],
   alphaCSR[ 133 ][ 237 ],
   alphaCSR[ 133 ][ 238 ],
   alphaCSR[ 133 ][ 239 ],
   alphaCSR[ 133 ][ 240 ],
   alphaCSR[ 133 ][ 241 ],
   alphaCSR[ 133 ][ 242 ],
   alphaCSR[ 133 ][ 243 ],
   alphaCSR[ 133 ][ 244 ],
   alphaCSR[ 133 ][ 245 ],
   alphaCSR[ 133 ][ 246 ],
   alphaCSR[ 133 ][ 247 ],
   alphaCSR[ 133 ][ 248 ],
   alphaCSR[ 133 ][ 249 ],
   alphaCSR[ 133 ][ 250 ],
   alphaCSR[ 133 ][ 251 ],
   alphaCSR[ 133 ][ 252 ],
   alphaCSR[ 133 ][ 253 ],
   alphaCSR[ 133 ][ 254 ],
   alphaCSR[ 133 ][ 255 ],
   alphaCSR[ 133 ][ 256 ],
   alphaCSR[ 133 ][ 257 ],
   alphaCSR[ 133 ][ 258 ],
   alphaCSR[ 133 ][ 259 ],
   alphaCSR[ 133 ][ 260 ],
   alphaCSR[ 133 ][ 261 ],
   alphaCSR[ 133 ][ 262 ],
   alphaCSR[ 133 ][ 263 ],
   alphaCSR[ 133 ][ 264 ],
   alphaCSR[ 133 ][ 265 ],
   alphaCSR[ 133 ][ 266 ],
   alphaCSR[ 133 ][ 267 ],
   alphaCSR[ 133 ][ 268 ],
   alphaCSR[ 133 ][ 269 ],
   alphaCSR[ 133 ][ 270 ],
   alphaCSR[ 133 ][ 271 ],
   alphaCSR[ 133 ][ 272 ],
   alphaCSR[ 133 ][ 273 ],
   alphaCSR[ 133 ][ 274 ],
   alphaCSR[ 133 ][ 275 ],
   alphaCSR[ 133 ][ 276 ],
   alphaCSR[ 133 ][ 277 ],
   alphaCSR[ 133 ][ 278 ],
   alphaCSR[ 133 ][ 279 ],
   alphaCSR[ 133 ][ 280 ],
   alphaCSR[ 133 ][ 281 ],
   alphaCSR[ 133 ][ 282 ],
   alphaCSR[ 133 ][ 283 ],
   alphaCSR[ 133 ][ 284 ],
   alphaCSR[ 133 ][ 285 ],
   alphaCSR[ 133 ][ 286 ],
   alphaCSR[ 133 ][ 287 ],
   alphaCSR[ 133 ][ 288 ],
   alphaCSR[ 133 ][ 289 ],
   alphaCSR[ 133 ][ 290 ],
   alphaCSR[ 133 ][ 291 ],
   alphaCSR[ 133 ][ 292 ],
   alphaCSR[ 133 ][ 293 ],
   alphaCSR[ 133 ][ 294 ],
   alphaCSR[ 133 ][ 295 ],
   alphaCSR[ 133 ][ 296 ],
   alphaCSR[ 133 ][ 297 ],
   alphaCSR[ 133 ][ 298 ],
   alphaCSR[ 133 ][ 299 ],
   alphaCSR[ 133 ][ 300 ],
   alphaCSR[ 133 ][ 301 ],
   alphaCSR[ 133 ][ 302 ],
   alphaCSR[ 133 ][ 303 ],
   alphaCSR[ 133 ][ 304 ],
   alphaCSR[ 133 ][ 305 ],
   alphaCSR[ 133 ][ 306 ],
   alphaCSR[ 133 ][ 307 ],
   alphaCSR[ 133 ][ 308 ],
   alphaCSR[ 133 ][ 309 ],
   alphaCSR[ 133 ][ 310 ],
   alphaCSR[ 133 ][ 311 ],
   alphaCSR[ 133 ][ 312 ],
   alphaCSR[ 133 ][ 313 ],
   alphaCSR[ 133 ][ 314 ],
   alphaCSR[ 133 ][ 315 ],
   alphaCSR[ 133 ][ 316 ],
   alphaCSR[ 133 ][ 317 ],
   alphaCSR[ 133 ][ 318 ],
   alphaCSR[ 133 ][ 319 ],
   alphaCSR[ 133 ][ 320 ],
   alphaCSR[ 133 ][ 321 ],
   alphaCSR[ 133 ][ 322 ],
   alphaCSR[ 133 ][ 323 ],
   alphaCSR[ 133 ][ 324 ],
   alphaCSR[ 133 ][ 325 ],
   alphaCSR[ 133 ][ 326 ],
   alphaCSR[ 133 ][ 327 ],
   alphaCSR[ 133 ][ 328 ],
   alphaCSR[ 133 ][ 329 ],
   alphaCSR[ 133 ][ 330 ],
   alphaCSR[ 133 ][ 331 ],
   alphaCSR[ 133 ][ 332 ],
   alphaCSR[ 133 ][ 333 ],
   alphaCSR[ 133 ][ 334 ],
   alphaCSR[ 133 ][ 335 ],
   alphaCSR[ 133 ][ 336 ],
   alphaCSR[ 133 ][ 337 ],
   alphaCSR[ 133 ][ 338 ],
   alphaCSR[ 133 ][ 339 ],
   alphaCSR[ 133 ][ 340 ],
   alphaCSR[ 133 ][ 341 ],
   alphaCSR[ 133 ][ 342 ],
   alphaCSR[ 133 ][ 343 ],
   alphaCSR[ 133 ][ 344 ],
   alphaCSR[ 133 ][ 345 ],
   alphaCSR[ 133 ][ 346 ],
   alphaCSR[ 133 ][ 347 ],
   alphaCSR[ 133 ][ 348 ],
   alphaCSR[ 133 ][ 349 ],
   alphaCSR[ 133 ][ 350 ],
   alphaCSR[ 133 ][ 351 ],
   alphaCSR[ 133 ][ 352 ],
   alphaCSR[ 133 ][ 353 ],
   alphaCSR[ 133 ][ 354 ],
   alphaCSR[ 133 ][ 355 ],
   alphaCSR[ 133 ][ 356 ],
   alphaCSR[ 133 ][ 357 ],
   alphaCSR[ 133 ][ 358 ],
   alphaCSR[ 133 ][ 359 ],
   alphaCSR[ 133 ][ 360 ],
   alphaCSR[ 133 ][ 361 ],
   alphaCSR[ 133 ][ 362 ],
   alphaCSR[ 133 ][ 363 ],
   alphaCSR[ 133 ][ 364 ],
   alphaCSR[ 133 ][ 365 ],
   alphaCSR[ 133 ][ 366 ],
   alphaCSR[ 133 ][ 367 ],
   alphaCSR[ 133 ][ 368 ],
   alphaCSR[ 133 ][ 369 ],
   alphaCSR[ 133 ][ 370 ],
   alphaCSR[ 133 ][ 371 ],
   alphaCSR[ 133 ][ 372 ],
   alphaCSR[ 133 ][ 373 ],
   alphaCSR[ 133 ][ 374 ],
   alphaCSR[ 133 ][ 375 ],
   alphaCSR[ 133 ][ 376 ],
   alphaCSR[ 133 ][ 377 ],
   alphaCSR[ 133 ][ 378 ],
   alphaCSR[ 133 ][ 379 ],
   alphaCSR[ 133 ][ 380 ],
   alphaCSR[ 133 ][ 381 ],
   alphaCSR[ 133 ][ 382 ],
   alphaCSR[ 133 ][ 383 ],
   alphaCSR[ 134 ][ 0 ],
   alphaCSR[ 134 ][ 1 ],
   alphaCSR[ 134 ][ 2 ],
   alphaCSR[ 134 ][ 3 ],
   alphaCSR[ 134 ][ 4 ],
   alphaCSR[ 134 ][ 5 ],
   alphaCSR[ 134 ][ 6 ],
   alphaCSR[ 134 ][ 7 ],
   alphaCSR[ 134 ][ 8 ],
   alphaCSR[ 134 ][ 9 ],
   alphaCSR[ 134 ][ 10 ],
   alphaCSR[ 134 ][ 11 ],
   alphaCSR[ 134 ][ 12 ],
   alphaCSR[ 134 ][ 13 ],
   alphaCSR[ 134 ][ 14 ],
   alphaCSR[ 134 ][ 15 ],
   alphaCSR[ 134 ][ 16 ],
   alphaCSR[ 134 ][ 17 ],
   alphaCSR[ 134 ][ 18 ],
   alphaCSR[ 134 ][ 19 ],
   alphaCSR[ 134 ][ 20 ],
   alphaCSR[ 134 ][ 21 ],
   alphaCSR[ 134 ][ 22 ],
   alphaCSR[ 134 ][ 23 ],
   alphaCSR[ 134 ][ 24 ],
   alphaCSR[ 134 ][ 25 ],
   alphaCSR[ 134 ][ 26 ],
   alphaCSR[ 134 ][ 27 ],
   alphaCSR[ 134 ][ 28 ],
   alphaCSR[ 134 ][ 29 ],
   alphaCSR[ 134 ][ 30 ],
   alphaCSR[ 134 ][ 31 ],
   alphaCSR[ 134 ][ 32 ],
   alphaCSR[ 134 ][ 33 ],
   alphaCSR[ 134 ][ 34 ],
   alphaCSR[ 134 ][ 35 ],
   alphaCSR[ 134 ][ 36 ],
   alphaCSR[ 134 ][ 37 ],
   alphaCSR[ 134 ][ 38 ],
   alphaCSR[ 134 ][ 39 ],
   alphaCSR[ 134 ][ 40 ],
   alphaCSR[ 134 ][ 41 ],
   alphaCSR[ 134 ][ 42 ],
   alphaCSR[ 134 ][ 43 ],
   alphaCSR[ 134 ][ 44 ],
   alphaCSR[ 134 ][ 45 ],
   alphaCSR[ 134 ][ 46 ],
   alphaCSR[ 134 ][ 47 ],
   alphaCSR[ 134 ][ 48 ],
   alphaCSR[ 134 ][ 49 ],
   alphaCSR[ 134 ][ 50 ],
   alphaCSR[ 134 ][ 51 ],
   alphaCSR[ 134 ][ 52 ],
   alphaCSR[ 134 ][ 53 ],
   alphaCSR[ 134 ][ 54 ],
   alphaCSR[ 134 ][ 55 ],
   alphaCSR[ 134 ][ 56 ],
   alphaCSR[ 134 ][ 57 ],
   alphaCSR[ 134 ][ 58 ],
   alphaCSR[ 134 ][ 59 ],
   alphaCSR[ 134 ][ 60 ],
   alphaCSR[ 134 ][ 61 ],
   alphaCSR[ 134 ][ 62 ],
   alphaCSR[ 134 ][ 63 ],
   alphaCSR[ 134 ][ 64 ],
   alphaCSR[ 134 ][ 65 ],
   alphaCSR[ 134 ][ 66 ],
   alphaCSR[ 134 ][ 67 ],
   alphaCSR[ 134 ][ 68 ],
   alphaCSR[ 134 ][ 69 ],
   alphaCSR[ 134 ][ 70 ],
   alphaCSR[ 134 ][ 71 ],
   alphaCSR[ 134 ][ 72 ],
   alphaCSR[ 134 ][ 73 ],
   alphaCSR[ 134 ][ 74 ],
   alphaCSR[ 134 ][ 75 ],
   alphaCSR[ 134 ][ 76 ],
   alphaCSR[ 134 ][ 77 ],
   alphaCSR[ 134 ][ 78 ],
   alphaCSR[ 134 ][ 79 ],
   alphaCSR[ 134 ][ 80 ],
   alphaCSR[ 134 ][ 81 ],
   alphaCSR[ 134 ][ 82 ],
   alphaCSR[ 134 ][ 83 ],
   alphaCSR[ 134 ][ 84 ],
   alphaCSR[ 134 ][ 85 ],
   alphaCSR[ 134 ][ 86 ],
   alphaCSR[ 134 ][ 87 ],
   alphaCSR[ 134 ][ 88 ],
   alphaCSR[ 134 ][ 89 ],
   alphaCSR[ 134 ][ 90 ],
   alphaCSR[ 134 ][ 91 ],
   alphaCSR[ 134 ][ 92 ],
   alphaCSR[ 134 ][ 93 ],
   alphaCSR[ 134 ][ 94 ],
   alphaCSR[ 134 ][ 95 ],
   alphaCSR[ 134 ][ 96 ],
   alphaCSR[ 134 ][ 97 ],
   alphaCSR[ 134 ][ 98 ],
   alphaCSR[ 134 ][ 99 ],
   alphaCSR[ 134 ][ 100 ],
   alphaCSR[ 134 ][ 101 ],
   alphaCSR[ 134 ][ 102 ],
   alphaCSR[ 134 ][ 103 ],
   alphaCSR[ 134 ][ 104 ],
   alphaCSR[ 134 ][ 105 ],
   alphaCSR[ 134 ][ 106 ],
   alphaCSR[ 134 ][ 107 ],
   alphaCSR[ 134 ][ 108 ],
   alphaCSR[ 134 ][ 109 ],
   alphaCSR[ 134 ][ 110 ],
   alphaCSR[ 134 ][ 111 ],
   alphaCSR[ 134 ][ 112 ],
   alphaCSR[ 134 ][ 113 ],
   alphaCSR[ 134 ][ 114 ],
   alphaCSR[ 134 ][ 115 ],
   alphaCSR[ 134 ][ 116 ],
   alphaCSR[ 134 ][ 117 ],
   alphaCSR[ 134 ][ 118 ],
   alphaCSR[ 134 ][ 119 ],
   alphaCSR[ 134 ][ 120 ],
   alphaCSR[ 134 ][ 121 ],
   alphaCSR[ 134 ][ 122 ],
   alphaCSR[ 134 ][ 123 ],
   alphaCSR[ 134 ][ 124 ],
   alphaCSR[ 134 ][ 125 ],
   alphaCSR[ 134 ][ 126 ],
   alphaCSR[ 134 ][ 127 ],
   alphaCSR[ 134 ][ 128 ],
   alphaCSR[ 134 ][ 129 ],
   alphaCSR[ 134 ][ 130 ],
   alphaCSR[ 134 ][ 131 ],
   alphaCSR[ 134 ][ 132 ],
   alphaCSR[ 134 ][ 133 ],
   alphaCSR[ 134 ][ 134 ],
   alphaCSR[ 134 ][ 135 ],
   alphaCSR[ 134 ][ 136 ],
   alphaCSR[ 134 ][ 137 ],
   alphaCSR[ 134 ][ 138 ],
   alphaCSR[ 134 ][ 139 ],
   alphaCSR[ 134 ][ 140 ],
   alphaCSR[ 134 ][ 141 ],
   alphaCSR[ 134 ][ 142 ],
   alphaCSR[ 134 ][ 143 ],
   alphaCSR[ 134 ][ 144 ],
   alphaCSR[ 134 ][ 145 ],
   alphaCSR[ 134 ][ 146 ],
   alphaCSR[ 134 ][ 147 ],
   alphaCSR[ 134 ][ 148 ],
   alphaCSR[ 134 ][ 149 ],
   alphaCSR[ 134 ][ 150 ],
   alphaCSR[ 134 ][ 151 ],
   alphaCSR[ 134 ][ 152 ],
   alphaCSR[ 134 ][ 153 ],
   alphaCSR[ 134 ][ 154 ],
   alphaCSR[ 134 ][ 155 ],
   alphaCSR[ 134 ][ 156 ],
   alphaCSR[ 134 ][ 157 ],
   alphaCSR[ 134 ][ 158 ],
   alphaCSR[ 134 ][ 159 ],
   alphaCSR[ 134 ][ 160 ],
   alphaCSR[ 134 ][ 161 ],
   alphaCSR[ 134 ][ 162 ],
   alphaCSR[ 134 ][ 163 ],
   alphaCSR[ 134 ][ 164 ],
   alphaCSR[ 134 ][ 165 ],
   alphaCSR[ 134 ][ 166 ],
   alphaCSR[ 134 ][ 167 ],
   alphaCSR[ 134 ][ 168 ],
   alphaCSR[ 134 ][ 169 ],
   alphaCSR[ 134 ][ 170 ],
   alphaCSR[ 134 ][ 171 ],
   alphaCSR[ 134 ][ 172 ],
   alphaCSR[ 134 ][ 173 ],
   alphaCSR[ 134 ][ 174 ],
   alphaCSR[ 134 ][ 175 ],
   alphaCSR[ 134 ][ 176 ],
   alphaCSR[ 134 ][ 177 ],
   alphaCSR[ 134 ][ 178 ],
   alphaCSR[ 134 ][ 179 ],
   alphaCSR[ 134 ][ 180 ],
   alphaCSR[ 134 ][ 181 ],
   alphaCSR[ 134 ][ 182 ],
   alphaCSR[ 134 ][ 183 ],
   alphaCSR[ 134 ][ 184 ],
   alphaCSR[ 134 ][ 185 ],
   alphaCSR[ 134 ][ 186 ],
   alphaCSR[ 134 ][ 187 ],
   alphaCSR[ 134 ][ 188 ],
   alphaCSR[ 134 ][ 189 ],
   alphaCSR[ 134 ][ 190 ],
   alphaCSR[ 134 ][ 191 ],
   alphaCSR[ 134 ][ 192 ],
   alphaCSR[ 134 ][ 193 ],
   alphaCSR[ 134 ][ 194 ],
   alphaCSR[ 134 ][ 195 ],
   alphaCSR[ 134 ][ 196 ],
   alphaCSR[ 134 ][ 197 ],
   alphaCSR[ 134 ][ 198 ],
   alphaCSR[ 134 ][ 199 ],
   alphaCSR[ 134 ][ 200 ],
   alphaCSR[ 134 ][ 201 ],
   alphaCSR[ 134 ][ 202 ],
   alphaCSR[ 134 ][ 203 ],
   alphaCSR[ 134 ][ 204 ],
   alphaCSR[ 134 ][ 205 ],
   alphaCSR[ 134 ][ 206 ],
   alphaCSR[ 134 ][ 207 ],
   alphaCSR[ 134 ][ 208 ],
   alphaCSR[ 134 ][ 209 ],
   alphaCSR[ 134 ][ 210 ],
   alphaCSR[ 134 ][ 211 ],
   alphaCSR[ 134 ][ 212 ],
   alphaCSR[ 134 ][ 213 ],
   alphaCSR[ 134 ][ 214 ],
   alphaCSR[ 134 ][ 215 ],
   alphaCSR[ 134 ][ 216 ],
   alphaCSR[ 134 ][ 217 ],
   alphaCSR[ 134 ][ 218 ],
   alphaCSR[ 134 ][ 219 ],
   alphaCSR[ 134 ][ 220 ],
   alphaCSR[ 134 ][ 221 ],
   alphaCSR[ 134 ][ 222 ],
   alphaCSR[ 134 ][ 223 ],
   alphaCSR[ 134 ][ 224 ],
   alphaCSR[ 134 ][ 225 ],
   alphaCSR[ 134 ][ 226 ],
   alphaCSR[ 134 ][ 227 ],
   alphaCSR[ 134 ][ 228 ],
   alphaCSR[ 134 ][ 229 ],
   alphaCSR[ 134 ][ 230 ],
   alphaCSR[ 134 ][ 231 ],
   alphaCSR[ 134 ][ 232 ],
   alphaCSR[ 134 ][ 233 ],
   alphaCSR[ 134 ][ 234 ],
   alphaCSR[ 134 ][ 235 ],
   alphaCSR[ 134 ][ 236 ],
   alphaCSR[ 134 ][ 237 ],
   alphaCSR[ 134 ][ 238 ],
   alphaCSR[ 134 ][ 239 ],
   alphaCSR[ 134 ][ 240 ],
   alphaCSR[ 134 ][ 241 ],
   alphaCSR[ 134 ][ 242 ],
   alphaCSR[ 134 ][ 243 ],
   alphaCSR[ 134 ][ 244 ],
   alphaCSR[ 134 ][ 245 ],
   alphaCSR[ 134 ][ 246 ],
   alphaCSR[ 134 ][ 247 ],
   alphaCSR[ 134 ][ 248 ],
   alphaCSR[ 134 ][ 249 ],
   alphaCSR[ 134 ][ 250 ],
   alphaCSR[ 134 ][ 251 ],
   alphaCSR[ 134 ][ 252 ],
   alphaCSR[ 134 ][ 253 ],
   alphaCSR[ 134 ][ 254 ],
   alphaCSR[ 134 ][ 255 ],
   alphaCSR[ 134 ][ 256 ],
   alphaCSR[ 134 ][ 257 ],
   alphaCSR[ 134 ][ 258 ],
   alphaCSR[ 134 ][ 259 ],
   alphaCSR[ 134 ][ 260 ],
   alphaCSR[ 134 ][ 261 ],
   alphaCSR[ 134 ][ 262 ],
   alphaCSR[ 134 ][ 263 ],
   alphaCSR[ 134 ][ 264 ],
   alphaCSR[ 134 ][ 265 ],
   alphaCSR[ 134 ][ 266 ],
   alphaCSR[ 134 ][ 267 ],
   alphaCSR[ 134 ][ 268 ],
   alphaCSR[ 134 ][ 269 ],
   alphaCSR[ 134 ][ 270 ],
   alphaCSR[ 134 ][ 271 ],
   alphaCSR[ 134 ][ 272 ],
   alphaCSR[ 134 ][ 273 ],
   alphaCSR[ 134 ][ 274 ],
   alphaCSR[ 134 ][ 275 ],
   alphaCSR[ 134 ][ 276 ],
   alphaCSR[ 134 ][ 277 ],
   alphaCSR[ 134 ][ 278 ],
   alphaCSR[ 134 ][ 279 ],
   alphaCSR[ 134 ][ 280 ],
   alphaCSR[ 134 ][ 281 ],
   alphaCSR[ 134 ][ 282 ],
   alphaCSR[ 134 ][ 283 ],
   alphaCSR[ 134 ][ 284 ],
   alphaCSR[ 134 ][ 285 ],
   alphaCSR[ 134 ][ 286 ],
   alphaCSR[ 134 ][ 287 ],
   alphaCSR[ 134 ][ 288 ],
   alphaCSR[ 134 ][ 289 ],
   alphaCSR[ 134 ][ 290 ],
   alphaCSR[ 134 ][ 291 ],
   alphaCSR[ 134 ][ 292 ],
   alphaCSR[ 134 ][ 293 ],
   alphaCSR[ 134 ][ 294 ],
   alphaCSR[ 134 ][ 295 ],
   alphaCSR[ 134 ][ 296 ],
   alphaCSR[ 134 ][ 297 ],
   alphaCSR[ 134 ][ 298 ],
   alphaCSR[ 134 ][ 299 ],
   alphaCSR[ 134 ][ 300 ],
   alphaCSR[ 134 ][ 301 ],
   alphaCSR[ 134 ][ 302 ],
   alphaCSR[ 134 ][ 303 ],
   alphaCSR[ 134 ][ 304 ],
   alphaCSR[ 134 ][ 305 ],
   alphaCSR[ 134 ][ 306 ],
   alphaCSR[ 134 ][ 307 ],
   alphaCSR[ 134 ][ 308 ],
   alphaCSR[ 134 ][ 309 ],
   alphaCSR[ 134 ][ 310 ],
   alphaCSR[ 134 ][ 311 ],
   alphaCSR[ 134 ][ 312 ],
   alphaCSR[ 134 ][ 313 ],
   alphaCSR[ 134 ][ 314 ],
   alphaCSR[ 134 ][ 315 ],
   alphaCSR[ 134 ][ 316 ],
   alphaCSR[ 134 ][ 317 ],
   alphaCSR[ 134 ][ 318 ],
   alphaCSR[ 134 ][ 319 ],
   alphaCSR[ 134 ][ 320 ],
   alphaCSR[ 134 ][ 321 ],
   alphaCSR[ 134 ][ 322 ],
   alphaCSR[ 134 ][ 323 ],
   alphaCSR[ 134 ][ 324 ],
   alphaCSR[ 134 ][ 325 ],
   alphaCSR[ 134 ][ 326 ],
   alphaCSR[ 134 ][ 327 ],
   alphaCSR[ 134 ][ 328 ],
   alphaCSR[ 134 ][ 329 ],
   alphaCSR[ 134 ][ 330 ],
   alphaCSR[ 134 ][ 331 ],
   alphaCSR[ 134 ][ 332 ],
   alphaCSR[ 134 ][ 333 ],
   alphaCSR[ 134 ][ 334 ],
   alphaCSR[ 134 ][ 335 ],
   alphaCSR[ 134 ][ 336 ],
   alphaCSR[ 134 ][ 337 ],
   alphaCSR[ 134 ][ 338 ],
   alphaCSR[ 134 ][ 339 ],
   alphaCSR[ 134 ][ 340 ],
   alphaCSR[ 134 ][ 341 ],
   alphaCSR[ 134 ][ 342 ],
   alphaCSR[ 134 ][ 343 ],
   alphaCSR[ 134 ][ 344 ],
   alphaCSR[ 134 ][ 345 ],
   alphaCSR[ 134 ][ 346 ],
   alphaCSR[ 134 ][ 347 ],
   alphaCSR[ 134 ][ 348 ],
   alphaCSR[ 134 ][ 349 ],
   alphaCSR[ 134 ][ 350 ],
   alphaCSR[ 134 ][ 351 ],
   alphaCSR[ 134 ][ 352 ],
   alphaCSR[ 134 ][ 353 ],
   alphaCSR[ 134 ][ 354 ],
   alphaCSR[ 134 ][ 355 ],
   alphaCSR[ 134 ][ 356 ],
   alphaCSR[ 134 ][ 357 ],
   alphaCSR[ 134 ][ 358 ],
   alphaCSR[ 134 ][ 359 ],
   alphaCSR[ 134 ][ 360 ],
   alphaCSR[ 134 ][ 361 ],
   alphaCSR[ 134 ][ 362 ],
   alphaCSR[ 134 ][ 363 ],
   alphaCSR[ 134 ][ 364 ],
   alphaCSR[ 134 ][ 365 ],
   alphaCSR[ 134 ][ 366 ],
   alphaCSR[ 134 ][ 367 ],
   alphaCSR[ 134 ][ 368 ],
   alphaCSR[ 134 ][ 369 ],
   alphaCSR[ 134 ][ 370 ],
   alphaCSR[ 134 ][ 371 ],
   alphaCSR[ 134 ][ 372 ],
   alphaCSR[ 134 ][ 373 ],
   alphaCSR[ 134 ][ 374 ],
   alphaCSR[ 134 ][ 375 ],
   alphaCSR[ 134 ][ 376 ],
   alphaCSR[ 134 ][ 377 ],
   alphaCSR[ 134 ][ 378 ],
   alphaCSR[ 134 ][ 379 ],
   alphaCSR[ 134 ][ 380 ],
   alphaCSR[ 134 ][ 381 ],
   alphaCSR[ 134 ][ 382 ],
   alphaCSR[ 134 ][ 383 ],
   alphaCSR[ 135 ][ 0 ],
   alphaCSR[ 135 ][ 1 ],
   alphaCSR[ 135 ][ 2 ],
   alphaCSR[ 135 ][ 3 ],
   alphaCSR[ 135 ][ 4 ],
   alphaCSR[ 135 ][ 5 ],
   alphaCSR[ 135 ][ 6 ],
   alphaCSR[ 135 ][ 7 ],
   alphaCSR[ 135 ][ 8 ],
   alphaCSR[ 135 ][ 9 ],
   alphaCSR[ 135 ][ 10 ],
   alphaCSR[ 135 ][ 11 ],
   alphaCSR[ 135 ][ 12 ],
   alphaCSR[ 135 ][ 13 ],
   alphaCSR[ 135 ][ 14 ],
   alphaCSR[ 135 ][ 15 ],
   alphaCSR[ 135 ][ 16 ],
   alphaCSR[ 135 ][ 17 ],
   alphaCSR[ 135 ][ 18 ],
   alphaCSR[ 135 ][ 19 ],
   alphaCSR[ 135 ][ 20 ],
   alphaCSR[ 135 ][ 21 ],
   alphaCSR[ 135 ][ 22 ],
   alphaCSR[ 135 ][ 23 ],
   alphaCSR[ 135 ][ 24 ],
   alphaCSR[ 135 ][ 25 ],
   alphaCSR[ 135 ][ 26 ],
   alphaCSR[ 135 ][ 27 ],
   alphaCSR[ 135 ][ 28 ],
   alphaCSR[ 135 ][ 29 ],
   alphaCSR[ 135 ][ 30 ],
   alphaCSR[ 135 ][ 31 ],
   alphaCSR[ 135 ][ 32 ],
   alphaCSR[ 135 ][ 33 ],
   alphaCSR[ 135 ][ 34 ],
   alphaCSR[ 135 ][ 35 ],
   alphaCSR[ 135 ][ 36 ],
   alphaCSR[ 135 ][ 37 ],
   alphaCSR[ 135 ][ 38 ],
   alphaCSR[ 135 ][ 39 ],
   alphaCSR[ 135 ][ 40 ],
   alphaCSR[ 135 ][ 41 ],
   alphaCSR[ 135 ][ 42 ],
   alphaCSR[ 135 ][ 43 ],
   alphaCSR[ 135 ][ 44 ],
   alphaCSR[ 135 ][ 45 ],
   alphaCSR[ 135 ][ 46 ],
   alphaCSR[ 135 ][ 47 ],
   alphaCSR[ 135 ][ 48 ],
   alphaCSR[ 135 ][ 49 ],
   alphaCSR[ 135 ][ 50 ],
   alphaCSR[ 135 ][ 51 ],
   alphaCSR[ 135 ][ 52 ],
   alphaCSR[ 135 ][ 53 ],
   alphaCSR[ 135 ][ 54 ],
   alphaCSR[ 135 ][ 55 ],
   alphaCSR[ 135 ][ 56 ],
   alphaCSR[ 135 ][ 57 ],
   alphaCSR[ 135 ][ 58 ],
   alphaCSR[ 135 ][ 59 ],
   alphaCSR[ 135 ][ 60 ],
   alphaCSR[ 135 ][ 61 ],
   alphaCSR[ 135 ][ 62 ],
   alphaCSR[ 135 ][ 63 ],
   alphaCSR[ 135 ][ 64 ],
   alphaCSR[ 135 ][ 65 ],
   alphaCSR[ 135 ][ 66 ],
   alphaCSR[ 135 ][ 67 ],
   alphaCSR[ 135 ][ 68 ],
   alphaCSR[ 135 ][ 69 ],
   alphaCSR[ 135 ][ 70 ],
   alphaCSR[ 135 ][ 71 ],
   alphaCSR[ 135 ][ 72 ],
   alphaCSR[ 135 ][ 73 ],
   alphaCSR[ 135 ][ 74 ],
   alphaCSR[ 135 ][ 75 ],
   alphaCSR[ 135 ][ 76 ],
   alphaCSR[ 135 ][ 77 ],
   alphaCSR[ 135 ][ 78 ],
   alphaCSR[ 135 ][ 79 ],
   alphaCSR[ 135 ][ 80 ],
   alphaCSR[ 135 ][ 81 ],
   alphaCSR[ 135 ][ 82 ],
   alphaCSR[ 135 ][ 83 ],
   alphaCSR[ 135 ][ 84 ],
   alphaCSR[ 135 ][ 85 ],
   alphaCSR[ 135 ][ 86 ],
   alphaCSR[ 135 ][ 87 ],
   alphaCSR[ 135 ][ 88 ],
   alphaCSR[ 135 ][ 89 ],
   alphaCSR[ 135 ][ 90 ],
   alphaCSR[ 135 ][ 91 ],
   alphaCSR[ 135 ][ 92 ],
   alphaCSR[ 135 ][ 93 ],
   alphaCSR[ 135 ][ 94 ],
   alphaCSR[ 135 ][ 95 ],
   alphaCSR[ 135 ][ 96 ],
   alphaCSR[ 135 ][ 97 ],
   alphaCSR[ 135 ][ 98 ],
   alphaCSR[ 135 ][ 99 ],
   alphaCSR[ 135 ][ 100 ],
   alphaCSR[ 135 ][ 101 ],
   alphaCSR[ 135 ][ 102 ],
   alphaCSR[ 135 ][ 103 ],
   alphaCSR[ 135 ][ 104 ],
   alphaCSR[ 135 ][ 105 ],
   alphaCSR[ 135 ][ 106 ],
   alphaCSR[ 135 ][ 107 ],
   alphaCSR[ 135 ][ 108 ],
   alphaCSR[ 135 ][ 109 ],
   alphaCSR[ 135 ][ 110 ],
   alphaCSR[ 135 ][ 111 ],
   alphaCSR[ 135 ][ 112 ],
   alphaCSR[ 135 ][ 113 ],
   alphaCSR[ 135 ][ 114 ],
   alphaCSR[ 135 ][ 115 ],
   alphaCSR[ 135 ][ 116 ],
   alphaCSR[ 135 ][ 117 ],
   alphaCSR[ 135 ][ 118 ],
   alphaCSR[ 135 ][ 119 ],
   alphaCSR[ 135 ][ 120 ],
   alphaCSR[ 135 ][ 121 ],
   alphaCSR[ 135 ][ 122 ],
   alphaCSR[ 135 ][ 123 ],
   alphaCSR[ 135 ][ 124 ],
   alphaCSR[ 135 ][ 125 ],
   alphaCSR[ 135 ][ 126 ],
   alphaCSR[ 135 ][ 127 ],
   alphaCSR[ 135 ][ 128 ],
   alphaCSR[ 135 ][ 129 ],
   alphaCSR[ 135 ][ 130 ],
   alphaCSR[ 135 ][ 131 ],
   alphaCSR[ 135 ][ 132 ],
   alphaCSR[ 135 ][ 133 ],
   alphaCSR[ 135 ][ 134 ],
   alphaCSR[ 135 ][ 135 ],
   alphaCSR[ 135 ][ 136 ],
   alphaCSR[ 135 ][ 137 ],
   alphaCSR[ 135 ][ 138 ],
   alphaCSR[ 135 ][ 139 ],
   alphaCSR[ 135 ][ 140 ],
   alphaCSR[ 135 ][ 141 ],
   alphaCSR[ 135 ][ 142 ],
   alphaCSR[ 135 ][ 143 ],
   alphaCSR[ 135 ][ 144 ],
   alphaCSR[ 135 ][ 145 ],
   alphaCSR[ 135 ][ 146 ],
   alphaCSR[ 135 ][ 147 ],
   alphaCSR[ 135 ][ 148 ],
   alphaCSR[ 135 ][ 149 ],
   alphaCSR[ 135 ][ 150 ],
   alphaCSR[ 135 ][ 151 ],
   alphaCSR[ 135 ][ 152 ],
   alphaCSR[ 135 ][ 153 ],
   alphaCSR[ 135 ][ 154 ],
   alphaCSR[ 135 ][ 155 ],
   alphaCSR[ 135 ][ 156 ],
   alphaCSR[ 135 ][ 157 ],
   alphaCSR[ 135 ][ 158 ],
   alphaCSR[ 135 ][ 159 ],
   alphaCSR[ 135 ][ 160 ],
   alphaCSR[ 135 ][ 161 ],
   alphaCSR[ 135 ][ 162 ],
   alphaCSR[ 135 ][ 163 ],
   alphaCSR[ 135 ][ 164 ],
   alphaCSR[ 135 ][ 165 ],
   alphaCSR[ 135 ][ 166 ],
   alphaCSR[ 135 ][ 167 ],
   alphaCSR[ 135 ][ 168 ],
   alphaCSR[ 135 ][ 169 ],
   alphaCSR[ 135 ][ 170 ],
   alphaCSR[ 135 ][ 171 ],
   alphaCSR[ 135 ][ 172 ],
   alphaCSR[ 135 ][ 173 ],
   alphaCSR[ 135 ][ 174 ],
   alphaCSR[ 135 ][ 175 ],
   alphaCSR[ 135 ][ 176 ],
   alphaCSR[ 135 ][ 177 ],
   alphaCSR[ 135 ][ 178 ],
   alphaCSR[ 135 ][ 179 ],
   alphaCSR[ 135 ][ 180 ],
   alphaCSR[ 135 ][ 181 ],
   alphaCSR[ 135 ][ 182 ],
   alphaCSR[ 135 ][ 183 ],
   alphaCSR[ 135 ][ 184 ],
   alphaCSR[ 135 ][ 185 ],
   alphaCSR[ 135 ][ 186 ],
   alphaCSR[ 135 ][ 187 ],
   alphaCSR[ 135 ][ 188 ],
   alphaCSR[ 135 ][ 189 ],
   alphaCSR[ 135 ][ 190 ],
   alphaCSR[ 135 ][ 191 ],
   alphaCSR[ 135 ][ 192 ],
   alphaCSR[ 135 ][ 193 ],
   alphaCSR[ 135 ][ 194 ],
   alphaCSR[ 135 ][ 195 ],
   alphaCSR[ 135 ][ 196 ],
   alphaCSR[ 135 ][ 197 ],
   alphaCSR[ 135 ][ 198 ],
   alphaCSR[ 135 ][ 199 ],
   alphaCSR[ 135 ][ 200 ],
   alphaCSR[ 135 ][ 201 ],
   alphaCSR[ 135 ][ 202 ],
   alphaCSR[ 135 ][ 203 ],
   alphaCSR[ 135 ][ 204 ],
   alphaCSR[ 135 ][ 205 ],
   alphaCSR[ 135 ][ 206 ],
   alphaCSR[ 135 ][ 207 ],
   alphaCSR[ 135 ][ 208 ],
   alphaCSR[ 135 ][ 209 ],
   alphaCSR[ 135 ][ 210 ],
   alphaCSR[ 135 ][ 211 ],
   alphaCSR[ 135 ][ 212 ],
   alphaCSR[ 135 ][ 213 ],
   alphaCSR[ 135 ][ 214 ],
   alphaCSR[ 135 ][ 215 ],
   alphaCSR[ 135 ][ 216 ],
   alphaCSR[ 135 ][ 217 ],
   alphaCSR[ 135 ][ 218 ],
   alphaCSR[ 135 ][ 219 ],
   alphaCSR[ 135 ][ 220 ],
   alphaCSR[ 135 ][ 221 ],
   alphaCSR[ 135 ][ 222 ],
   alphaCSR[ 135 ][ 223 ],
   alphaCSR[ 135 ][ 224 ],
   alphaCSR[ 135 ][ 225 ],
   alphaCSR[ 135 ][ 226 ],
   alphaCSR[ 135 ][ 227 ],
   alphaCSR[ 135 ][ 228 ],
   alphaCSR[ 135 ][ 229 ],
   alphaCSR[ 135 ][ 230 ],
   alphaCSR[ 135 ][ 231 ],
   alphaCSR[ 135 ][ 232 ],
   alphaCSR[ 135 ][ 233 ],
   alphaCSR[ 135 ][ 234 ],
   alphaCSR[ 135 ][ 235 ],
   alphaCSR[ 135 ][ 236 ],
   alphaCSR[ 135 ][ 237 ],
   alphaCSR[ 135 ][ 238 ],
   alphaCSR[ 135 ][ 239 ],
   alphaCSR[ 135 ][ 240 ],
   alphaCSR[ 135 ][ 241 ],
   alphaCSR[ 135 ][ 242 ],
   alphaCSR[ 135 ][ 243 ],
   alphaCSR[ 135 ][ 244 ],
   alphaCSR[ 135 ][ 245 ],
   alphaCSR[ 135 ][ 246 ],
   alphaCSR[ 135 ][ 247 ],
   alphaCSR[ 135 ][ 248 ],
   alphaCSR[ 135 ][ 249 ],
   alphaCSR[ 135 ][ 250 ],
   alphaCSR[ 135 ][ 251 ],
   alphaCSR[ 135 ][ 252 ],
   alphaCSR[ 135 ][ 253 ],
   alphaCSR[ 135 ][ 254 ],
   alphaCSR[ 135 ][ 255 ],
   alphaCSR[ 135 ][ 256 ],
   alphaCSR[ 135 ][ 257 ],
   alphaCSR[ 135 ][ 258 ],
   alphaCSR[ 135 ][ 259 ],
   alphaCSR[ 135 ][ 260 ],
   alphaCSR[ 135 ][ 261 ],
   alphaCSR[ 135 ][ 262 ],
   alphaCSR[ 135 ][ 263 ],
   alphaCSR[ 135 ][ 264 ],
   alphaCSR[ 135 ][ 265 ],
   alphaCSR[ 135 ][ 266 ],
   alphaCSR[ 135 ][ 267 ],
   alphaCSR[ 135 ][ 268 ],
   alphaCSR[ 135 ][ 269 ],
   alphaCSR[ 135 ][ 270 ],
   alphaCSR[ 135 ][ 271 ],
   alphaCSR[ 135 ][ 272 ],
   alphaCSR[ 135 ][ 273 ],
   alphaCSR[ 135 ][ 274 ],
   alphaCSR[ 135 ][ 275 ],
   alphaCSR[ 135 ][ 276 ],
   alphaCSR[ 135 ][ 277 ],
   alphaCSR[ 135 ][ 278 ],
   alphaCSR[ 135 ][ 279 ],
   alphaCSR[ 135 ][ 280 ],
   alphaCSR[ 135 ][ 281 ],
   alphaCSR[ 135 ][ 282 ],
   alphaCSR[ 135 ][ 283 ],
   alphaCSR[ 135 ][ 284 ],
   alphaCSR[ 135 ][ 285 ],
   alphaCSR[ 135 ][ 286 ],
   alphaCSR[ 135 ][ 287 ],
   alphaCSR[ 135 ][ 288 ],
   alphaCSR[ 135 ][ 289 ],
   alphaCSR[ 135 ][ 290 ],
   alphaCSR[ 135 ][ 291 ],
   alphaCSR[ 135 ][ 292 ],
   alphaCSR[ 135 ][ 293 ],
   alphaCSR[ 135 ][ 294 ],
   alphaCSR[ 135 ][ 295 ],
   alphaCSR[ 135 ][ 296 ],
   alphaCSR[ 135 ][ 297 ],
   alphaCSR[ 135 ][ 298 ],
   alphaCSR[ 135 ][ 299 ],
   alphaCSR[ 135 ][ 300 ],
   alphaCSR[ 135 ][ 301 ],
   alphaCSR[ 135 ][ 302 ],
   alphaCSR[ 135 ][ 303 ],
   alphaCSR[ 135 ][ 304 ],
   alphaCSR[ 135 ][ 305 ],
   alphaCSR[ 135 ][ 306 ],
   alphaCSR[ 135 ][ 307 ],
   alphaCSR[ 135 ][ 308 ],
   alphaCSR[ 135 ][ 309 ],
   alphaCSR[ 135 ][ 310 ],
   alphaCSR[ 135 ][ 311 ],
   alphaCSR[ 135 ][ 312 ],
   alphaCSR[ 135 ][ 313 ],
   alphaCSR[ 135 ][ 314 ],
   alphaCSR[ 135 ][ 315 ],
   alphaCSR[ 135 ][ 316 ],
   alphaCSR[ 135 ][ 317 ],
   alphaCSR[ 135 ][ 318 ],
   alphaCSR[ 135 ][ 319 ],
   alphaCSR[ 135 ][ 320 ],
   alphaCSR[ 135 ][ 321 ],
   alphaCSR[ 135 ][ 322 ],
   alphaCSR[ 135 ][ 323 ],
   alphaCSR[ 135 ][ 324 ],
   alphaCSR[ 135 ][ 325 ],
   alphaCSR[ 135 ][ 326 ],
   alphaCSR[ 135 ][ 327 ],
   alphaCSR[ 135 ][ 328 ],
   alphaCSR[ 135 ][ 329 ],
   alphaCSR[ 135 ][ 330 ],
   alphaCSR[ 135 ][ 331 ],
   alphaCSR[ 135 ][ 332 ],
   alphaCSR[ 135 ][ 333 ],
   alphaCSR[ 135 ][ 334 ],
   alphaCSR[ 135 ][ 335 ],
   alphaCSR[ 135 ][ 336 ],
   alphaCSR[ 135 ][ 337 ],
   alphaCSR[ 135 ][ 338 ],
   alphaCSR[ 135 ][ 339 ],
   alphaCSR[ 135 ][ 340 ],
   alphaCSR[ 135 ][ 341 ],
   alphaCSR[ 135 ][ 342 ],
   alphaCSR[ 135 ][ 343 ],
   alphaCSR[ 135 ][ 344 ],
   alphaCSR[ 135 ][ 345 ],
   alphaCSR[ 135 ][ 346 ],
   alphaCSR[ 135 ][ 347 ],
   alphaCSR[ 135 ][ 348 ],
   alphaCSR[ 135 ][ 349 ],
   alphaCSR[ 135 ][ 350 ],
   alphaCSR[ 135 ][ 351 ],
   alphaCSR[ 135 ][ 352 ],
   alphaCSR[ 135 ][ 353 ],
   alphaCSR[ 135 ][ 354 ],
   alphaCSR[ 135 ][ 355 ],
   alphaCSR[ 135 ][ 356 ],
   alphaCSR[ 135 ][ 357 ],
   alphaCSR[ 135 ][ 358 ],
   alphaCSR[ 135 ][ 359 ],
   alphaCSR[ 135 ][ 360 ],
   alphaCSR[ 135 ][ 361 ],
   alphaCSR[ 135 ][ 362 ],
   alphaCSR[ 135 ][ 363 ],
   alphaCSR[ 135 ][ 364 ],
   alphaCSR[ 135 ][ 365 ],
   alphaCSR[ 135 ][ 366 ],
   alphaCSR[ 135 ][ 367 ],
   alphaCSR[ 135 ][ 368 ],
   alphaCSR[ 135 ][ 369 ],
   alphaCSR[ 135 ][ 370 ],
   alphaCSR[ 135 ][ 371 ],
   alphaCSR[ 135 ][ 372 ],
   alphaCSR[ 135 ][ 373 ],
   alphaCSR[ 135 ][ 374 ],
   alphaCSR[ 135 ][ 375 ],
   alphaCSR[ 135 ][ 376 ],
   alphaCSR[ 135 ][ 377 ],
   alphaCSR[ 135 ][ 378 ],
   alphaCSR[ 135 ][ 379 ],
   alphaCSR[ 135 ][ 380 ],
   alphaCSR[ 135 ][ 381 ],
   alphaCSR[ 135 ][ 382 ],
   alphaCSR[ 135 ][ 383 ],
   alphaCSR[ 136 ][ 0 ],
   alphaCSR[ 136 ][ 1 ],
   alphaCSR[ 136 ][ 2 ],
   alphaCSR[ 136 ][ 3 ],
   alphaCSR[ 136 ][ 4 ],
   alphaCSR[ 136 ][ 5 ],
   alphaCSR[ 136 ][ 6 ],
   alphaCSR[ 136 ][ 7 ],
   alphaCSR[ 136 ][ 8 ],
   alphaCSR[ 136 ][ 9 ],
   alphaCSR[ 136 ][ 10 ],
   alphaCSR[ 136 ][ 11 ],
   alphaCSR[ 136 ][ 12 ],
   alphaCSR[ 136 ][ 13 ],
   alphaCSR[ 136 ][ 14 ],
   alphaCSR[ 136 ][ 15 ],
   alphaCSR[ 136 ][ 16 ],
   alphaCSR[ 136 ][ 17 ],
   alphaCSR[ 136 ][ 18 ],
   alphaCSR[ 136 ][ 19 ],
   alphaCSR[ 136 ][ 20 ],
   alphaCSR[ 136 ][ 21 ],
   alphaCSR[ 136 ][ 22 ],
   alphaCSR[ 136 ][ 23 ],
   alphaCSR[ 136 ][ 24 ],
   alphaCSR[ 136 ][ 25 ],
   alphaCSR[ 136 ][ 26 ],
   alphaCSR[ 136 ][ 27 ],
   alphaCSR[ 136 ][ 28 ],
   alphaCSR[ 136 ][ 29 ],
   alphaCSR[ 136 ][ 30 ],
   alphaCSR[ 136 ][ 31 ],
   alphaCSR[ 136 ][ 32 ],
   alphaCSR[ 136 ][ 33 ],
   alphaCSR[ 136 ][ 34 ],
   alphaCSR[ 136 ][ 35 ],
   alphaCSR[ 136 ][ 36 ],
   alphaCSR[ 136 ][ 37 ],
   alphaCSR[ 136 ][ 38 ],
   alphaCSR[ 136 ][ 39 ],
   alphaCSR[ 136 ][ 40 ],
   alphaCSR[ 136 ][ 41 ],
   alphaCSR[ 136 ][ 42 ],
   alphaCSR[ 136 ][ 43 ],
   alphaCSR[ 136 ][ 44 ],
   alphaCSR[ 136 ][ 45 ],
   alphaCSR[ 136 ][ 46 ],
   alphaCSR[ 136 ][ 47 ],
   alphaCSR[ 136 ][ 48 ],
   alphaCSR[ 136 ][ 49 ],
   alphaCSR[ 136 ][ 50 ],
   alphaCSR[ 136 ][ 51 ],
   alphaCSR[ 136 ][ 52 ],
   alphaCSR[ 136 ][ 53 ],
   alphaCSR[ 136 ][ 54 ],
   alphaCSR[ 136 ][ 55 ],
   alphaCSR[ 136 ][ 56 ],
   alphaCSR[ 136 ][ 57 ],
   alphaCSR[ 136 ][ 58 ],
   alphaCSR[ 136 ][ 59 ],
   alphaCSR[ 136 ][ 60 ],
   alphaCSR[ 136 ][ 61 ],
   alphaCSR[ 136 ][ 62 ],
   alphaCSR[ 136 ][ 63 ],
   alphaCSR[ 136 ][ 64 ],
   alphaCSR[ 136 ][ 65 ],
   alphaCSR[ 136 ][ 66 ],
   alphaCSR[ 136 ][ 67 ],
   alphaCSR[ 136 ][ 68 ],
   alphaCSR[ 136 ][ 69 ],
   alphaCSR[ 136 ][ 70 ],
   alphaCSR[ 136 ][ 71 ],
   alphaCSR[ 136 ][ 72 ],
   alphaCSR[ 136 ][ 73 ],
   alphaCSR[ 136 ][ 74 ],
   alphaCSR[ 136 ][ 75 ],
   alphaCSR[ 136 ][ 76 ],
   alphaCSR[ 136 ][ 77 ],
   alphaCSR[ 136 ][ 78 ],
   alphaCSR[ 136 ][ 79 ],
   alphaCSR[ 136 ][ 80 ],
   alphaCSR[ 136 ][ 81 ],
   alphaCSR[ 136 ][ 82 ],
   alphaCSR[ 136 ][ 83 ],
   alphaCSR[ 136 ][ 84 ],
   alphaCSR[ 136 ][ 85 ],
   alphaCSR[ 136 ][ 86 ],
   alphaCSR[ 136 ][ 87 ],
   alphaCSR[ 136 ][ 88 ],
   alphaCSR[ 136 ][ 89 ],
   alphaCSR[ 136 ][ 90 ],
   alphaCSR[ 136 ][ 91 ],
   alphaCSR[ 136 ][ 92 ],
   alphaCSR[ 136 ][ 93 ],
   alphaCSR[ 136 ][ 94 ],
   alphaCSR[ 136 ][ 95 ],
   alphaCSR[ 136 ][ 96 ],
   alphaCSR[ 136 ][ 97 ],
   alphaCSR[ 136 ][ 98 ],
   alphaCSR[ 136 ][ 99 ],
   alphaCSR[ 136 ][ 100 ],
   alphaCSR[ 136 ][ 101 ],
   alphaCSR[ 136 ][ 102 ],
   alphaCSR[ 136 ][ 103 ],
   alphaCSR[ 136 ][ 104 ],
   alphaCSR[ 136 ][ 105 ],
   alphaCSR[ 136 ][ 106 ],
   alphaCSR[ 136 ][ 107 ],
   alphaCSR[ 136 ][ 108 ],
   alphaCSR[ 136 ][ 109 ],
   alphaCSR[ 136 ][ 110 ],
   alphaCSR[ 136 ][ 111 ],
   alphaCSR[ 136 ][ 112 ],
   alphaCSR[ 136 ][ 113 ],
   alphaCSR[ 136 ][ 114 ],
   alphaCSR[ 136 ][ 115 ],
   alphaCSR[ 136 ][ 116 ],
   alphaCSR[ 136 ][ 117 ],
   alphaCSR[ 136 ][ 118 ],
   alphaCSR[ 136 ][ 119 ],
   alphaCSR[ 136 ][ 120 ],
   alphaCSR[ 136 ][ 121 ],
   alphaCSR[ 136 ][ 122 ],
   alphaCSR[ 136 ][ 123 ],
   alphaCSR[ 136 ][ 124 ],
   alphaCSR[ 136 ][ 125 ],
   alphaCSR[ 136 ][ 126 ],
   alphaCSR[ 136 ][ 127 ],
   alphaCSR[ 136 ][ 128 ],
   alphaCSR[ 136 ][ 129 ],
   alphaCSR[ 136 ][ 130 ],
   alphaCSR[ 136 ][ 131 ],
   alphaCSR[ 136 ][ 132 ],
   alphaCSR[ 136 ][ 133 ],
   alphaCSR[ 136 ][ 134 ],
   alphaCSR[ 136 ][ 135 ],
   alphaCSR[ 136 ][ 136 ],
   alphaCSR[ 136 ][ 137 ],
   alphaCSR[ 136 ][ 138 ],
   alphaCSR[ 136 ][ 139 ],
   alphaCSR[ 136 ][ 140 ],
   alphaCSR[ 136 ][ 141 ],
   alphaCSR[ 136 ][ 142 ],
   alphaCSR[ 136 ][ 143 ],
   alphaCSR[ 136 ][ 144 ],
   alphaCSR[ 136 ][ 145 ],
   alphaCSR[ 136 ][ 146 ],
   alphaCSR[ 136 ][ 147 ],
   alphaCSR[ 136 ][ 148 ],
   alphaCSR[ 136 ][ 149 ],
   alphaCSR[ 136 ][ 150 ],
   alphaCSR[ 136 ][ 151 ],
   alphaCSR[ 136 ][ 152 ],
   alphaCSR[ 136 ][ 153 ],
   alphaCSR[ 136 ][ 154 ],
   alphaCSR[ 136 ][ 155 ],
   alphaCSR[ 136 ][ 156 ],
   alphaCSR[ 136 ][ 157 ],
   alphaCSR[ 136 ][ 158 ],
   alphaCSR[ 136 ][ 159 ],
   alphaCSR[ 136 ][ 160 ],
   alphaCSR[ 136 ][ 161 ],
   alphaCSR[ 136 ][ 162 ],
   alphaCSR[ 136 ][ 163 ],
   alphaCSR[ 136 ][ 164 ],
   alphaCSR[ 136 ][ 165 ],
   alphaCSR[ 136 ][ 166 ],
   alphaCSR[ 136 ][ 167 ],
   alphaCSR[ 136 ][ 168 ],
   alphaCSR[ 136 ][ 169 ],
   alphaCSR[ 136 ][ 170 ],
   alphaCSR[ 136 ][ 171 ],
   alphaCSR[ 136 ][ 172 ],
   alphaCSR[ 136 ][ 173 ],
   alphaCSR[ 136 ][ 174 ],
   alphaCSR[ 136 ][ 175 ],
   alphaCSR[ 136 ][ 176 ],
   alphaCSR[ 136 ][ 177 ],
   alphaCSR[ 136 ][ 178 ],
   alphaCSR[ 136 ][ 179 ],
   alphaCSR[ 136 ][ 180 ],
   alphaCSR[ 136 ][ 181 ],
   alphaCSR[ 136 ][ 182 ],
   alphaCSR[ 136 ][ 183 ],
   alphaCSR[ 136 ][ 184 ],
   alphaCSR[ 136 ][ 185 ],
   alphaCSR[ 136 ][ 186 ],
   alphaCSR[ 136 ][ 187 ],
   alphaCSR[ 136 ][ 188 ],
   alphaCSR[ 136 ][ 189 ],
   alphaCSR[ 136 ][ 190 ],
   alphaCSR[ 136 ][ 191 ],
   alphaCSR[ 136 ][ 192 ],
   alphaCSR[ 136 ][ 193 ],
   alphaCSR[ 136 ][ 194 ],
   alphaCSR[ 136 ][ 195 ],
   alphaCSR[ 136 ][ 196 ],
   alphaCSR[ 136 ][ 197 ],
   alphaCSR[ 136 ][ 198 ],
   alphaCSR[ 136 ][ 199 ],
   alphaCSR[ 136 ][ 200 ],
   alphaCSR[ 136 ][ 201 ],
   alphaCSR[ 136 ][ 202 ],
   alphaCSR[ 136 ][ 203 ],
   alphaCSR[ 136 ][ 204 ],
   alphaCSR[ 136 ][ 205 ],
   alphaCSR[ 136 ][ 206 ],
   alphaCSR[ 136 ][ 207 ],
   alphaCSR[ 136 ][ 208 ],
   alphaCSR[ 136 ][ 209 ],
   alphaCSR[ 136 ][ 210 ],
   alphaCSR[ 136 ][ 211 ],
   alphaCSR[ 136 ][ 212 ],
   alphaCSR[ 136 ][ 213 ],
   alphaCSR[ 136 ][ 214 ],
   alphaCSR[ 136 ][ 215 ],
   alphaCSR[ 136 ][ 216 ],
   alphaCSR[ 136 ][ 217 ],
   alphaCSR[ 136 ][ 218 ],
   alphaCSR[ 136 ][ 219 ],
   alphaCSR[ 136 ][ 220 ],
   alphaCSR[ 136 ][ 221 ],
   alphaCSR[ 136 ][ 222 ],
   alphaCSR[ 136 ][ 223 ],
   alphaCSR[ 136 ][ 224 ],
   alphaCSR[ 136 ][ 225 ],
   alphaCSR[ 136 ][ 226 ],
   alphaCSR[ 136 ][ 227 ],
   alphaCSR[ 136 ][ 228 ],
   alphaCSR[ 136 ][ 229 ],
   alphaCSR[ 136 ][ 230 ],
   alphaCSR[ 136 ][ 231 ],
   alphaCSR[ 136 ][ 232 ],
   alphaCSR[ 136 ][ 233 ],
   alphaCSR[ 136 ][ 234 ],
   alphaCSR[ 136 ][ 235 ],
   alphaCSR[ 136 ][ 236 ],
   alphaCSR[ 136 ][ 237 ],
   alphaCSR[ 136 ][ 238 ],
   alphaCSR[ 136 ][ 239 ],
   alphaCSR[ 136 ][ 240 ],
   alphaCSR[ 136 ][ 241 ],
   alphaCSR[ 136 ][ 242 ],
   alphaCSR[ 136 ][ 243 ],
   alphaCSR[ 136 ][ 244 ],
   alphaCSR[ 136 ][ 245 ],
   alphaCSR[ 136 ][ 246 ],
   alphaCSR[ 136 ][ 247 ],
   alphaCSR[ 136 ][ 248 ],
   alphaCSR[ 136 ][ 249 ],
   alphaCSR[ 136 ][ 250 ],
   alphaCSR[ 136 ][ 251 ],
   alphaCSR[ 136 ][ 252 ],
   alphaCSR[ 136 ][ 253 ],
   alphaCSR[ 136 ][ 254 ],
   alphaCSR[ 136 ][ 255 ],
   alphaCSR[ 136 ][ 256 ],
   alphaCSR[ 136 ][ 257 ],
   alphaCSR[ 136 ][ 258 ],
   alphaCSR[ 136 ][ 259 ],
   alphaCSR[ 136 ][ 260 ],
   alphaCSR[ 136 ][ 261 ],
   alphaCSR[ 136 ][ 262 ],
   alphaCSR[ 136 ][ 263 ],
   alphaCSR[ 136 ][ 264 ],
   alphaCSR[ 136 ][ 265 ],
   alphaCSR[ 136 ][ 266 ],
   alphaCSR[ 136 ][ 267 ],
   alphaCSR[ 136 ][ 268 ],
   alphaCSR[ 136 ][ 269 ],
   alphaCSR[ 136 ][ 270 ],
   alphaCSR[ 136 ][ 271 ],
   alphaCSR[ 136 ][ 272 ],
   alphaCSR[ 136 ][ 273 ],
   alphaCSR[ 136 ][ 274 ],
   alphaCSR[ 136 ][ 275 ],
   alphaCSR[ 136 ][ 276 ],
   alphaCSR[ 136 ][ 277 ],
   alphaCSR[ 136 ][ 278 ],
   alphaCSR[ 136 ][ 279 ],
   alphaCSR[ 136 ][ 280 ],
   alphaCSR[ 136 ][ 281 ],
   alphaCSR[ 136 ][ 282 ],
   alphaCSR[ 136 ][ 283 ],
   alphaCSR[ 136 ][ 284 ],
   alphaCSR[ 136 ][ 285 ],
   alphaCSR[ 136 ][ 286 ],
   alphaCSR[ 136 ][ 287 ],
   alphaCSR[ 136 ][ 288 ],
   alphaCSR[ 136 ][ 289 ],
   alphaCSR[ 136 ][ 290 ],
   alphaCSR[ 136 ][ 291 ],
   alphaCSR[ 136 ][ 292 ],
   alphaCSR[ 136 ][ 293 ],
   alphaCSR[ 136 ][ 294 ],
   alphaCSR[ 136 ][ 295 ],
   alphaCSR[ 136 ][ 296 ],
   alphaCSR[ 136 ][ 297 ],
   alphaCSR[ 136 ][ 298 ],
   alphaCSR[ 136 ][ 299 ],
   alphaCSR[ 136 ][ 300 ],
   alphaCSR[ 136 ][ 301 ],
   alphaCSR[ 136 ][ 302 ],
   alphaCSR[ 136 ][ 303 ],
   alphaCSR[ 136 ][ 304 ],
   alphaCSR[ 136 ][ 305 ],
   alphaCSR[ 136 ][ 306 ],
   alphaCSR[ 136 ][ 307 ],
   alphaCSR[ 136 ][ 308 ],
   alphaCSR[ 136 ][ 309 ],
   alphaCSR[ 136 ][ 310 ],
   alphaCSR[ 136 ][ 311 ],
   alphaCSR[ 136 ][ 312 ],
   alphaCSR[ 136 ][ 313 ],
   alphaCSR[ 136 ][ 314 ],
   alphaCSR[ 136 ][ 315 ],
   alphaCSR[ 136 ][ 316 ],
   alphaCSR[ 136 ][ 317 ],
   alphaCSR[ 136 ][ 318 ],
   alphaCSR[ 136 ][ 319 ],
   alphaCSR[ 136 ][ 320 ],
   alphaCSR[ 136 ][ 321 ],
   alphaCSR[ 136 ][ 322 ],
   alphaCSR[ 136 ][ 323 ],
   alphaCSR[ 136 ][ 324 ],
   alphaCSR[ 136 ][ 325 ],
   alphaCSR[ 136 ][ 326 ],
   alphaCSR[ 136 ][ 327 ],
   alphaCSR[ 136 ][ 328 ],
   alphaCSR[ 136 ][ 329 ],
   alphaCSR[ 136 ][ 330 ],
   alphaCSR[ 136 ][ 331 ],
   alphaCSR[ 136 ][ 332 ],
   alphaCSR[ 136 ][ 333 ],
   alphaCSR[ 136 ][ 334 ],
   alphaCSR[ 136 ][ 335 ],
   alphaCSR[ 136 ][ 336 ],
   alphaCSR[ 136 ][ 337 ],
   alphaCSR[ 136 ][ 338 ],
   alphaCSR[ 136 ][ 339 ],
   alphaCSR[ 136 ][ 340 ],
   alphaCSR[ 136 ][ 341 ],
   alphaCSR[ 136 ][ 342 ],
   alphaCSR[ 136 ][ 343 ],
   alphaCSR[ 136 ][ 344 ],
   alphaCSR[ 136 ][ 345 ],
   alphaCSR[ 136 ][ 346 ],
   alphaCSR[ 136 ][ 347 ],
   alphaCSR[ 136 ][ 348 ],
   alphaCSR[ 136 ][ 349 ],
   alphaCSR[ 136 ][ 350 ],
   alphaCSR[ 136 ][ 351 ],
   alphaCSR[ 136 ][ 352 ],
   alphaCSR[ 136 ][ 353 ],
   alphaCSR[ 136 ][ 354 ],
   alphaCSR[ 136 ][ 355 ],
   alphaCSR[ 136 ][ 356 ],
   alphaCSR[ 136 ][ 357 ],
   alphaCSR[ 136 ][ 358 ],
   alphaCSR[ 136 ][ 359 ],
   alphaCSR[ 136 ][ 360 ],
   alphaCSR[ 136 ][ 361 ],
   alphaCSR[ 136 ][ 362 ],
   alphaCSR[ 136 ][ 363 ],
   alphaCSR[ 136 ][ 364 ],
   alphaCSR[ 136 ][ 365 ],
   alphaCSR[ 136 ][ 366 ],
   alphaCSR[ 136 ][ 367 ],
   alphaCSR[ 136 ][ 368 ],
   alphaCSR[ 136 ][ 369 ],
   alphaCSR[ 136 ][ 370 ],
   alphaCSR[ 136 ][ 371 ],
   alphaCSR[ 136 ][ 372 ],
   alphaCSR[ 136 ][ 373 ],
   alphaCSR[ 136 ][ 374 ],
   alphaCSR[ 136 ][ 375 ],
   alphaCSR[ 136 ][ 376 ],
   alphaCSR[ 136 ][ 377 ],
   alphaCSR[ 136 ][ 378 ],
   alphaCSR[ 136 ][ 379 ],
   alphaCSR[ 136 ][ 380 ],
   alphaCSR[ 136 ][ 381 ],
   alphaCSR[ 136 ][ 382 ],
   alphaCSR[ 136 ][ 383 ],
   alphaCSR[ 137 ][ 0 ],
   alphaCSR[ 137 ][ 1 ],
   alphaCSR[ 137 ][ 2 ],
   alphaCSR[ 137 ][ 3 ],
   alphaCSR[ 137 ][ 4 ],
   alphaCSR[ 137 ][ 5 ],
   alphaCSR[ 137 ][ 6 ],
   alphaCSR[ 137 ][ 7 ],
   alphaCSR[ 137 ][ 8 ],
   alphaCSR[ 137 ][ 9 ],
   alphaCSR[ 137 ][ 10 ],
   alphaCSR[ 137 ][ 11 ],
   alphaCSR[ 137 ][ 12 ],
   alphaCSR[ 137 ][ 13 ],
   alphaCSR[ 137 ][ 14 ],
   alphaCSR[ 137 ][ 15 ],
   alphaCSR[ 137 ][ 16 ],
   alphaCSR[ 137 ][ 17 ],
   alphaCSR[ 137 ][ 18 ],
   alphaCSR[ 137 ][ 19 ],
   alphaCSR[ 137 ][ 20 ],
   alphaCSR[ 137 ][ 21 ],
   alphaCSR[ 137 ][ 22 ],
   alphaCSR[ 137 ][ 23 ],
   alphaCSR[ 137 ][ 24 ],
   alphaCSR[ 137 ][ 25 ],
   alphaCSR[ 137 ][ 26 ],
   alphaCSR[ 137 ][ 27 ],
   alphaCSR[ 137 ][ 28 ],
   alphaCSR[ 137 ][ 29 ],
   alphaCSR[ 137 ][ 30 ],
   alphaCSR[ 137 ][ 31 ],
   alphaCSR[ 137 ][ 32 ],
   alphaCSR[ 137 ][ 33 ],
   alphaCSR[ 137 ][ 34 ],
   alphaCSR[ 137 ][ 35 ],
   alphaCSR[ 137 ][ 36 ],
   alphaCSR[ 137 ][ 37 ],
   alphaCSR[ 137 ][ 38 ],
   alphaCSR[ 137 ][ 39 ],
   alphaCSR[ 137 ][ 40 ],
   alphaCSR[ 137 ][ 41 ],
   alphaCSR[ 137 ][ 42 ],
   alphaCSR[ 137 ][ 43 ],
   alphaCSR[ 137 ][ 44 ],
   alphaCSR[ 137 ][ 45 ],
   alphaCSR[ 137 ][ 46 ],
   alphaCSR[ 137 ][ 47 ],
   alphaCSR[ 137 ][ 48 ],
   alphaCSR[ 137 ][ 49 ],
   alphaCSR[ 137 ][ 50 ],
   alphaCSR[ 137 ][ 51 ],
   alphaCSR[ 137 ][ 52 ],
   alphaCSR[ 137 ][ 53 ],
   alphaCSR[ 137 ][ 54 ],
   alphaCSR[ 137 ][ 55 ],
   alphaCSR[ 137 ][ 56 ],
   alphaCSR[ 137 ][ 57 ],
   alphaCSR[ 137 ][ 58 ],
   alphaCSR[ 137 ][ 59 ],
   alphaCSR[ 137 ][ 60 ],
   alphaCSR[ 137 ][ 61 ],
   alphaCSR[ 137 ][ 62 ],
   alphaCSR[ 137 ][ 63 ],
   alphaCSR[ 137 ][ 64 ],
   alphaCSR[ 137 ][ 65 ],
   alphaCSR[ 137 ][ 66 ],
   alphaCSR[ 137 ][ 67 ],
   alphaCSR[ 137 ][ 68 ],
   alphaCSR[ 137 ][ 69 ],
   alphaCSR[ 137 ][ 70 ],
   alphaCSR[ 137 ][ 71 ],
   alphaCSR[ 137 ][ 72 ],
   alphaCSR[ 137 ][ 73 ],
   alphaCSR[ 137 ][ 74 ],
   alphaCSR[ 137 ][ 75 ],
   alphaCSR[ 137 ][ 76 ],
   alphaCSR[ 137 ][ 77 ],
   alphaCSR[ 137 ][ 78 ],
   alphaCSR[ 137 ][ 79 ],
   alphaCSR[ 137 ][ 80 ],
   alphaCSR[ 137 ][ 81 ],
   alphaCSR[ 137 ][ 82 ],
   alphaCSR[ 137 ][ 83 ],
   alphaCSR[ 137 ][ 84 ],
   alphaCSR[ 137 ][ 85 ],
   alphaCSR[ 137 ][ 86 ],
   alphaCSR[ 137 ][ 87 ],
   alphaCSR[ 137 ][ 88 ],
   alphaCSR[ 137 ][ 89 ],
   alphaCSR[ 137 ][ 90 ],
   alphaCSR[ 137 ][ 91 ],
   alphaCSR[ 137 ][ 92 ],
   alphaCSR[ 137 ][ 93 ],
   alphaCSR[ 137 ][ 94 ],
   alphaCSR[ 137 ][ 95 ],
   alphaCSR[ 137 ][ 96 ],
   alphaCSR[ 137 ][ 97 ],
   alphaCSR[ 137 ][ 98 ],
   alphaCSR[ 137 ][ 99 ],
   alphaCSR[ 137 ][ 100 ],
   alphaCSR[ 137 ][ 101 ],
   alphaCSR[ 137 ][ 102 ],
   alphaCSR[ 137 ][ 103 ],
   alphaCSR[ 137 ][ 104 ],
   alphaCSR[ 137 ][ 105 ],
   alphaCSR[ 137 ][ 106 ],
   alphaCSR[ 137 ][ 107 ],
   alphaCSR[ 137 ][ 108 ],
   alphaCSR[ 137 ][ 109 ],
   alphaCSR[ 137 ][ 110 ],
   alphaCSR[ 137 ][ 111 ],
   alphaCSR[ 137 ][ 112 ],
   alphaCSR[ 137 ][ 113 ],
   alphaCSR[ 137 ][ 114 ],
   alphaCSR[ 137 ][ 115 ],
   alphaCSR[ 137 ][ 116 ],
   alphaCSR[ 137 ][ 117 ],
   alphaCSR[ 137 ][ 118 ],
   alphaCSR[ 137 ][ 119 ],
   alphaCSR[ 137 ][ 120 ],
   alphaCSR[ 137 ][ 121 ],
   alphaCSR[ 137 ][ 122 ],
   alphaCSR[ 137 ][ 123 ],
   alphaCSR[ 137 ][ 124 ],
   alphaCSR[ 137 ][ 125 ],
   alphaCSR[ 137 ][ 126 ],
   alphaCSR[ 137 ][ 127 ],
   alphaCSR[ 137 ][ 128 ],
   alphaCSR[ 137 ][ 129 ],
   alphaCSR[ 137 ][ 130 ],
   alphaCSR[ 137 ][ 131 ],
   alphaCSR[ 137 ][ 132 ],
   alphaCSR[ 137 ][ 133 ],
   alphaCSR[ 137 ][ 134 ],
   alphaCSR[ 137 ][ 135 ],
   alphaCSR[ 137 ][ 136 ],
   alphaCSR[ 137 ][ 137 ],
   alphaCSR[ 137 ][ 138 ],
   alphaCSR[ 137 ][ 139 ],
   alphaCSR[ 137 ][ 140 ],
   alphaCSR[ 137 ][ 141 ],
   alphaCSR[ 137 ][ 142 ],
   alphaCSR[ 137 ][ 143 ],
   alphaCSR[ 137 ][ 144 ],
   alphaCSR[ 137 ][ 145 ],
   alphaCSR[ 137 ][ 146 ],
   alphaCSR[ 137 ][ 147 ],
   alphaCSR[ 137 ][ 148 ],
   alphaCSR[ 137 ][ 149 ],
   alphaCSR[ 137 ][ 150 ],
   alphaCSR[ 137 ][ 151 ],
   alphaCSR[ 137 ][ 152 ],
   alphaCSR[ 137 ][ 153 ],
   alphaCSR[ 137 ][ 154 ],
   alphaCSR[ 137 ][ 155 ],
   alphaCSR[ 137 ][ 156 ],
   alphaCSR[ 137 ][ 157 ],
   alphaCSR[ 137 ][ 158 ],
   alphaCSR[ 137 ][ 159 ],
   alphaCSR[ 137 ][ 160 ],
   alphaCSR[ 137 ][ 161 ],
   alphaCSR[ 137 ][ 162 ],
   alphaCSR[ 137 ][ 163 ],
   alphaCSR[ 137 ][ 164 ],
   alphaCSR[ 137 ][ 165 ],
   alphaCSR[ 137 ][ 166 ],
   alphaCSR[ 137 ][ 167 ],
   alphaCSR[ 137 ][ 168 ],
   alphaCSR[ 137 ][ 169 ],
   alphaCSR[ 137 ][ 170 ],
   alphaCSR[ 137 ][ 171 ],
   alphaCSR[ 137 ][ 172 ],
   alphaCSR[ 137 ][ 173 ],
   alphaCSR[ 137 ][ 174 ],
   alphaCSR[ 137 ][ 175 ],
   alphaCSR[ 137 ][ 176 ],
   alphaCSR[ 137 ][ 177 ],
   alphaCSR[ 137 ][ 178 ],
   alphaCSR[ 137 ][ 179 ],
   alphaCSR[ 137 ][ 180 ],
   alphaCSR[ 137 ][ 181 ],
   alphaCSR[ 137 ][ 182 ],
   alphaCSR[ 137 ][ 183 ],
   alphaCSR[ 137 ][ 184 ],
   alphaCSR[ 137 ][ 185 ],
   alphaCSR[ 137 ][ 186 ],
   alphaCSR[ 137 ][ 187 ],
   alphaCSR[ 137 ][ 188 ],
   alphaCSR[ 137 ][ 189 ],
   alphaCSR[ 137 ][ 190 ],
   alphaCSR[ 137 ][ 191 ],
   alphaCSR[ 137 ][ 192 ],
   alphaCSR[ 137 ][ 193 ],
   alphaCSR[ 137 ][ 194 ],
   alphaCSR[ 137 ][ 195 ],
   alphaCSR[ 137 ][ 196 ],
   alphaCSR[ 137 ][ 197 ],
   alphaCSR[ 137 ][ 198 ],
   alphaCSR[ 137 ][ 199 ],
   alphaCSR[ 137 ][ 200 ],
   alphaCSR[ 137 ][ 201 ],
   alphaCSR[ 137 ][ 202 ],
   alphaCSR[ 137 ][ 203 ],
   alphaCSR[ 137 ][ 204 ],
   alphaCSR[ 137 ][ 205 ],
   alphaCSR[ 137 ][ 206 ],
   alphaCSR[ 137 ][ 207 ],
   alphaCSR[ 137 ][ 208 ],
   alphaCSR[ 137 ][ 209 ],
   alphaCSR[ 137 ][ 210 ],
   alphaCSR[ 137 ][ 211 ],
   alphaCSR[ 137 ][ 212 ],
   alphaCSR[ 137 ][ 213 ],
   alphaCSR[ 137 ][ 214 ],
   alphaCSR[ 137 ][ 215 ],
   alphaCSR[ 137 ][ 216 ],
   alphaCSR[ 137 ][ 217 ],
   alphaCSR[ 137 ][ 218 ],
   alphaCSR[ 137 ][ 219 ],
   alphaCSR[ 137 ][ 220 ],
   alphaCSR[ 137 ][ 221 ],
   alphaCSR[ 137 ][ 222 ],
   alphaCSR[ 137 ][ 223 ],
   alphaCSR[ 137 ][ 224 ],
   alphaCSR[ 137 ][ 225 ],
   alphaCSR[ 137 ][ 226 ],
   alphaCSR[ 137 ][ 227 ],
   alphaCSR[ 137 ][ 228 ],
   alphaCSR[ 137 ][ 229 ],
   alphaCSR[ 137 ][ 230 ],
   alphaCSR[ 137 ][ 231 ],
   alphaCSR[ 137 ][ 232 ],
   alphaCSR[ 137 ][ 233 ],
   alphaCSR[ 137 ][ 234 ],
   alphaCSR[ 137 ][ 235 ],
   alphaCSR[ 137 ][ 236 ],
   alphaCSR[ 137 ][ 237 ],
   alphaCSR[ 137 ][ 238 ],
   alphaCSR[ 137 ][ 239 ],
   alphaCSR[ 137 ][ 240 ],
   alphaCSR[ 137 ][ 241 ],
   alphaCSR[ 137 ][ 242 ],
   alphaCSR[ 137 ][ 243 ],
   alphaCSR[ 137 ][ 244 ],
   alphaCSR[ 137 ][ 245 ],
   alphaCSR[ 137 ][ 246 ],
   alphaCSR[ 137 ][ 247 ],
   alphaCSR[ 137 ][ 248 ],
   alphaCSR[ 137 ][ 249 ],
   alphaCSR[ 137 ][ 250 ],
   alphaCSR[ 137 ][ 251 ],
   alphaCSR[ 137 ][ 252 ],
   alphaCSR[ 137 ][ 253 ],
   alphaCSR[ 137 ][ 254 ],
   alphaCSR[ 137 ][ 255 ],
   alphaCSR[ 137 ][ 256 ],
   alphaCSR[ 137 ][ 257 ],
   alphaCSR[ 137 ][ 258 ],
   alphaCSR[ 137 ][ 259 ],
   alphaCSR[ 137 ][ 260 ],
   alphaCSR[ 137 ][ 261 ],
   alphaCSR[ 137 ][ 262 ],
   alphaCSR[ 137 ][ 263 ],
   alphaCSR[ 137 ][ 264 ],
   alphaCSR[ 137 ][ 265 ],
   alphaCSR[ 137 ][ 266 ],
   alphaCSR[ 137 ][ 267 ],
   alphaCSR[ 137 ][ 268 ],
   alphaCSR[ 137 ][ 269 ],
   alphaCSR[ 137 ][ 270 ],
   alphaCSR[ 137 ][ 271 ],
   alphaCSR[ 137 ][ 272 ],
   alphaCSR[ 137 ][ 273 ],
   alphaCSR[ 137 ][ 274 ],
   alphaCSR[ 137 ][ 275 ],
   alphaCSR[ 137 ][ 276 ],
   alphaCSR[ 137 ][ 277 ],
   alphaCSR[ 137 ][ 278 ],
   alphaCSR[ 137 ][ 279 ],
   alphaCSR[ 137 ][ 280 ],
   alphaCSR[ 137 ][ 281 ],
   alphaCSR[ 137 ][ 282 ],
   alphaCSR[ 137 ][ 283 ],
   alphaCSR[ 137 ][ 284 ],
   alphaCSR[ 137 ][ 285 ],
   alphaCSR[ 137 ][ 286 ],
   alphaCSR[ 137 ][ 287 ],
   alphaCSR[ 137 ][ 288 ],
   alphaCSR[ 137 ][ 289 ],
   alphaCSR[ 137 ][ 290 ],
   alphaCSR[ 137 ][ 291 ],
   alphaCSR[ 137 ][ 292 ],
   alphaCSR[ 137 ][ 293 ],
   alphaCSR[ 137 ][ 294 ],
   alphaCSR[ 137 ][ 295 ],
   alphaCSR[ 137 ][ 296 ],
   alphaCSR[ 137 ][ 297 ],
   alphaCSR[ 137 ][ 298 ],
   alphaCSR[ 137 ][ 299 ],
   alphaCSR[ 137 ][ 300 ],
   alphaCSR[ 137 ][ 301 ],
   alphaCSR[ 137 ][ 302 ],
   alphaCSR[ 137 ][ 303 ],
   alphaCSR[ 137 ][ 304 ],
   alphaCSR[ 137 ][ 305 ],
   alphaCSR[ 137 ][ 306 ],
   alphaCSR[ 137 ][ 307 ],
   alphaCSR[ 137 ][ 308 ],
   alphaCSR[ 137 ][ 309 ],
   alphaCSR[ 137 ][ 310 ],
   alphaCSR[ 137 ][ 311 ],
   alphaCSR[ 137 ][ 312 ],
   alphaCSR[ 137 ][ 313 ],
   alphaCSR[ 137 ][ 314 ],
   alphaCSR[ 137 ][ 315 ],
   alphaCSR[ 137 ][ 316 ],
   alphaCSR[ 137 ][ 317 ],
   alphaCSR[ 137 ][ 318 ],
   alphaCSR[ 137 ][ 319 ],
   alphaCSR[ 137 ][ 320 ],
   alphaCSR[ 137 ][ 321 ],
   alphaCSR[ 137 ][ 322 ],
   alphaCSR[ 137 ][ 323 ],
   alphaCSR[ 137 ][ 324 ],
   alphaCSR[ 137 ][ 325 ],
   alphaCSR[ 137 ][ 326 ],
   alphaCSR[ 137 ][ 327 ],
   alphaCSR[ 137 ][ 328 ],
   alphaCSR[ 137 ][ 329 ],
   alphaCSR[ 137 ][ 330 ],
   alphaCSR[ 137 ][ 331 ],
   alphaCSR[ 137 ][ 332 ],
   alphaCSR[ 137 ][ 333 ],
   alphaCSR[ 137 ][ 334 ],
   alphaCSR[ 137 ][ 335 ],
   alphaCSR[ 137 ][ 336 ],
   alphaCSR[ 137 ][ 337 ],
   alphaCSR[ 137 ][ 338 ],
   alphaCSR[ 137 ][ 339 ],
   alphaCSR[ 137 ][ 340 ],
   alphaCSR[ 137 ][ 341 ],
   alphaCSR[ 137 ][ 342 ],
   alphaCSR[ 137 ][ 343 ],
   alphaCSR[ 137 ][ 344 ],
   alphaCSR[ 137 ][ 345 ],
   alphaCSR[ 137 ][ 346 ],
   alphaCSR[ 137 ][ 347 ],
   alphaCSR[ 137 ][ 348 ],
   alphaCSR[ 137 ][ 349 ],
   alphaCSR[ 137 ][ 350 ],
   alphaCSR[ 137 ][ 351 ],
   alphaCSR[ 137 ][ 352 ],
   alphaCSR[ 137 ][ 353 ],
   alphaCSR[ 137 ][ 354 ],
   alphaCSR[ 137 ][ 355 ],
   alphaCSR[ 137 ][ 356 ],
   alphaCSR[ 137 ][ 357 ],
   alphaCSR[ 137 ][ 358 ],
   alphaCSR[ 137 ][ 359 ],
   alphaCSR[ 137 ][ 360 ],
   alphaCSR[ 137 ][ 361 ],
   alphaCSR[ 137 ][ 362 ],
   alphaCSR[ 137 ][ 363 ],
   alphaCSR[ 137 ][ 364 ],
   alphaCSR[ 137 ][ 365 ],
   alphaCSR[ 137 ][ 366 ],
   alphaCSR[ 137 ][ 367 ],
   alphaCSR[ 137 ][ 368 ],
   alphaCSR[ 137 ][ 369 ],
   alphaCSR[ 137 ][ 370 ],
   alphaCSR[ 137 ][ 371 ],
   alphaCSR[ 137 ][ 372 ],
   alphaCSR[ 137 ][ 373 ],
   alphaCSR[ 137 ][ 374 ],
   alphaCSR[ 137 ][ 375 ],
   alphaCSR[ 137 ][ 376 ],
   alphaCSR[ 137 ][ 377 ],
   alphaCSR[ 137 ][ 378 ],
   alphaCSR[ 137 ][ 379 ],
   alphaCSR[ 137 ][ 380 ],
   alphaCSR[ 137 ][ 381 ],
   alphaCSR[ 137 ][ 382 ],
   alphaCSR[ 137 ][ 383 ],
   alphaCSR[ 138 ][ 0 ],
   alphaCSR[ 138 ][ 1 ],
   alphaCSR[ 138 ][ 2 ],
   alphaCSR[ 138 ][ 3 ],
   alphaCSR[ 138 ][ 4 ],
   alphaCSR[ 138 ][ 5 ],
   alphaCSR[ 138 ][ 6 ],
   alphaCSR[ 138 ][ 7 ],
   alphaCSR[ 138 ][ 8 ],
   alphaCSR[ 138 ][ 9 ],
   alphaCSR[ 138 ][ 10 ],
   alphaCSR[ 138 ][ 11 ],
   alphaCSR[ 138 ][ 12 ],
   alphaCSR[ 138 ][ 13 ],
   alphaCSR[ 138 ][ 14 ],
   alphaCSR[ 138 ][ 15 ],
   alphaCSR[ 138 ][ 16 ],
   alphaCSR[ 138 ][ 17 ],
   alphaCSR[ 138 ][ 18 ],
   alphaCSR[ 138 ][ 19 ],
   alphaCSR[ 138 ][ 20 ],
   alphaCSR[ 138 ][ 21 ],
   alphaCSR[ 138 ][ 22 ],
   alphaCSR[ 138 ][ 23 ],
   alphaCSR[ 138 ][ 24 ],
   alphaCSR[ 138 ][ 25 ],
   alphaCSR[ 138 ][ 26 ],
   alphaCSR[ 138 ][ 27 ],
   alphaCSR[ 138 ][ 28 ],
   alphaCSR[ 138 ][ 29 ],
   alphaCSR[ 138 ][ 30 ],
   alphaCSR[ 138 ][ 31 ],
   alphaCSR[ 138 ][ 32 ],
   alphaCSR[ 138 ][ 33 ],
   alphaCSR[ 138 ][ 34 ],
   alphaCSR[ 138 ][ 35 ],
   alphaCSR[ 138 ][ 36 ],
   alphaCSR[ 138 ][ 37 ],
   alphaCSR[ 138 ][ 38 ],
   alphaCSR[ 138 ][ 39 ],
   alphaCSR[ 138 ][ 40 ],
   alphaCSR[ 138 ][ 41 ],
   alphaCSR[ 138 ][ 42 ],
   alphaCSR[ 138 ][ 43 ],
   alphaCSR[ 138 ][ 44 ],
   alphaCSR[ 138 ][ 45 ],
   alphaCSR[ 138 ][ 46 ],
   alphaCSR[ 138 ][ 47 ],
   alphaCSR[ 138 ][ 48 ],
   alphaCSR[ 138 ][ 49 ],
   alphaCSR[ 138 ][ 50 ],
   alphaCSR[ 138 ][ 51 ],
   alphaCSR[ 138 ][ 52 ],
   alphaCSR[ 138 ][ 53 ],
   alphaCSR[ 138 ][ 54 ],
   alphaCSR[ 138 ][ 55 ],
   alphaCSR[ 138 ][ 56 ],
   alphaCSR[ 138 ][ 57 ],
   alphaCSR[ 138 ][ 58 ],
   alphaCSR[ 138 ][ 59 ],
   alphaCSR[ 138 ][ 60 ],
   alphaCSR[ 138 ][ 61 ],
   alphaCSR[ 138 ][ 62 ],
   alphaCSR[ 138 ][ 63 ],
   alphaCSR[ 138 ][ 64 ],
   alphaCSR[ 138 ][ 65 ],
   alphaCSR[ 138 ][ 66 ],
   alphaCSR[ 138 ][ 67 ],
   alphaCSR[ 138 ][ 68 ],
   alphaCSR[ 138 ][ 69 ],
   alphaCSR[ 138 ][ 70 ],
   alphaCSR[ 138 ][ 71 ],
   alphaCSR[ 138 ][ 72 ],
   alphaCSR[ 138 ][ 73 ],
   alphaCSR[ 138 ][ 74 ],
   alphaCSR[ 138 ][ 75 ],
   alphaCSR[ 138 ][ 76 ],
   alphaCSR[ 138 ][ 77 ],
   alphaCSR[ 138 ][ 78 ],
   alphaCSR[ 138 ][ 79 ],
   alphaCSR[ 138 ][ 80 ],
   alphaCSR[ 138 ][ 81 ],
   alphaCSR[ 138 ][ 82 ],
   alphaCSR[ 138 ][ 83 ],
   alphaCSR[ 138 ][ 84 ],
   alphaCSR[ 138 ][ 85 ],
   alphaCSR[ 138 ][ 86 ],
   alphaCSR[ 138 ][ 87 ],
   alphaCSR[ 138 ][ 88 ],
   alphaCSR[ 138 ][ 89 ],
   alphaCSR[ 138 ][ 90 ],
   alphaCSR[ 138 ][ 91 ],
   alphaCSR[ 138 ][ 92 ],
   alphaCSR[ 138 ][ 93 ],
   alphaCSR[ 138 ][ 94 ],
   alphaCSR[ 138 ][ 95 ],
   alphaCSR[ 138 ][ 96 ],
   alphaCSR[ 138 ][ 97 ],
   alphaCSR[ 138 ][ 98 ],
   alphaCSR[ 138 ][ 99 ],
   alphaCSR[ 138 ][ 100 ],
   alphaCSR[ 138 ][ 101 ],
   alphaCSR[ 138 ][ 102 ],
   alphaCSR[ 138 ][ 103 ],
   alphaCSR[ 138 ][ 104 ],
   alphaCSR[ 138 ][ 105 ],
   alphaCSR[ 138 ][ 106 ],
   alphaCSR[ 138 ][ 107 ],
   alphaCSR[ 138 ][ 108 ],
   alphaCSR[ 138 ][ 109 ],
   alphaCSR[ 138 ][ 110 ],
   alphaCSR[ 138 ][ 111 ],
   alphaCSR[ 138 ][ 112 ],
   alphaCSR[ 138 ][ 113 ],
   alphaCSR[ 138 ][ 114 ],
   alphaCSR[ 138 ][ 115 ],
   alphaCSR[ 138 ][ 116 ],
   alphaCSR[ 138 ][ 117 ],
   alphaCSR[ 138 ][ 118 ],
   alphaCSR[ 138 ][ 119 ],
   alphaCSR[ 138 ][ 120 ],
   alphaCSR[ 138 ][ 121 ],
   alphaCSR[ 138 ][ 122 ],
   alphaCSR[ 138 ][ 123 ],
   alphaCSR[ 138 ][ 124 ],
   alphaCSR[ 138 ][ 125 ],
   alphaCSR[ 138 ][ 126 ],
   alphaCSR[ 138 ][ 127 ],
   alphaCSR[ 138 ][ 128 ],
   alphaCSR[ 138 ][ 129 ],
   alphaCSR[ 138 ][ 130 ],
   alphaCSR[ 138 ][ 131 ],
   alphaCSR[ 138 ][ 132 ],
   alphaCSR[ 138 ][ 133 ],
   alphaCSR[ 138 ][ 134 ],
   alphaCSR[ 138 ][ 135 ],
   alphaCSR[ 138 ][ 136 ],
   alphaCSR[ 138 ][ 137 ],
   alphaCSR[ 138 ][ 138 ],
   alphaCSR[ 138 ][ 139 ],
   alphaCSR[ 138 ][ 140 ],
   alphaCSR[ 138 ][ 141 ],
   alphaCSR[ 138 ][ 142 ],
   alphaCSR[ 138 ][ 143 ],
   alphaCSR[ 138 ][ 144 ],
   alphaCSR[ 138 ][ 145 ],
   alphaCSR[ 138 ][ 146 ],
   alphaCSR[ 138 ][ 147 ],
   alphaCSR[ 138 ][ 148 ],
   alphaCSR[ 138 ][ 149 ],
   alphaCSR[ 138 ][ 150 ],
   alphaCSR[ 138 ][ 151 ],
   alphaCSR[ 138 ][ 152 ],
   alphaCSR[ 138 ][ 153 ],
   alphaCSR[ 138 ][ 154 ],
   alphaCSR[ 138 ][ 155 ],
   alphaCSR[ 138 ][ 156 ],
   alphaCSR[ 138 ][ 157 ],
   alphaCSR[ 138 ][ 158 ],
   alphaCSR[ 138 ][ 159 ],
   alphaCSR[ 138 ][ 160 ],
   alphaCSR[ 138 ][ 161 ],
   alphaCSR[ 138 ][ 162 ],
   alphaCSR[ 138 ][ 163 ],
   alphaCSR[ 138 ][ 164 ],
   alphaCSR[ 138 ][ 165 ],
   alphaCSR[ 138 ][ 166 ],
   alphaCSR[ 138 ][ 167 ],
   alphaCSR[ 138 ][ 168 ],
   alphaCSR[ 138 ][ 169 ],
   alphaCSR[ 138 ][ 170 ],
   alphaCSR[ 138 ][ 171 ],
   alphaCSR[ 138 ][ 172 ],
   alphaCSR[ 138 ][ 173 ],
   alphaCSR[ 138 ][ 174 ],
   alphaCSR[ 138 ][ 175 ],
   alphaCSR[ 138 ][ 176 ],
   alphaCSR[ 138 ][ 177 ],
   alphaCSR[ 138 ][ 178 ],
   alphaCSR[ 138 ][ 179 ],
   alphaCSR[ 138 ][ 180 ],
   alphaCSR[ 138 ][ 181 ],
   alphaCSR[ 138 ][ 182 ],
   alphaCSR[ 138 ][ 183 ],
   alphaCSR[ 138 ][ 184 ],
   alphaCSR[ 138 ][ 185 ],
   alphaCSR[ 138 ][ 186 ],
   alphaCSR[ 138 ][ 187 ],
   alphaCSR[ 138 ][ 188 ],
   alphaCSR[ 138 ][ 189 ],
   alphaCSR[ 138 ][ 190 ],
   alphaCSR[ 138 ][ 191 ],
   alphaCSR[ 138 ][ 192 ],
   alphaCSR[ 138 ][ 193 ],
   alphaCSR[ 138 ][ 194 ],
   alphaCSR[ 138 ][ 195 ],
   alphaCSR[ 138 ][ 196 ],
   alphaCSR[ 138 ][ 197 ],
   alphaCSR[ 138 ][ 198 ],
   alphaCSR[ 138 ][ 199 ],
   alphaCSR[ 138 ][ 200 ],
   alphaCSR[ 138 ][ 201 ],
   alphaCSR[ 138 ][ 202 ],
   alphaCSR[ 138 ][ 203 ],
   alphaCSR[ 138 ][ 204 ],
   alphaCSR[ 138 ][ 205 ],
   alphaCSR[ 138 ][ 206 ],
   alphaCSR[ 138 ][ 207 ],
   alphaCSR[ 138 ][ 208 ],
   alphaCSR[ 138 ][ 209 ],
   alphaCSR[ 138 ][ 210 ],
   alphaCSR[ 138 ][ 211 ],
   alphaCSR[ 138 ][ 212 ],
   alphaCSR[ 138 ][ 213 ],
   alphaCSR[ 138 ][ 214 ],
   alphaCSR[ 138 ][ 215 ],
   alphaCSR[ 138 ][ 216 ],
   alphaCSR[ 138 ][ 217 ],
   alphaCSR[ 138 ][ 218 ],
   alphaCSR[ 138 ][ 219 ],
   alphaCSR[ 138 ][ 220 ],
   alphaCSR[ 138 ][ 221 ],
   alphaCSR[ 138 ][ 222 ],
   alphaCSR[ 138 ][ 223 ],
   alphaCSR[ 138 ][ 224 ],
   alphaCSR[ 138 ][ 225 ],
   alphaCSR[ 138 ][ 226 ],
   alphaCSR[ 138 ][ 227 ],
   alphaCSR[ 138 ][ 228 ],
   alphaCSR[ 138 ][ 229 ],
   alphaCSR[ 138 ][ 230 ],
   alphaCSR[ 138 ][ 231 ],
   alphaCSR[ 138 ][ 232 ],
   alphaCSR[ 138 ][ 233 ],
   alphaCSR[ 138 ][ 234 ],
   alphaCSR[ 138 ][ 235 ],
   alphaCSR[ 138 ][ 236 ],
   alphaCSR[ 138 ][ 237 ],
   alphaCSR[ 138 ][ 238 ],
   alphaCSR[ 138 ][ 239 ],
   alphaCSR[ 138 ][ 240 ],
   alphaCSR[ 138 ][ 241 ],
   alphaCSR[ 138 ][ 242 ],
   alphaCSR[ 138 ][ 243 ],
   alphaCSR[ 138 ][ 244 ],
   alphaCSR[ 138 ][ 245 ],
   alphaCSR[ 138 ][ 246 ],
   alphaCSR[ 138 ][ 247 ],
   alphaCSR[ 138 ][ 248 ],
   alphaCSR[ 138 ][ 249 ],
   alphaCSR[ 138 ][ 250 ],
   alphaCSR[ 138 ][ 251 ],
   alphaCSR[ 138 ][ 252 ],
   alphaCSR[ 138 ][ 253 ],
   alphaCSR[ 138 ][ 254 ],
   alphaCSR[ 138 ][ 255 ],
   alphaCSR[ 138 ][ 256 ],
   alphaCSR[ 138 ][ 257 ],
   alphaCSR[ 138 ][ 258 ],
   alphaCSR[ 138 ][ 259 ],
   alphaCSR[ 138 ][ 260 ],
   alphaCSR[ 138 ][ 261 ],
   alphaCSR[ 138 ][ 262 ],
   alphaCSR[ 138 ][ 263 ],
   alphaCSR[ 138 ][ 264 ],
   alphaCSR[ 138 ][ 265 ],
   alphaCSR[ 138 ][ 266 ],
   alphaCSR[ 138 ][ 267 ],
   alphaCSR[ 138 ][ 268 ],
   alphaCSR[ 138 ][ 269 ],
   alphaCSR[ 138 ][ 270 ],
   alphaCSR[ 138 ][ 271 ],
   alphaCSR[ 138 ][ 272 ],
   alphaCSR[ 138 ][ 273 ],
   alphaCSR[ 138 ][ 274 ],
   alphaCSR[ 138 ][ 275 ],
   alphaCSR[ 138 ][ 276 ],
   alphaCSR[ 138 ][ 277 ],
   alphaCSR[ 138 ][ 278 ],
   alphaCSR[ 138 ][ 279 ],
   alphaCSR[ 138 ][ 280 ],
   alphaCSR[ 138 ][ 281 ],
   alphaCSR[ 138 ][ 282 ],
   alphaCSR[ 138 ][ 283 ],
   alphaCSR[ 138 ][ 284 ],
   alphaCSR[ 138 ][ 285 ],
   alphaCSR[ 138 ][ 286 ],
   alphaCSR[ 138 ][ 287 ],
   alphaCSR[ 138 ][ 288 ],
   alphaCSR[ 138 ][ 289 ],
   alphaCSR[ 138 ][ 290 ],
   alphaCSR[ 138 ][ 291 ],
   alphaCSR[ 138 ][ 292 ],
   alphaCSR[ 138 ][ 293 ],
   alphaCSR[ 138 ][ 294 ],
   alphaCSR[ 138 ][ 295 ],
   alphaCSR[ 138 ][ 296 ],
   alphaCSR[ 138 ][ 297 ],
   alphaCSR[ 138 ][ 298 ],
   alphaCSR[ 138 ][ 299 ],
   alphaCSR[ 138 ][ 300 ],
   alphaCSR[ 138 ][ 301 ],
   alphaCSR[ 138 ][ 302 ],
   alphaCSR[ 138 ][ 303 ],
   alphaCSR[ 138 ][ 304 ],
   alphaCSR[ 138 ][ 305 ],
   alphaCSR[ 138 ][ 306 ],
   alphaCSR[ 138 ][ 307 ],
   alphaCSR[ 138 ][ 308 ],
   alphaCSR[ 138 ][ 309 ],
   alphaCSR[ 138 ][ 310 ],
   alphaCSR[ 138 ][ 311 ],
   alphaCSR[ 138 ][ 312 ],
   alphaCSR[ 138 ][ 313 ],
   alphaCSR[ 138 ][ 314 ],
   alphaCSR[ 138 ][ 315 ],
   alphaCSR[ 138 ][ 316 ],
   alphaCSR[ 138 ][ 317 ],
   alphaCSR[ 138 ][ 318 ],
   alphaCSR[ 138 ][ 319 ],
   alphaCSR[ 138 ][ 320 ],
   alphaCSR[ 138 ][ 321 ],
   alphaCSR[ 138 ][ 322 ],
   alphaCSR[ 138 ][ 323 ],
   alphaCSR[ 138 ][ 324 ],
   alphaCSR[ 138 ][ 325 ],
   alphaCSR[ 138 ][ 326 ],
   alphaCSR[ 138 ][ 327 ],
   alphaCSR[ 138 ][ 328 ],
   alphaCSR[ 138 ][ 329 ],
   alphaCSR[ 138 ][ 330 ],
   alphaCSR[ 138 ][ 331 ],
   alphaCSR[ 138 ][ 332 ],
   alphaCSR[ 138 ][ 333 ],
   alphaCSR[ 138 ][ 334 ],
   alphaCSR[ 138 ][ 335 ],
   alphaCSR[ 138 ][ 336 ],
   alphaCSR[ 138 ][ 337 ],
   alphaCSR[ 138 ][ 338 ],
   alphaCSR[ 138 ][ 339 ],
   alphaCSR[ 138 ][ 340 ],
   alphaCSR[ 138 ][ 341 ],
   alphaCSR[ 138 ][ 342 ],
   alphaCSR[ 138 ][ 343 ],
   alphaCSR[ 138 ][ 344 ],
   alphaCSR[ 138 ][ 345 ],
   alphaCSR[ 138 ][ 346 ],
   alphaCSR[ 138 ][ 347 ],
   alphaCSR[ 138 ][ 348 ],
   alphaCSR[ 138 ][ 349 ],
   alphaCSR[ 138 ][ 350 ],
   alphaCSR[ 138 ][ 351 ],
   alphaCSR[ 138 ][ 352 ],
   alphaCSR[ 138 ][ 353 ],
   alphaCSR[ 138 ][ 354 ],
   alphaCSR[ 138 ][ 355 ],
   alphaCSR[ 138 ][ 356 ],
   alphaCSR[ 138 ][ 357 ],
   alphaCSR[ 138 ][ 358 ],
   alphaCSR[ 138 ][ 359 ],
   alphaCSR[ 138 ][ 360 ],
   alphaCSR[ 138 ][ 361 ],
   alphaCSR[ 138 ][ 362 ],
   alphaCSR[ 138 ][ 363 ],
   alphaCSR[ 138 ][ 364 ],
   alphaCSR[ 138 ][ 365 ],
   alphaCSR[ 138 ][ 366 ],
   alphaCSR[ 138 ][ 367 ],
   alphaCSR[ 138 ][ 368 ],
   alphaCSR[ 138 ][ 369 ],
   alphaCSR[ 138 ][ 370 ],
   alphaCSR[ 138 ][ 371 ],
   alphaCSR[ 138 ][ 372 ],
   alphaCSR[ 138 ][ 373 ],
   alphaCSR[ 138 ][ 374 ],
   alphaCSR[ 138 ][ 375 ],
   alphaCSR[ 138 ][ 376 ],
   alphaCSR[ 138 ][ 377 ],
   alphaCSR[ 138 ][ 378 ],
   alphaCSR[ 138 ][ 379 ],
   alphaCSR[ 138 ][ 380 ],
   alphaCSR[ 138 ][ 381 ],
   alphaCSR[ 138 ][ 382 ],
   alphaCSR[ 138 ][ 383 ],
   alphaCSR[ 139 ][ 0 ],
   alphaCSR[ 139 ][ 1 ],
   alphaCSR[ 139 ][ 2 ],
   alphaCSR[ 139 ][ 3 ],
   alphaCSR[ 139 ][ 4 ],
   alphaCSR[ 139 ][ 5 ],
   alphaCSR[ 139 ][ 6 ],
   alphaCSR[ 139 ][ 7 ],
   alphaCSR[ 139 ][ 8 ],
   alphaCSR[ 139 ][ 9 ],
   alphaCSR[ 139 ][ 10 ],
   alphaCSR[ 139 ][ 11 ],
   alphaCSR[ 139 ][ 12 ],
   alphaCSR[ 139 ][ 13 ],
   alphaCSR[ 139 ][ 14 ],
   alphaCSR[ 139 ][ 15 ],
   alphaCSR[ 139 ][ 16 ],
   alphaCSR[ 139 ][ 17 ],
   alphaCSR[ 139 ][ 18 ],
   alphaCSR[ 139 ][ 19 ],
   alphaCSR[ 139 ][ 20 ],
   alphaCSR[ 139 ][ 21 ],
   alphaCSR[ 139 ][ 22 ],
   alphaCSR[ 139 ][ 23 ],
   alphaCSR[ 139 ][ 24 ],
   alphaCSR[ 139 ][ 25 ],
   alphaCSR[ 139 ][ 26 ],
   alphaCSR[ 139 ][ 27 ],
   alphaCSR[ 139 ][ 28 ],
   alphaCSR[ 139 ][ 29 ],
   alphaCSR[ 139 ][ 30 ],
   alphaCSR[ 139 ][ 31 ],
   alphaCSR[ 139 ][ 32 ],
   alphaCSR[ 139 ][ 33 ],
   alphaCSR[ 139 ][ 34 ],
   alphaCSR[ 139 ][ 35 ],
   alphaCSR[ 139 ][ 36 ],
   alphaCSR[ 139 ][ 37 ],
   alphaCSR[ 139 ][ 38 ],
   alphaCSR[ 139 ][ 39 ],
   alphaCSR[ 139 ][ 40 ],
   alphaCSR[ 139 ][ 41 ],
   alphaCSR[ 139 ][ 42 ],
   alphaCSR[ 139 ][ 43 ],
   alphaCSR[ 139 ][ 44 ],
   alphaCSR[ 139 ][ 45 ],
   alphaCSR[ 139 ][ 46 ],
   alphaCSR[ 139 ][ 47 ],
   alphaCSR[ 139 ][ 48 ],
   alphaCSR[ 139 ][ 49 ],
   alphaCSR[ 139 ][ 50 ],
   alphaCSR[ 139 ][ 51 ],
   alphaCSR[ 139 ][ 52 ],
   alphaCSR[ 139 ][ 53 ],
   alphaCSR[ 139 ][ 54 ],
   alphaCSR[ 139 ][ 55 ],
   alphaCSR[ 139 ][ 56 ],
   alphaCSR[ 139 ][ 57 ],
   alphaCSR[ 139 ][ 58 ],
   alphaCSR[ 139 ][ 59 ],
   alphaCSR[ 139 ][ 60 ],
   alphaCSR[ 139 ][ 61 ],
   alphaCSR[ 139 ][ 62 ],
   alphaCSR[ 139 ][ 63 ],
   alphaCSR[ 139 ][ 64 ],
   alphaCSR[ 139 ][ 65 ],
   alphaCSR[ 139 ][ 66 ],
   alphaCSR[ 139 ][ 67 ],
   alphaCSR[ 139 ][ 68 ],
   alphaCSR[ 139 ][ 69 ],
   alphaCSR[ 139 ][ 70 ],
   alphaCSR[ 139 ][ 71 ],
   alphaCSR[ 139 ][ 72 ],
   alphaCSR[ 139 ][ 73 ],
   alphaCSR[ 139 ][ 74 ],
   alphaCSR[ 139 ][ 75 ],
   alphaCSR[ 139 ][ 76 ],
   alphaCSR[ 139 ][ 77 ],
   alphaCSR[ 139 ][ 78 ],
   alphaCSR[ 139 ][ 79 ],
   alphaCSR[ 139 ][ 80 ],
   alphaCSR[ 139 ][ 81 ],
   alphaCSR[ 139 ][ 82 ],
   alphaCSR[ 139 ][ 83 ],
   alphaCSR[ 139 ][ 84 ],
   alphaCSR[ 139 ][ 85 ],
   alphaCSR[ 139 ][ 86 ],
   alphaCSR[ 139 ][ 87 ],
   alphaCSR[ 139 ][ 88 ],
   alphaCSR[ 139 ][ 89 ],
   alphaCSR[ 139 ][ 90 ],
   alphaCSR[ 139 ][ 91 ],
   alphaCSR[ 139 ][ 92 ],
   alphaCSR[ 139 ][ 93 ],
   alphaCSR[ 139 ][ 94 ],
   alphaCSR[ 139 ][ 95 ],
   alphaCSR[ 139 ][ 96 ],
   alphaCSR[ 139 ][ 97 ],
   alphaCSR[ 139 ][ 98 ],
   alphaCSR[ 139 ][ 99 ],
   alphaCSR[ 139 ][ 100 ],
   alphaCSR[ 139 ][ 101 ],
   alphaCSR[ 139 ][ 102 ],
   alphaCSR[ 139 ][ 103 ],
   alphaCSR[ 139 ][ 104 ],
   alphaCSR[ 139 ][ 105 ],
   alphaCSR[ 139 ][ 106 ],
   alphaCSR[ 139 ][ 107 ],
   alphaCSR[ 139 ][ 108 ],
   alphaCSR[ 139 ][ 109 ],
   alphaCSR[ 139 ][ 110 ],
   alphaCSR[ 139 ][ 111 ],
   alphaCSR[ 139 ][ 112 ],
   alphaCSR[ 139 ][ 113 ],
   alphaCSR[ 139 ][ 114 ],
   alphaCSR[ 139 ][ 115 ],
   alphaCSR[ 139 ][ 116 ],
   alphaCSR[ 139 ][ 117 ],
   alphaCSR[ 139 ][ 118 ],
   alphaCSR[ 139 ][ 119 ],
   alphaCSR[ 139 ][ 120 ],
   alphaCSR[ 139 ][ 121 ],
   alphaCSR[ 139 ][ 122 ],
   alphaCSR[ 139 ][ 123 ],
   alphaCSR[ 139 ][ 124 ],
   alphaCSR[ 139 ][ 125 ],
   alphaCSR[ 139 ][ 126 ],
   alphaCSR[ 139 ][ 127 ],
   alphaCSR[ 139 ][ 128 ],
   alphaCSR[ 139 ][ 129 ],
   alphaCSR[ 139 ][ 130 ],
   alphaCSR[ 139 ][ 131 ],
   alphaCSR[ 139 ][ 132 ],
   alphaCSR[ 139 ][ 133 ],
   alphaCSR[ 139 ][ 134 ],
   alphaCSR[ 139 ][ 135 ],
   alphaCSR[ 139 ][ 136 ],
   alphaCSR[ 139 ][ 137 ],
   alphaCSR[ 139 ][ 138 ],
   alphaCSR[ 139 ][ 139 ],
   alphaCSR[ 139 ][ 140 ],
   alphaCSR[ 139 ][ 141 ],
   alphaCSR[ 139 ][ 142 ],
   alphaCSR[ 139 ][ 143 ],
   alphaCSR[ 139 ][ 144 ],
   alphaCSR[ 139 ][ 145 ],
   alphaCSR[ 139 ][ 146 ],
   alphaCSR[ 139 ][ 147 ],
   alphaCSR[ 139 ][ 148 ],
   alphaCSR[ 139 ][ 149 ],
   alphaCSR[ 139 ][ 150 ],
   alphaCSR[ 139 ][ 151 ],
   alphaCSR[ 139 ][ 152 ],
   alphaCSR[ 139 ][ 153 ],
   alphaCSR[ 139 ][ 154 ],
   alphaCSR[ 139 ][ 155 ],
   alphaCSR[ 139 ][ 156 ],
   alphaCSR[ 139 ][ 157 ],
   alphaCSR[ 139 ][ 158 ],
   alphaCSR[ 139 ][ 159 ],
   alphaCSR[ 139 ][ 160 ],
   alphaCSR[ 139 ][ 161 ],
   alphaCSR[ 139 ][ 162 ],
   alphaCSR[ 139 ][ 163 ],
   alphaCSR[ 139 ][ 164 ],
   alphaCSR[ 139 ][ 165 ],
   alphaCSR[ 139 ][ 166 ],
   alphaCSR[ 139 ][ 167 ],
   alphaCSR[ 139 ][ 168 ],
   alphaCSR[ 139 ][ 169 ],
   alphaCSR[ 139 ][ 170 ],
   alphaCSR[ 139 ][ 171 ],
   alphaCSR[ 139 ][ 172 ],
   alphaCSR[ 139 ][ 173 ],
   alphaCSR[ 139 ][ 174 ],
   alphaCSR[ 139 ][ 175 ],
   alphaCSR[ 139 ][ 176 ],
   alphaCSR[ 139 ][ 177 ],
   alphaCSR[ 139 ][ 178 ],
   alphaCSR[ 139 ][ 179 ],
   alphaCSR[ 139 ][ 180 ],
   alphaCSR[ 139 ][ 181 ],
   alphaCSR[ 139 ][ 182 ],
   alphaCSR[ 139 ][ 183 ],
   alphaCSR[ 139 ][ 184 ],
   alphaCSR[ 139 ][ 185 ],
   alphaCSR[ 139 ][ 186 ],
   alphaCSR[ 139 ][ 187 ],
   alphaCSR[ 139 ][ 188 ],
   alphaCSR[ 139 ][ 189 ],
   alphaCSR[ 139 ][ 190 ],
   alphaCSR[ 139 ][ 191 ],
   alphaCSR[ 139 ][ 192 ],
   alphaCSR[ 139 ][ 193 ],
   alphaCSR[ 139 ][ 194 ],
   alphaCSR[ 139 ][ 195 ],
   alphaCSR[ 139 ][ 196 ],
   alphaCSR[ 139 ][ 197 ],
   alphaCSR[ 139 ][ 198 ],
   alphaCSR[ 139 ][ 199 ],
   alphaCSR[ 139 ][ 200 ],
   alphaCSR[ 139 ][ 201 ],
   alphaCSR[ 139 ][ 202 ],
   alphaCSR[ 139 ][ 203 ],
   alphaCSR[ 139 ][ 204 ],
   alphaCSR[ 139 ][ 205 ],
   alphaCSR[ 139 ][ 206 ],
   alphaCSR[ 139 ][ 207 ],
   alphaCSR[ 139 ][ 208 ],
   alphaCSR[ 139 ][ 209 ],
   alphaCSR[ 139 ][ 210 ],
   alphaCSR[ 139 ][ 211 ],
   alphaCSR[ 139 ][ 212 ],
   alphaCSR[ 139 ][ 213 ],
   alphaCSR[ 139 ][ 214 ],
   alphaCSR[ 139 ][ 215 ],
   alphaCSR[ 139 ][ 216 ],
   alphaCSR[ 139 ][ 217 ],
   alphaCSR[ 139 ][ 218 ],
   alphaCSR[ 139 ][ 219 ],
   alphaCSR[ 139 ][ 220 ],
   alphaCSR[ 139 ][ 221 ],
   alphaCSR[ 139 ][ 222 ],
   alphaCSR[ 139 ][ 223 ],
   alphaCSR[ 139 ][ 224 ],
   alphaCSR[ 139 ][ 225 ],
   alphaCSR[ 139 ][ 226 ],
   alphaCSR[ 139 ][ 227 ],
   alphaCSR[ 139 ][ 228 ],
   alphaCSR[ 139 ][ 229 ],
   alphaCSR[ 139 ][ 230 ],
   alphaCSR[ 139 ][ 231 ],
   alphaCSR[ 139 ][ 232 ],
   alphaCSR[ 139 ][ 233 ],
   alphaCSR[ 139 ][ 234 ],
   alphaCSR[ 139 ][ 235 ],
   alphaCSR[ 139 ][ 236 ],
   alphaCSR[ 139 ][ 237 ],
   alphaCSR[ 139 ][ 238 ],
   alphaCSR[ 139 ][ 239 ],
   alphaCSR[ 139 ][ 240 ],
   alphaCSR[ 139 ][ 241 ],
   alphaCSR[ 139 ][ 242 ],
   alphaCSR[ 139 ][ 243 ],
   alphaCSR[ 139 ][ 244 ],
   alphaCSR[ 139 ][ 245 ],
   alphaCSR[ 139 ][ 246 ],
   alphaCSR[ 139 ][ 247 ],
   alphaCSR[ 139 ][ 248 ],
   alphaCSR[ 139 ][ 249 ],
   alphaCSR[ 139 ][ 250 ],
   alphaCSR[ 139 ][ 251 ],
   alphaCSR[ 139 ][ 252 ],
   alphaCSR[ 139 ][ 253 ],
   alphaCSR[ 139 ][ 254 ],
   alphaCSR[ 139 ][ 255 ],
   alphaCSR[ 139 ][ 256 ],
   alphaCSR[ 139 ][ 257 ],
   alphaCSR[ 139 ][ 258 ],
   alphaCSR[ 139 ][ 259 ],
   alphaCSR[ 139 ][ 260 ],
   alphaCSR[ 139 ][ 261 ],
   alphaCSR[ 139 ][ 262 ],
   alphaCSR[ 139 ][ 263 ],
   alphaCSR[ 139 ][ 264 ],
   alphaCSR[ 139 ][ 265 ],
   alphaCSR[ 139 ][ 266 ],
   alphaCSR[ 139 ][ 267 ],
   alphaCSR[ 139 ][ 268 ],
   alphaCSR[ 139 ][ 269 ],
   alphaCSR[ 139 ][ 270 ],
   alphaCSR[ 139 ][ 271 ],
   alphaCSR[ 139 ][ 272 ],
   alphaCSR[ 139 ][ 273 ],
   alphaCSR[ 139 ][ 274 ],
   alphaCSR[ 139 ][ 275 ],
   alphaCSR[ 139 ][ 276 ],
   alphaCSR[ 139 ][ 277 ],
   alphaCSR[ 139 ][ 278 ],
   alphaCSR[ 139 ][ 279 ],
   alphaCSR[ 139 ][ 280 ],
   alphaCSR[ 139 ][ 281 ],
   alphaCSR[ 139 ][ 282 ],
   alphaCSR[ 139 ][ 283 ],
   alphaCSR[ 139 ][ 284 ],
   alphaCSR[ 139 ][ 285 ],
   alphaCSR[ 139 ][ 286 ],
   alphaCSR[ 139 ][ 287 ],
   alphaCSR[ 139 ][ 288 ],
   alphaCSR[ 139 ][ 289 ],
   alphaCSR[ 139 ][ 290 ],
   alphaCSR[ 139 ][ 291 ],
   alphaCSR[ 139 ][ 292 ],
   alphaCSR[ 139 ][ 293 ],
   alphaCSR[ 139 ][ 294 ],
   alphaCSR[ 139 ][ 295 ],
   alphaCSR[ 139 ][ 296 ],
   alphaCSR[ 139 ][ 297 ],
   alphaCSR[ 139 ][ 298 ],
   alphaCSR[ 139 ][ 299 ],
   alphaCSR[ 139 ][ 300 ],
   alphaCSR[ 139 ][ 301 ],
   alphaCSR[ 139 ][ 302 ],
   alphaCSR[ 139 ][ 303 ],
   alphaCSR[ 139 ][ 304 ],
   alphaCSR[ 139 ][ 305 ],
   alphaCSR[ 139 ][ 306 ],
   alphaCSR[ 139 ][ 307 ],
   alphaCSR[ 139 ][ 308 ],
   alphaCSR[ 139 ][ 309 ],
   alphaCSR[ 139 ][ 310 ],
   alphaCSR[ 139 ][ 311 ],
   alphaCSR[ 139 ][ 312 ],
   alphaCSR[ 139 ][ 313 ],
   alphaCSR[ 139 ][ 314 ],
   alphaCSR[ 139 ][ 315 ],
   alphaCSR[ 139 ][ 316 ],
   alphaCSR[ 139 ][ 317 ],
   alphaCSR[ 139 ][ 318 ],
   alphaCSR[ 139 ][ 319 ],
   alphaCSR[ 139 ][ 320 ],
   alphaCSR[ 139 ][ 321 ],
   alphaCSR[ 139 ][ 322 ],
   alphaCSR[ 139 ][ 323 ],
   alphaCSR[ 139 ][ 324 ],
   alphaCSR[ 139 ][ 325 ],
   alphaCSR[ 139 ][ 326 ],
   alphaCSR[ 139 ][ 327 ],
   alphaCSR[ 139 ][ 328 ],
   alphaCSR[ 139 ][ 329 ],
   alphaCSR[ 139 ][ 330 ],
   alphaCSR[ 139 ][ 331 ],
   alphaCSR[ 139 ][ 332 ],
   alphaCSR[ 139 ][ 333 ],
   alphaCSR[ 139 ][ 334 ],
   alphaCSR[ 139 ][ 335 ],
   alphaCSR[ 139 ][ 336 ],
   alphaCSR[ 139 ][ 337 ],
   alphaCSR[ 139 ][ 338 ],
   alphaCSR[ 139 ][ 339 ],
   alphaCSR[ 139 ][ 340 ],
   alphaCSR[ 139 ][ 341 ],
   alphaCSR[ 139 ][ 342 ],
   alphaCSR[ 139 ][ 343 ],
   alphaCSR[ 139 ][ 344 ],
   alphaCSR[ 139 ][ 345 ],
   alphaCSR[ 139 ][ 346 ],
   alphaCSR[ 139 ][ 347 ],
   alphaCSR[ 139 ][ 348 ],
   alphaCSR[ 139 ][ 349 ],
   alphaCSR[ 139 ][ 350 ],
   alphaCSR[ 139 ][ 351 ],
   alphaCSR[ 139 ][ 352 ],
   alphaCSR[ 139 ][ 353 ],
   alphaCSR[ 139 ][ 354 ],
   alphaCSR[ 139 ][ 355 ],
   alphaCSR[ 139 ][ 356 ],
   alphaCSR[ 139 ][ 357 ],
   alphaCSR[ 139 ][ 358 ],
   alphaCSR[ 139 ][ 359 ],
   alphaCSR[ 139 ][ 360 ],
   alphaCSR[ 139 ][ 361 ],
   alphaCSR[ 139 ][ 362 ],
   alphaCSR[ 139 ][ 363 ],
   alphaCSR[ 139 ][ 364 ],
   alphaCSR[ 139 ][ 365 ],
   alphaCSR[ 139 ][ 366 ],
   alphaCSR[ 139 ][ 367 ],
   alphaCSR[ 139 ][ 368 ],
   alphaCSR[ 139 ][ 369 ],
   alphaCSR[ 139 ][ 370 ],
   alphaCSR[ 139 ][ 371 ],
   alphaCSR[ 139 ][ 372 ],
   alphaCSR[ 139 ][ 373 ],
   alphaCSR[ 139 ][ 374 ],
   alphaCSR[ 139 ][ 375 ],
   alphaCSR[ 139 ][ 376 ],
   alphaCSR[ 139 ][ 377 ],
   alphaCSR[ 139 ][ 378 ],
   alphaCSR[ 139 ][ 379 ],
   alphaCSR[ 139 ][ 380 ],
   alphaCSR[ 139 ][ 381 ],
   alphaCSR[ 139 ][ 382 ],
   alphaCSR[ 139 ][ 383 ],
   alphaCSR[ 140 ][ 0 ],
   alphaCSR[ 140 ][ 1 ],
   alphaCSR[ 140 ][ 2 ],
   alphaCSR[ 140 ][ 3 ],
   alphaCSR[ 140 ][ 4 ],
   alphaCSR[ 140 ][ 5 ],
   alphaCSR[ 140 ][ 6 ],
   alphaCSR[ 140 ][ 7 ],
   alphaCSR[ 140 ][ 8 ],
   alphaCSR[ 140 ][ 9 ],
   alphaCSR[ 140 ][ 10 ],
   alphaCSR[ 140 ][ 11 ],
   alphaCSR[ 140 ][ 12 ],
   alphaCSR[ 140 ][ 13 ],
   alphaCSR[ 140 ][ 14 ],
   alphaCSR[ 140 ][ 15 ],
   alphaCSR[ 140 ][ 16 ],
   alphaCSR[ 140 ][ 17 ],
   alphaCSR[ 140 ][ 18 ],
   alphaCSR[ 140 ][ 19 ],
   alphaCSR[ 140 ][ 20 ],
   alphaCSR[ 140 ][ 21 ],
   alphaCSR[ 140 ][ 22 ],
   alphaCSR[ 140 ][ 23 ],
   alphaCSR[ 140 ][ 24 ],
   alphaCSR[ 140 ][ 25 ],
   alphaCSR[ 140 ][ 26 ],
   alphaCSR[ 140 ][ 27 ],
   alphaCSR[ 140 ][ 28 ],
   alphaCSR[ 140 ][ 29 ],
   alphaCSR[ 140 ][ 30 ],
   alphaCSR[ 140 ][ 31 ],
   alphaCSR[ 140 ][ 32 ],
   alphaCSR[ 140 ][ 33 ],
   alphaCSR[ 140 ][ 34 ],
   alphaCSR[ 140 ][ 35 ],
   alphaCSR[ 140 ][ 36 ],
   alphaCSR[ 140 ][ 37 ],
   alphaCSR[ 140 ][ 38 ],
   alphaCSR[ 140 ][ 39 ],
   alphaCSR[ 140 ][ 40 ],
   alphaCSR[ 140 ][ 41 ],
   alphaCSR[ 140 ][ 42 ],
   alphaCSR[ 140 ][ 43 ],
   alphaCSR[ 140 ][ 44 ],
   alphaCSR[ 140 ][ 45 ],
   alphaCSR[ 140 ][ 46 ],
   alphaCSR[ 140 ][ 47 ],
   alphaCSR[ 140 ][ 48 ],
   alphaCSR[ 140 ][ 49 ],
   alphaCSR[ 140 ][ 50 ],
   alphaCSR[ 140 ][ 51 ],
   alphaCSR[ 140 ][ 52 ],
   alphaCSR[ 140 ][ 53 ],
   alphaCSR[ 140 ][ 54 ],
   alphaCSR[ 140 ][ 55 ],
   alphaCSR[ 140 ][ 56 ],
   alphaCSR[ 140 ][ 57 ],
   alphaCSR[ 140 ][ 58 ],
   alphaCSR[ 140 ][ 59 ],
   alphaCSR[ 140 ][ 60 ],
   alphaCSR[ 140 ][ 61 ],
   alphaCSR[ 140 ][ 62 ],
   alphaCSR[ 140 ][ 63 ],
   alphaCSR[ 140 ][ 64 ],
   alphaCSR[ 140 ][ 65 ],
   alphaCSR[ 140 ][ 66 ],
   alphaCSR[ 140 ][ 67 ],
   alphaCSR[ 140 ][ 68 ],
   alphaCSR[ 140 ][ 69 ],
   alphaCSR[ 140 ][ 70 ],
   alphaCSR[ 140 ][ 71 ],
   alphaCSR[ 140 ][ 72 ],
   alphaCSR[ 140 ][ 73 ],
   alphaCSR[ 140 ][ 74 ],
   alphaCSR[ 140 ][ 75 ],
   alphaCSR[ 140 ][ 76 ],
   alphaCSR[ 140 ][ 77 ],
   alphaCSR[ 140 ][ 78 ],
   alphaCSR[ 140 ][ 79 ],
   alphaCSR[ 140 ][ 80 ],
   alphaCSR[ 140 ][ 81 ],
   alphaCSR[ 140 ][ 82 ],
   alphaCSR[ 140 ][ 83 ],
   alphaCSR[ 140 ][ 84 ],
   alphaCSR[ 140 ][ 85 ],
   alphaCSR[ 140 ][ 86 ],
   alphaCSR[ 140 ][ 87 ],
   alphaCSR[ 140 ][ 88 ],
   alphaCSR[ 140 ][ 89 ],
   alphaCSR[ 140 ][ 90 ],
   alphaCSR[ 140 ][ 91 ],
   alphaCSR[ 140 ][ 92 ],
   alphaCSR[ 140 ][ 93 ],
   alphaCSR[ 140 ][ 94 ],
   alphaCSR[ 140 ][ 95 ],
   alphaCSR[ 140 ][ 96 ],
   alphaCSR[ 140 ][ 97 ],
   alphaCSR[ 140 ][ 98 ],
   alphaCSR[ 140 ][ 99 ],
   alphaCSR[ 140 ][ 100 ],
   alphaCSR[ 140 ][ 101 ],
   alphaCSR[ 140 ][ 102 ],
   alphaCSR[ 140 ][ 103 ],
   alphaCSR[ 140 ][ 104 ],
   alphaCSR[ 140 ][ 105 ],
   alphaCSR[ 140 ][ 106 ],
   alphaCSR[ 140 ][ 107 ],
   alphaCSR[ 140 ][ 108 ],
   alphaCSR[ 140 ][ 109 ],
   alphaCSR[ 140 ][ 110 ],
   alphaCSR[ 140 ][ 111 ],
   alphaCSR[ 140 ][ 112 ],
   alphaCSR[ 140 ][ 113 ],
   alphaCSR[ 140 ][ 114 ],
   alphaCSR[ 140 ][ 115 ],
   alphaCSR[ 140 ][ 116 ],
   alphaCSR[ 140 ][ 117 ],
   alphaCSR[ 140 ][ 118 ],
   alphaCSR[ 140 ][ 119 ],
   alphaCSR[ 140 ][ 120 ],
   alphaCSR[ 140 ][ 121 ],
   alphaCSR[ 140 ][ 122 ],
   alphaCSR[ 140 ][ 123 ],
   alphaCSR[ 140 ][ 124 ],
   alphaCSR[ 140 ][ 125 ],
   alphaCSR[ 140 ][ 126 ],
   alphaCSR[ 140 ][ 127 ],
   alphaCSR[ 140 ][ 128 ],
   alphaCSR[ 140 ][ 129 ],
   alphaCSR[ 140 ][ 130 ],
   alphaCSR[ 140 ][ 131 ],
   alphaCSR[ 140 ][ 132 ],
   alphaCSR[ 140 ][ 133 ],
   alphaCSR[ 140 ][ 134 ],
   alphaCSR[ 140 ][ 135 ],
   alphaCSR[ 140 ][ 136 ],
   alphaCSR[ 140 ][ 137 ],
   alphaCSR[ 140 ][ 138 ],
   alphaCSR[ 140 ][ 139 ],
   alphaCSR[ 140 ][ 140 ],
   alphaCSR[ 140 ][ 141 ],
   alphaCSR[ 140 ][ 142 ],
   alphaCSR[ 140 ][ 143 ],
   alphaCSR[ 140 ][ 144 ],
   alphaCSR[ 140 ][ 145 ],
   alphaCSR[ 140 ][ 146 ],
   alphaCSR[ 140 ][ 147 ],
   alphaCSR[ 140 ][ 148 ],
   alphaCSR[ 140 ][ 149 ],
   alphaCSR[ 140 ][ 150 ],
   alphaCSR[ 140 ][ 151 ],
   alphaCSR[ 140 ][ 152 ],
   alphaCSR[ 140 ][ 153 ],
   alphaCSR[ 140 ][ 154 ],
   alphaCSR[ 140 ][ 155 ],
   alphaCSR[ 140 ][ 156 ],
   alphaCSR[ 140 ][ 157 ],
   alphaCSR[ 140 ][ 158 ],
   alphaCSR[ 140 ][ 159 ],
   alphaCSR[ 140 ][ 160 ],
   alphaCSR[ 140 ][ 161 ],
   alphaCSR[ 140 ][ 162 ],
   alphaCSR[ 140 ][ 163 ],
   alphaCSR[ 140 ][ 164 ],
   alphaCSR[ 140 ][ 165 ],
   alphaCSR[ 140 ][ 166 ],
   alphaCSR[ 140 ][ 167 ],
   alphaCSR[ 140 ][ 168 ],
   alphaCSR[ 140 ][ 169 ],
   alphaCSR[ 140 ][ 170 ],
   alphaCSR[ 140 ][ 171 ],
   alphaCSR[ 140 ][ 172 ],
   alphaCSR[ 140 ][ 173 ],
   alphaCSR[ 140 ][ 174 ],
   alphaCSR[ 140 ][ 175 ],
   alphaCSR[ 140 ][ 176 ],
   alphaCSR[ 140 ][ 177 ],
   alphaCSR[ 140 ][ 178 ],
   alphaCSR[ 140 ][ 179 ],
   alphaCSR[ 140 ][ 180 ],
   alphaCSR[ 140 ][ 181 ],
   alphaCSR[ 140 ][ 182 ],
   alphaCSR[ 140 ][ 183 ],
   alphaCSR[ 140 ][ 184 ],
   alphaCSR[ 140 ][ 185 ],
   alphaCSR[ 140 ][ 186 ],
   alphaCSR[ 140 ][ 187 ],
   alphaCSR[ 140 ][ 188 ],
   alphaCSR[ 140 ][ 189 ],
   alphaCSR[ 140 ][ 190 ],
   alphaCSR[ 140 ][ 191 ],
   alphaCSR[ 140 ][ 192 ],
   alphaCSR[ 140 ][ 193 ],
   alphaCSR[ 140 ][ 194 ],
   alphaCSR[ 140 ][ 195 ],
   alphaCSR[ 140 ][ 196 ],
   alphaCSR[ 140 ][ 197 ],
   alphaCSR[ 140 ][ 198 ],
   alphaCSR[ 140 ][ 199 ],
   alphaCSR[ 140 ][ 200 ],
   alphaCSR[ 140 ][ 201 ],
   alphaCSR[ 140 ][ 202 ],
   alphaCSR[ 140 ][ 203 ],
   alphaCSR[ 140 ][ 204 ],
   alphaCSR[ 140 ][ 205 ],
   alphaCSR[ 140 ][ 206 ],
   alphaCSR[ 140 ][ 207 ],
   alphaCSR[ 140 ][ 208 ],
   alphaCSR[ 140 ][ 209 ],
   alphaCSR[ 140 ][ 210 ],
   alphaCSR[ 140 ][ 211 ],
   alphaCSR[ 140 ][ 212 ],
   alphaCSR[ 140 ][ 213 ],
   alphaCSR[ 140 ][ 214 ],
   alphaCSR[ 140 ][ 215 ],
   alphaCSR[ 140 ][ 216 ],
   alphaCSR[ 140 ][ 217 ],
   alphaCSR[ 140 ][ 218 ],
   alphaCSR[ 140 ][ 219 ],
   alphaCSR[ 140 ][ 220 ],
   alphaCSR[ 140 ][ 221 ],
   alphaCSR[ 140 ][ 222 ],
   alphaCSR[ 140 ][ 223 ],
   alphaCSR[ 140 ][ 224 ],
   alphaCSR[ 140 ][ 225 ],
   alphaCSR[ 140 ][ 226 ],
   alphaCSR[ 140 ][ 227 ],
   alphaCSR[ 140 ][ 228 ],
   alphaCSR[ 140 ][ 229 ],
   alphaCSR[ 140 ][ 230 ],
   alphaCSR[ 140 ][ 231 ],
   alphaCSR[ 140 ][ 232 ],
   alphaCSR[ 140 ][ 233 ],
   alphaCSR[ 140 ][ 234 ],
   alphaCSR[ 140 ][ 235 ],
   alphaCSR[ 140 ][ 236 ],
   alphaCSR[ 140 ][ 237 ],
   alphaCSR[ 140 ][ 238 ],
   alphaCSR[ 140 ][ 239 ],
   alphaCSR[ 140 ][ 240 ],
   alphaCSR[ 140 ][ 241 ],
   alphaCSR[ 140 ][ 242 ],
   alphaCSR[ 140 ][ 243 ],
   alphaCSR[ 140 ][ 244 ],
   alphaCSR[ 140 ][ 245 ],
   alphaCSR[ 140 ][ 246 ],
   alphaCSR[ 140 ][ 247 ],
   alphaCSR[ 140 ][ 248 ],
   alphaCSR[ 140 ][ 249 ],
   alphaCSR[ 140 ][ 250 ],
   alphaCSR[ 140 ][ 251 ],
   alphaCSR[ 140 ][ 252 ],
   alphaCSR[ 140 ][ 253 ],
   alphaCSR[ 140 ][ 254 ],
   alphaCSR[ 140 ][ 255 ],
   alphaCSR[ 140 ][ 256 ],
   alphaCSR[ 140 ][ 257 ],
   alphaCSR[ 140 ][ 258 ],
   alphaCSR[ 140 ][ 259 ],
   alphaCSR[ 140 ][ 260 ],
   alphaCSR[ 140 ][ 261 ],
   alphaCSR[ 140 ][ 262 ],
   alphaCSR[ 140 ][ 263 ],
   alphaCSR[ 140 ][ 264 ],
   alphaCSR[ 140 ][ 265 ],
   alphaCSR[ 140 ][ 266 ],
   alphaCSR[ 140 ][ 267 ],
   alphaCSR[ 140 ][ 268 ],
   alphaCSR[ 140 ][ 269 ],
   alphaCSR[ 140 ][ 270 ],
   alphaCSR[ 140 ][ 271 ],
   alphaCSR[ 140 ][ 272 ],
   alphaCSR[ 140 ][ 273 ],
   alphaCSR[ 140 ][ 274 ],
   alphaCSR[ 140 ][ 275 ],
   alphaCSR[ 140 ][ 276 ],
   alphaCSR[ 140 ][ 277 ],
   alphaCSR[ 140 ][ 278 ],
   alphaCSR[ 140 ][ 279 ],
   alphaCSR[ 140 ][ 280 ],
   alphaCSR[ 140 ][ 281 ],
   alphaCSR[ 140 ][ 282 ],
   alphaCSR[ 140 ][ 283 ],
   alphaCSR[ 140 ][ 284 ],
   alphaCSR[ 140 ][ 285 ],
   alphaCSR[ 140 ][ 286 ],
   alphaCSR[ 140 ][ 287 ],
   alphaCSR[ 140 ][ 288 ],
   alphaCSR[ 140 ][ 289 ],
   alphaCSR[ 140 ][ 290 ],
   alphaCSR[ 140 ][ 291 ],
   alphaCSR[ 140 ][ 292 ],
   alphaCSR[ 140 ][ 293 ],
   alphaCSR[ 140 ][ 294 ],
   alphaCSR[ 140 ][ 295 ],
   alphaCSR[ 140 ][ 296 ],
   alphaCSR[ 140 ][ 297 ],
   alphaCSR[ 140 ][ 298 ],
   alphaCSR[ 140 ][ 299 ],
   alphaCSR[ 140 ][ 300 ],
   alphaCSR[ 140 ][ 301 ],
   alphaCSR[ 140 ][ 302 ],
   alphaCSR[ 140 ][ 303 ],
   alphaCSR[ 140 ][ 304 ],
   alphaCSR[ 140 ][ 305 ],
   alphaCSR[ 140 ][ 306 ],
   alphaCSR[ 140 ][ 307 ],
   alphaCSR[ 140 ][ 308 ],
   alphaCSR[ 140 ][ 309 ],
   alphaCSR[ 140 ][ 310 ],
   alphaCSR[ 140 ][ 311 ],
   alphaCSR[ 140 ][ 312 ],
   alphaCSR[ 140 ][ 313 ],
   alphaCSR[ 140 ][ 314 ],
   alphaCSR[ 140 ][ 315 ],
   alphaCSR[ 140 ][ 316 ],
   alphaCSR[ 140 ][ 317 ],
   alphaCSR[ 140 ][ 318 ],
   alphaCSR[ 140 ][ 319 ],
   alphaCSR[ 140 ][ 320 ],
   alphaCSR[ 140 ][ 321 ],
   alphaCSR[ 140 ][ 322 ],
   alphaCSR[ 140 ][ 323 ],
   alphaCSR[ 140 ][ 324 ],
   alphaCSR[ 140 ][ 325 ],
   alphaCSR[ 140 ][ 326 ],
   alphaCSR[ 140 ][ 327 ],
   alphaCSR[ 140 ][ 328 ],
   alphaCSR[ 140 ][ 329 ],
   alphaCSR[ 140 ][ 330 ],
   alphaCSR[ 140 ][ 331 ],
   alphaCSR[ 140 ][ 332 ],
   alphaCSR[ 140 ][ 333 ],
   alphaCSR[ 140 ][ 334 ],
   alphaCSR[ 140 ][ 335 ],
   alphaCSR[ 140 ][ 336 ],
   alphaCSR[ 140 ][ 337 ],
   alphaCSR[ 140 ][ 338 ],
   alphaCSR[ 140 ][ 339 ],
   alphaCSR[ 140 ][ 340 ],
   alphaCSR[ 140 ][ 341 ],
   alphaCSR[ 140 ][ 342 ],
   alphaCSR[ 140 ][ 343 ],
   alphaCSR[ 140 ][ 344 ],
   alphaCSR[ 140 ][ 345 ],
   alphaCSR[ 140 ][ 346 ],
   alphaCSR[ 140 ][ 347 ],
   alphaCSR[ 140 ][ 348 ],
   alphaCSR[ 140 ][ 349 ],
   alphaCSR[ 140 ][ 350 ],
   alphaCSR[ 140 ][ 351 ],
   alphaCSR[ 140 ][ 352 ],
   alphaCSR[ 140 ][ 353 ],
   alphaCSR[ 140 ][ 354 ],
   alphaCSR[ 140 ][ 355 ],
   alphaCSR[ 140 ][ 356 ],
   alphaCSR[ 140 ][ 357 ],
   alphaCSR[ 140 ][ 358 ],
   alphaCSR[ 140 ][ 359 ],
   alphaCSR[ 140 ][ 360 ],
   alphaCSR[ 140 ][ 361 ],
   alphaCSR[ 140 ][ 362 ],
   alphaCSR[ 140 ][ 363 ],
   alphaCSR[ 140 ][ 364 ],
   alphaCSR[ 140 ][ 365 ],
   alphaCSR[ 140 ][ 366 ],
   alphaCSR[ 140 ][ 367 ],
   alphaCSR[ 140 ][ 368 ],
   alphaCSR[ 140 ][ 369 ],
   alphaCSR[ 140 ][ 370 ],
   alphaCSR[ 140 ][ 371 ],
   alphaCSR[ 140 ][ 372 ],
   alphaCSR[ 140 ][ 373 ],
   alphaCSR[ 140 ][ 374 ],
   alphaCSR[ 140 ][ 375 ],
   alphaCSR[ 140 ][ 376 ],
   alphaCSR[ 140 ][ 377 ],
   alphaCSR[ 140 ][ 378 ],
   alphaCSR[ 140 ][ 379 ],
   alphaCSR[ 140 ][ 380 ],
   alphaCSR[ 140 ][ 381 ],
   alphaCSR[ 140 ][ 382 ],
   alphaCSR[ 140 ][ 383 ],
   alphaCSR[ 141 ][ 0 ],
   alphaCSR[ 141 ][ 1 ],
   alphaCSR[ 141 ][ 2 ],
   alphaCSR[ 141 ][ 3 ],
   alphaCSR[ 141 ][ 4 ],
   alphaCSR[ 141 ][ 5 ],
   alphaCSR[ 141 ][ 6 ],
   alphaCSR[ 141 ][ 7 ],
   alphaCSR[ 141 ][ 8 ],
   alphaCSR[ 141 ][ 9 ],
   alphaCSR[ 141 ][ 10 ],
   alphaCSR[ 141 ][ 11 ],
   alphaCSR[ 141 ][ 12 ],
   alphaCSR[ 141 ][ 13 ],
   alphaCSR[ 141 ][ 14 ],
   alphaCSR[ 141 ][ 15 ],
   alphaCSR[ 141 ][ 16 ],
   alphaCSR[ 141 ][ 17 ],
   alphaCSR[ 141 ][ 18 ],
   alphaCSR[ 141 ][ 19 ],
   alphaCSR[ 141 ][ 20 ],
   alphaCSR[ 141 ][ 21 ],
   alphaCSR[ 141 ][ 22 ],
   alphaCSR[ 141 ][ 23 ],
   alphaCSR[ 141 ][ 24 ],
   alphaCSR[ 141 ][ 25 ],
   alphaCSR[ 141 ][ 26 ],
   alphaCSR[ 141 ][ 27 ],
   alphaCSR[ 141 ][ 28 ],
   alphaCSR[ 141 ][ 29 ],
   alphaCSR[ 141 ][ 30 ],
   alphaCSR[ 141 ][ 31 ],
   alphaCSR[ 141 ][ 32 ],
   alphaCSR[ 141 ][ 33 ],
   alphaCSR[ 141 ][ 34 ],
   alphaCSR[ 141 ][ 35 ],
   alphaCSR[ 141 ][ 36 ],
   alphaCSR[ 141 ][ 37 ],
   alphaCSR[ 141 ][ 38 ],
   alphaCSR[ 141 ][ 39 ],
   alphaCSR[ 141 ][ 40 ],
   alphaCSR[ 141 ][ 41 ],
   alphaCSR[ 141 ][ 42 ],
   alphaCSR[ 141 ][ 43 ],
   alphaCSR[ 141 ][ 44 ],
   alphaCSR[ 141 ][ 45 ],
   alphaCSR[ 141 ][ 46 ],
   alphaCSR[ 141 ][ 47 ],
   alphaCSR[ 141 ][ 48 ],
   alphaCSR[ 141 ][ 49 ],
   alphaCSR[ 141 ][ 50 ],
   alphaCSR[ 141 ][ 51 ],
   alphaCSR[ 141 ][ 52 ],
   alphaCSR[ 141 ][ 53 ],
   alphaCSR[ 141 ][ 54 ],
   alphaCSR[ 141 ][ 55 ],
   alphaCSR[ 141 ][ 56 ],
   alphaCSR[ 141 ][ 57 ],
   alphaCSR[ 141 ][ 58 ],
   alphaCSR[ 141 ][ 59 ],
   alphaCSR[ 141 ][ 60 ],
   alphaCSR[ 141 ][ 61 ],
   alphaCSR[ 141 ][ 62 ],
   alphaCSR[ 141 ][ 63 ],
   alphaCSR[ 141 ][ 64 ],
   alphaCSR[ 141 ][ 65 ],
   alphaCSR[ 141 ][ 66 ],
   alphaCSR[ 141 ][ 67 ],
   alphaCSR[ 141 ][ 68 ],
   alphaCSR[ 141 ][ 69 ],
   alphaCSR[ 141 ][ 70 ],
   alphaCSR[ 141 ][ 71 ],
   alphaCSR[ 141 ][ 72 ],
   alphaCSR[ 141 ][ 73 ],
   alphaCSR[ 141 ][ 74 ],
   alphaCSR[ 141 ][ 75 ],
   alphaCSR[ 141 ][ 76 ],
   alphaCSR[ 141 ][ 77 ],
   alphaCSR[ 141 ][ 78 ],
   alphaCSR[ 141 ][ 79 ],
   alphaCSR[ 141 ][ 80 ],
   alphaCSR[ 141 ][ 81 ],
   alphaCSR[ 141 ][ 82 ],
   alphaCSR[ 141 ][ 83 ],
   alphaCSR[ 141 ][ 84 ],
   alphaCSR[ 141 ][ 85 ],
   alphaCSR[ 141 ][ 86 ],
   alphaCSR[ 141 ][ 87 ],
   alphaCSR[ 141 ][ 88 ],
   alphaCSR[ 141 ][ 89 ],
   alphaCSR[ 141 ][ 90 ],
   alphaCSR[ 141 ][ 91 ],
   alphaCSR[ 141 ][ 92 ],
   alphaCSR[ 141 ][ 93 ],
   alphaCSR[ 141 ][ 94 ],
   alphaCSR[ 141 ][ 95 ],
   alphaCSR[ 141 ][ 96 ],
   alphaCSR[ 141 ][ 97 ],
   alphaCSR[ 141 ][ 98 ],
   alphaCSR[ 141 ][ 99 ],
   alphaCSR[ 141 ][ 100 ],
   alphaCSR[ 141 ][ 101 ],
   alphaCSR[ 141 ][ 102 ],
   alphaCSR[ 141 ][ 103 ],
   alphaCSR[ 141 ][ 104 ],
   alphaCSR[ 141 ][ 105 ],
   alphaCSR[ 141 ][ 106 ],
   alphaCSR[ 141 ][ 107 ],
   alphaCSR[ 141 ][ 108 ],
   alphaCSR[ 141 ][ 109 ],
   alphaCSR[ 141 ][ 110 ],
   alphaCSR[ 141 ][ 111 ],
   alphaCSR[ 141 ][ 112 ],
   alphaCSR[ 141 ][ 113 ],
   alphaCSR[ 141 ][ 114 ],
   alphaCSR[ 141 ][ 115 ],
   alphaCSR[ 141 ][ 116 ],
   alphaCSR[ 141 ][ 117 ],
   alphaCSR[ 141 ][ 118 ],
   alphaCSR[ 141 ][ 119 ],
   alphaCSR[ 141 ][ 120 ],
   alphaCSR[ 141 ][ 121 ],
   alphaCSR[ 141 ][ 122 ],
   alphaCSR[ 141 ][ 123 ],
   alphaCSR[ 141 ][ 124 ],
   alphaCSR[ 141 ][ 125 ],
   alphaCSR[ 141 ][ 126 ],
   alphaCSR[ 141 ][ 127 ],
   alphaCSR[ 141 ][ 128 ],
   alphaCSR[ 141 ][ 129 ],
   alphaCSR[ 141 ][ 130 ],
   alphaCSR[ 141 ][ 131 ],
   alphaCSR[ 141 ][ 132 ],
   alphaCSR[ 141 ][ 133 ],
   alphaCSR[ 141 ][ 134 ],
   alphaCSR[ 141 ][ 135 ],
   alphaCSR[ 141 ][ 136 ],
   alphaCSR[ 141 ][ 137 ],
   alphaCSR[ 141 ][ 138 ],
   alphaCSR[ 141 ][ 139 ],
   alphaCSR[ 141 ][ 140 ],
   alphaCSR[ 141 ][ 141 ],
   alphaCSR[ 141 ][ 142 ],
   alphaCSR[ 141 ][ 143 ],
   alphaCSR[ 141 ][ 144 ],
   alphaCSR[ 141 ][ 145 ],
   alphaCSR[ 141 ][ 146 ],
   alphaCSR[ 141 ][ 147 ],
   alphaCSR[ 141 ][ 148 ],
   alphaCSR[ 141 ][ 149 ],
   alphaCSR[ 141 ][ 150 ],
   alphaCSR[ 141 ][ 151 ],
   alphaCSR[ 141 ][ 152 ],
   alphaCSR[ 141 ][ 153 ],
   alphaCSR[ 141 ][ 154 ],
   alphaCSR[ 141 ][ 155 ],
   alphaCSR[ 141 ][ 156 ],
   alphaCSR[ 141 ][ 157 ],
   alphaCSR[ 141 ][ 158 ],
   alphaCSR[ 141 ][ 159 ],
   alphaCSR[ 141 ][ 160 ],
   alphaCSR[ 141 ][ 161 ],
   alphaCSR[ 141 ][ 162 ],
   alphaCSR[ 141 ][ 163 ],
   alphaCSR[ 141 ][ 164 ],
   alphaCSR[ 141 ][ 165 ],
   alphaCSR[ 141 ][ 166 ],
   alphaCSR[ 141 ][ 167 ],
   alphaCSR[ 141 ][ 168 ],
   alphaCSR[ 141 ][ 169 ],
   alphaCSR[ 141 ][ 170 ],
   alphaCSR[ 141 ][ 171 ],
   alphaCSR[ 141 ][ 172 ],
   alphaCSR[ 141 ][ 173 ],
   alphaCSR[ 141 ][ 174 ],
   alphaCSR[ 141 ][ 175 ],
   alphaCSR[ 141 ][ 176 ],
   alphaCSR[ 141 ][ 177 ],
   alphaCSR[ 141 ][ 178 ],
   alphaCSR[ 141 ][ 179 ],
   alphaCSR[ 141 ][ 180 ],
   alphaCSR[ 141 ][ 181 ],
   alphaCSR[ 141 ][ 182 ],
   alphaCSR[ 141 ][ 183 ],
   alphaCSR[ 141 ][ 184 ],
   alphaCSR[ 141 ][ 185 ],
   alphaCSR[ 141 ][ 186 ],
   alphaCSR[ 141 ][ 187 ],
   alphaCSR[ 141 ][ 188 ],
   alphaCSR[ 141 ][ 189 ],
   alphaCSR[ 141 ][ 190 ],
   alphaCSR[ 141 ][ 191 ],
   alphaCSR[ 141 ][ 192 ],
   alphaCSR[ 141 ][ 193 ],
   alphaCSR[ 141 ][ 194 ],
   alphaCSR[ 141 ][ 195 ],
   alphaCSR[ 141 ][ 196 ],
   alphaCSR[ 141 ][ 197 ],
   alphaCSR[ 141 ][ 198 ],
   alphaCSR[ 141 ][ 199 ],
   alphaCSR[ 141 ][ 200 ],
   alphaCSR[ 141 ][ 201 ],
   alphaCSR[ 141 ][ 202 ],
   alphaCSR[ 141 ][ 203 ],
   alphaCSR[ 141 ][ 204 ],
   alphaCSR[ 141 ][ 205 ],
   alphaCSR[ 141 ][ 206 ],
   alphaCSR[ 141 ][ 207 ],
   alphaCSR[ 141 ][ 208 ],
   alphaCSR[ 141 ][ 209 ],
   alphaCSR[ 141 ][ 210 ],
   alphaCSR[ 141 ][ 211 ],
   alphaCSR[ 141 ][ 212 ],
   alphaCSR[ 141 ][ 213 ],
   alphaCSR[ 141 ][ 214 ],
   alphaCSR[ 141 ][ 215 ],
   alphaCSR[ 141 ][ 216 ],
   alphaCSR[ 141 ][ 217 ],
   alphaCSR[ 141 ][ 218 ],
   alphaCSR[ 141 ][ 219 ],
   alphaCSR[ 141 ][ 220 ],
   alphaCSR[ 141 ][ 221 ],
   alphaCSR[ 141 ][ 222 ],
   alphaCSR[ 141 ][ 223 ],
   alphaCSR[ 141 ][ 224 ],
   alphaCSR[ 141 ][ 225 ],
   alphaCSR[ 141 ][ 226 ],
   alphaCSR[ 141 ][ 227 ],
   alphaCSR[ 141 ][ 228 ],
   alphaCSR[ 141 ][ 229 ],
   alphaCSR[ 141 ][ 230 ],
   alphaCSR[ 141 ][ 231 ],
   alphaCSR[ 141 ][ 232 ],
   alphaCSR[ 141 ][ 233 ],
   alphaCSR[ 141 ][ 234 ],
   alphaCSR[ 141 ][ 235 ],
   alphaCSR[ 141 ][ 236 ],
   alphaCSR[ 141 ][ 237 ],
   alphaCSR[ 141 ][ 238 ],
   alphaCSR[ 141 ][ 239 ],
   alphaCSR[ 141 ][ 240 ],
   alphaCSR[ 141 ][ 241 ],
   alphaCSR[ 141 ][ 242 ],
   alphaCSR[ 141 ][ 243 ],
   alphaCSR[ 141 ][ 244 ],
   alphaCSR[ 141 ][ 245 ],
   alphaCSR[ 141 ][ 246 ],
   alphaCSR[ 141 ][ 247 ],
   alphaCSR[ 141 ][ 248 ],
   alphaCSR[ 141 ][ 249 ],
   alphaCSR[ 141 ][ 250 ],
   alphaCSR[ 141 ][ 251 ],
   alphaCSR[ 141 ][ 252 ],
   alphaCSR[ 141 ][ 253 ],
   alphaCSR[ 141 ][ 254 ],
   alphaCSR[ 141 ][ 255 ],
   alphaCSR[ 141 ][ 256 ],
   alphaCSR[ 141 ][ 257 ],
   alphaCSR[ 141 ][ 258 ],
   alphaCSR[ 141 ][ 259 ],
   alphaCSR[ 141 ][ 260 ],
   alphaCSR[ 141 ][ 261 ],
   alphaCSR[ 141 ][ 262 ],
   alphaCSR[ 141 ][ 263 ],
   alphaCSR[ 141 ][ 264 ],
   alphaCSR[ 141 ][ 265 ],
   alphaCSR[ 141 ][ 266 ],
   alphaCSR[ 141 ][ 267 ],
   alphaCSR[ 141 ][ 268 ],
   alphaCSR[ 141 ][ 269 ],
   alphaCSR[ 141 ][ 270 ],
   alphaCSR[ 141 ][ 271 ],
   alphaCSR[ 141 ][ 272 ],
   alphaCSR[ 141 ][ 273 ],
   alphaCSR[ 141 ][ 274 ],
   alphaCSR[ 141 ][ 275 ],
   alphaCSR[ 141 ][ 276 ],
   alphaCSR[ 141 ][ 277 ],
   alphaCSR[ 141 ][ 278 ],
   alphaCSR[ 141 ][ 279 ],
   alphaCSR[ 141 ][ 280 ],
   alphaCSR[ 141 ][ 281 ],
   alphaCSR[ 141 ][ 282 ],
   alphaCSR[ 141 ][ 283 ],
   alphaCSR[ 141 ][ 284 ],
   alphaCSR[ 141 ][ 285 ],
   alphaCSR[ 141 ][ 286 ],
   alphaCSR[ 141 ][ 287 ],
   alphaCSR[ 141 ][ 288 ],
   alphaCSR[ 141 ][ 289 ],
   alphaCSR[ 141 ][ 290 ],
   alphaCSR[ 141 ][ 291 ],
   alphaCSR[ 141 ][ 292 ],
   alphaCSR[ 141 ][ 293 ],
   alphaCSR[ 141 ][ 294 ],
   alphaCSR[ 141 ][ 295 ],
   alphaCSR[ 141 ][ 296 ],
   alphaCSR[ 141 ][ 297 ],
   alphaCSR[ 141 ][ 298 ],
   alphaCSR[ 141 ][ 299 ],
   alphaCSR[ 141 ][ 300 ],
   alphaCSR[ 141 ][ 301 ],
   alphaCSR[ 141 ][ 302 ],
   alphaCSR[ 141 ][ 303 ],
   alphaCSR[ 141 ][ 304 ],
   alphaCSR[ 141 ][ 305 ],
   alphaCSR[ 141 ][ 306 ],
   alphaCSR[ 141 ][ 307 ],
   alphaCSR[ 141 ][ 308 ],
   alphaCSR[ 141 ][ 309 ],
   alphaCSR[ 141 ][ 310 ],
   alphaCSR[ 141 ][ 311 ],
   alphaCSR[ 141 ][ 312 ],
   alphaCSR[ 141 ][ 313 ],
   alphaCSR[ 141 ][ 314 ],
   alphaCSR[ 141 ][ 315 ],
   alphaCSR[ 141 ][ 316 ],
   alphaCSR[ 141 ][ 317 ],
   alphaCSR[ 141 ][ 318 ],
   alphaCSR[ 141 ][ 319 ],
   alphaCSR[ 141 ][ 320 ],
   alphaCSR[ 141 ][ 321 ],
   alphaCSR[ 141 ][ 322 ],
   alphaCSR[ 141 ][ 323 ],
   alphaCSR[ 141 ][ 324 ],
   alphaCSR[ 141 ][ 325 ],
   alphaCSR[ 141 ][ 326 ],
   alphaCSR[ 141 ][ 327 ],
   alphaCSR[ 141 ][ 328 ],
   alphaCSR[ 141 ][ 329 ],
   alphaCSR[ 141 ][ 330 ],
   alphaCSR[ 141 ][ 331 ],
   alphaCSR[ 141 ][ 332 ],
   alphaCSR[ 141 ][ 333 ],
   alphaCSR[ 141 ][ 334 ],
   alphaCSR[ 141 ][ 335 ],
   alphaCSR[ 141 ][ 336 ],
   alphaCSR[ 141 ][ 337 ],
   alphaCSR[ 141 ][ 338 ],
   alphaCSR[ 141 ][ 339 ],
   alphaCSR[ 141 ][ 340 ],
   alphaCSR[ 141 ][ 341 ],
   alphaCSR[ 141 ][ 342 ],
   alphaCSR[ 141 ][ 343 ],
   alphaCSR[ 141 ][ 344 ],
   alphaCSR[ 141 ][ 345 ],
   alphaCSR[ 141 ][ 346 ],
   alphaCSR[ 141 ][ 347 ],
   alphaCSR[ 141 ][ 348 ],
   alphaCSR[ 141 ][ 349 ],
   alphaCSR[ 141 ][ 350 ],
   alphaCSR[ 141 ][ 351 ],
   alphaCSR[ 141 ][ 352 ],
   alphaCSR[ 141 ][ 353 ],
   alphaCSR[ 141 ][ 354 ],
   alphaCSR[ 141 ][ 355 ],
   alphaCSR[ 141 ][ 356 ],
   alphaCSR[ 141 ][ 357 ],
   alphaCSR[ 141 ][ 358 ],
   alphaCSR[ 141 ][ 359 ],
   alphaCSR[ 141 ][ 360 ],
   alphaCSR[ 141 ][ 361 ],
   alphaCSR[ 141 ][ 362 ],
   alphaCSR[ 141 ][ 363 ],
   alphaCSR[ 141 ][ 364 ],
   alphaCSR[ 141 ][ 365 ],
   alphaCSR[ 141 ][ 366 ],
   alphaCSR[ 141 ][ 367 ],
   alphaCSR[ 141 ][ 368 ],
   alphaCSR[ 141 ][ 369 ],
   alphaCSR[ 141 ][ 370 ],
   alphaCSR[ 141 ][ 371 ],
   alphaCSR[ 141 ][ 372 ],
   alphaCSR[ 141 ][ 373 ],
   alphaCSR[ 141 ][ 374 ],
   alphaCSR[ 141 ][ 375 ],
   alphaCSR[ 141 ][ 376 ],
   alphaCSR[ 141 ][ 377 ],
   alphaCSR[ 141 ][ 378 ],
   alphaCSR[ 141 ][ 379 ],
   alphaCSR[ 141 ][ 380 ],
   alphaCSR[ 141 ][ 381 ],
   alphaCSR[ 141 ][ 382 ],
   alphaCSR[ 141 ][ 383 ],
   alphaCSR[ 142 ][ 0 ],
   alphaCSR[ 142 ][ 1 ],
   alphaCSR[ 142 ][ 2 ],
   alphaCSR[ 142 ][ 3 ],
   alphaCSR[ 142 ][ 4 ],
   alphaCSR[ 142 ][ 5 ],
   alphaCSR[ 142 ][ 6 ],
   alphaCSR[ 142 ][ 7 ],
   alphaCSR[ 142 ][ 8 ],
   alphaCSR[ 142 ][ 9 ],
   alphaCSR[ 142 ][ 10 ],
   alphaCSR[ 142 ][ 11 ],
   alphaCSR[ 142 ][ 12 ],
   alphaCSR[ 142 ][ 13 ],
   alphaCSR[ 142 ][ 14 ],
   alphaCSR[ 142 ][ 15 ],
   alphaCSR[ 142 ][ 16 ],
   alphaCSR[ 142 ][ 17 ],
   alphaCSR[ 142 ][ 18 ],
   alphaCSR[ 142 ][ 19 ],
   alphaCSR[ 142 ][ 20 ],
   alphaCSR[ 142 ][ 21 ],
   alphaCSR[ 142 ][ 22 ],
   alphaCSR[ 142 ][ 23 ],
   alphaCSR[ 142 ][ 24 ],
   alphaCSR[ 142 ][ 25 ],
   alphaCSR[ 142 ][ 26 ],
   alphaCSR[ 142 ][ 27 ],
   alphaCSR[ 142 ][ 28 ],
   alphaCSR[ 142 ][ 29 ],
   alphaCSR[ 142 ][ 30 ],
   alphaCSR[ 142 ][ 31 ],
   alphaCSR[ 142 ][ 32 ],
   alphaCSR[ 142 ][ 33 ],
   alphaCSR[ 142 ][ 34 ],
   alphaCSR[ 142 ][ 35 ],
   alphaCSR[ 142 ][ 36 ],
   alphaCSR[ 142 ][ 37 ],
   alphaCSR[ 142 ][ 38 ],
   alphaCSR[ 142 ][ 39 ],
   alphaCSR[ 142 ][ 40 ],
   alphaCSR[ 142 ][ 41 ],
   alphaCSR[ 142 ][ 42 ],
   alphaCSR[ 142 ][ 43 ],
   alphaCSR[ 142 ][ 44 ],
   alphaCSR[ 142 ][ 45 ],
   alphaCSR[ 142 ][ 46 ],
   alphaCSR[ 142 ][ 47 ],
   alphaCSR[ 142 ][ 48 ],
   alphaCSR[ 142 ][ 49 ],
   alphaCSR[ 142 ][ 50 ],
   alphaCSR[ 142 ][ 51 ],
   alphaCSR[ 142 ][ 52 ],
   alphaCSR[ 142 ][ 53 ],
   alphaCSR[ 142 ][ 54 ],
   alphaCSR[ 142 ][ 55 ],
   alphaCSR[ 142 ][ 56 ],
   alphaCSR[ 142 ][ 57 ],
   alphaCSR[ 142 ][ 58 ],
   alphaCSR[ 142 ][ 59 ],
   alphaCSR[ 142 ][ 60 ],
   alphaCSR[ 142 ][ 61 ],
   alphaCSR[ 142 ][ 62 ],
   alphaCSR[ 142 ][ 63 ],
   alphaCSR[ 142 ][ 64 ],
   alphaCSR[ 142 ][ 65 ],
   alphaCSR[ 142 ][ 66 ],
   alphaCSR[ 142 ][ 67 ],
   alphaCSR[ 142 ][ 68 ],
   alphaCSR[ 142 ][ 69 ],
   alphaCSR[ 142 ][ 70 ],
   alphaCSR[ 142 ][ 71 ],
   alphaCSR[ 142 ][ 72 ],
   alphaCSR[ 142 ][ 73 ],
   alphaCSR[ 142 ][ 74 ],
   alphaCSR[ 142 ][ 75 ],
   alphaCSR[ 142 ][ 76 ],
   alphaCSR[ 142 ][ 77 ],
   alphaCSR[ 142 ][ 78 ],
   alphaCSR[ 142 ][ 79 ],
   alphaCSR[ 142 ][ 80 ],
   alphaCSR[ 142 ][ 81 ],
   alphaCSR[ 142 ][ 82 ],
   alphaCSR[ 142 ][ 83 ],
   alphaCSR[ 142 ][ 84 ],
   alphaCSR[ 142 ][ 85 ],
   alphaCSR[ 142 ][ 86 ],
   alphaCSR[ 142 ][ 87 ],
   alphaCSR[ 142 ][ 88 ],
   alphaCSR[ 142 ][ 89 ],
   alphaCSR[ 142 ][ 90 ],
   alphaCSR[ 142 ][ 91 ],
   alphaCSR[ 142 ][ 92 ],
   alphaCSR[ 142 ][ 93 ],
   alphaCSR[ 142 ][ 94 ],
   alphaCSR[ 142 ][ 95 ],
   alphaCSR[ 142 ][ 96 ],
   alphaCSR[ 142 ][ 97 ],
   alphaCSR[ 142 ][ 98 ],
   alphaCSR[ 142 ][ 99 ],
   alphaCSR[ 142 ][ 100 ],
   alphaCSR[ 142 ][ 101 ],
   alphaCSR[ 142 ][ 102 ],
   alphaCSR[ 142 ][ 103 ],
   alphaCSR[ 142 ][ 104 ],
   alphaCSR[ 142 ][ 105 ],
   alphaCSR[ 142 ][ 106 ],
   alphaCSR[ 142 ][ 107 ],
   alphaCSR[ 142 ][ 108 ],
   alphaCSR[ 142 ][ 109 ],
   alphaCSR[ 142 ][ 110 ],
   alphaCSR[ 142 ][ 111 ],
   alphaCSR[ 142 ][ 112 ],
   alphaCSR[ 142 ][ 113 ],
   alphaCSR[ 142 ][ 114 ],
   alphaCSR[ 142 ][ 115 ],
   alphaCSR[ 142 ][ 116 ],
   alphaCSR[ 142 ][ 117 ],
   alphaCSR[ 142 ][ 118 ],
   alphaCSR[ 142 ][ 119 ],
   alphaCSR[ 142 ][ 120 ],
   alphaCSR[ 142 ][ 121 ],
   alphaCSR[ 142 ][ 122 ],
   alphaCSR[ 142 ][ 123 ],
   alphaCSR[ 142 ][ 124 ],
   alphaCSR[ 142 ][ 125 ],
   alphaCSR[ 142 ][ 126 ],
   alphaCSR[ 142 ][ 127 ],
   alphaCSR[ 142 ][ 128 ],
   alphaCSR[ 142 ][ 129 ],
   alphaCSR[ 142 ][ 130 ],
   alphaCSR[ 142 ][ 131 ],
   alphaCSR[ 142 ][ 132 ],
   alphaCSR[ 142 ][ 133 ],
   alphaCSR[ 142 ][ 134 ],
   alphaCSR[ 142 ][ 135 ],
   alphaCSR[ 142 ][ 136 ],
   alphaCSR[ 142 ][ 137 ],
   alphaCSR[ 142 ][ 138 ],
   alphaCSR[ 142 ][ 139 ],
   alphaCSR[ 142 ][ 140 ],
   alphaCSR[ 142 ][ 141 ],
   alphaCSR[ 142 ][ 142 ],
   alphaCSR[ 142 ][ 143 ],
   alphaCSR[ 142 ][ 144 ],
   alphaCSR[ 142 ][ 145 ],
   alphaCSR[ 142 ][ 146 ],
   alphaCSR[ 142 ][ 147 ],
   alphaCSR[ 142 ][ 148 ],
   alphaCSR[ 142 ][ 149 ],
   alphaCSR[ 142 ][ 150 ],
   alphaCSR[ 142 ][ 151 ],
   alphaCSR[ 142 ][ 152 ],
   alphaCSR[ 142 ][ 153 ],
   alphaCSR[ 142 ][ 154 ],
   alphaCSR[ 142 ][ 155 ],
   alphaCSR[ 142 ][ 156 ],
   alphaCSR[ 142 ][ 157 ],
   alphaCSR[ 142 ][ 158 ],
   alphaCSR[ 142 ][ 159 ],
   alphaCSR[ 142 ][ 160 ],
   alphaCSR[ 142 ][ 161 ],
   alphaCSR[ 142 ][ 162 ],
   alphaCSR[ 142 ][ 163 ],
   alphaCSR[ 142 ][ 164 ],
   alphaCSR[ 142 ][ 165 ],
   alphaCSR[ 142 ][ 166 ],
   alphaCSR[ 142 ][ 167 ],
   alphaCSR[ 142 ][ 168 ],
   alphaCSR[ 142 ][ 169 ],
   alphaCSR[ 142 ][ 170 ],
   alphaCSR[ 142 ][ 171 ],
   alphaCSR[ 142 ][ 172 ],
   alphaCSR[ 142 ][ 173 ],
   alphaCSR[ 142 ][ 174 ],
   alphaCSR[ 142 ][ 175 ],
   alphaCSR[ 142 ][ 176 ],
   alphaCSR[ 142 ][ 177 ],
   alphaCSR[ 142 ][ 178 ],
   alphaCSR[ 142 ][ 179 ],
   alphaCSR[ 142 ][ 180 ],
   alphaCSR[ 142 ][ 181 ],
   alphaCSR[ 142 ][ 182 ],
   alphaCSR[ 142 ][ 183 ],
   alphaCSR[ 142 ][ 184 ],
   alphaCSR[ 142 ][ 185 ],
   alphaCSR[ 142 ][ 186 ],
   alphaCSR[ 142 ][ 187 ],
   alphaCSR[ 142 ][ 188 ],
   alphaCSR[ 142 ][ 189 ],
   alphaCSR[ 142 ][ 190 ],
   alphaCSR[ 142 ][ 191 ],
   alphaCSR[ 142 ][ 192 ],
   alphaCSR[ 142 ][ 193 ],
   alphaCSR[ 142 ][ 194 ],
   alphaCSR[ 142 ][ 195 ],
   alphaCSR[ 142 ][ 196 ],
   alphaCSR[ 142 ][ 197 ],
   alphaCSR[ 142 ][ 198 ],
   alphaCSR[ 142 ][ 199 ],
   alphaCSR[ 142 ][ 200 ],
   alphaCSR[ 142 ][ 201 ],
   alphaCSR[ 142 ][ 202 ],
   alphaCSR[ 142 ][ 203 ],
   alphaCSR[ 142 ][ 204 ],
   alphaCSR[ 142 ][ 205 ],
   alphaCSR[ 142 ][ 206 ],
   alphaCSR[ 142 ][ 207 ],
   alphaCSR[ 142 ][ 208 ],
   alphaCSR[ 142 ][ 209 ],
   alphaCSR[ 142 ][ 210 ],
   alphaCSR[ 142 ][ 211 ],
   alphaCSR[ 142 ][ 212 ],
   alphaCSR[ 142 ][ 213 ],
   alphaCSR[ 142 ][ 214 ],
   alphaCSR[ 142 ][ 215 ],
   alphaCSR[ 142 ][ 216 ],
   alphaCSR[ 142 ][ 217 ],
   alphaCSR[ 142 ][ 218 ],
   alphaCSR[ 142 ][ 219 ],
   alphaCSR[ 142 ][ 220 ],
   alphaCSR[ 142 ][ 221 ],
   alphaCSR[ 142 ][ 222 ],
   alphaCSR[ 142 ][ 223 ],
   alphaCSR[ 142 ][ 224 ],
   alphaCSR[ 142 ][ 225 ],
   alphaCSR[ 142 ][ 226 ],
   alphaCSR[ 142 ][ 227 ],
   alphaCSR[ 142 ][ 228 ],
   alphaCSR[ 142 ][ 229 ],
   alphaCSR[ 142 ][ 230 ],
   alphaCSR[ 142 ][ 231 ],
   alphaCSR[ 142 ][ 232 ],
   alphaCSR[ 142 ][ 233 ],
   alphaCSR[ 142 ][ 234 ],
   alphaCSR[ 142 ][ 235 ],
   alphaCSR[ 142 ][ 236 ],
   alphaCSR[ 142 ][ 237 ],
   alphaCSR[ 142 ][ 238 ],
   alphaCSR[ 142 ][ 239 ],
   alphaCSR[ 142 ][ 240 ],
   alphaCSR[ 142 ][ 241 ],
   alphaCSR[ 142 ][ 242 ],
   alphaCSR[ 142 ][ 243 ],
   alphaCSR[ 142 ][ 244 ],
   alphaCSR[ 142 ][ 245 ],
   alphaCSR[ 142 ][ 246 ],
   alphaCSR[ 142 ][ 247 ],
   alphaCSR[ 142 ][ 248 ],
   alphaCSR[ 142 ][ 249 ],
   alphaCSR[ 142 ][ 250 ],
   alphaCSR[ 142 ][ 251 ],
   alphaCSR[ 142 ][ 252 ],
   alphaCSR[ 142 ][ 253 ],
   alphaCSR[ 142 ][ 254 ],
   alphaCSR[ 142 ][ 255 ],
   alphaCSR[ 142 ][ 256 ],
   alphaCSR[ 142 ][ 257 ],
   alphaCSR[ 142 ][ 258 ],
   alphaCSR[ 142 ][ 259 ],
   alphaCSR[ 142 ][ 260 ],
   alphaCSR[ 142 ][ 261 ],
   alphaCSR[ 142 ][ 262 ],
   alphaCSR[ 142 ][ 263 ],
   alphaCSR[ 142 ][ 264 ],
   alphaCSR[ 142 ][ 265 ],
   alphaCSR[ 142 ][ 266 ],
   alphaCSR[ 142 ][ 267 ],
   alphaCSR[ 142 ][ 268 ],
   alphaCSR[ 142 ][ 269 ],
   alphaCSR[ 142 ][ 270 ],
   alphaCSR[ 142 ][ 271 ],
   alphaCSR[ 142 ][ 272 ],
   alphaCSR[ 142 ][ 273 ],
   alphaCSR[ 142 ][ 274 ],
   alphaCSR[ 142 ][ 275 ],
   alphaCSR[ 142 ][ 276 ],
   alphaCSR[ 142 ][ 277 ],
   alphaCSR[ 142 ][ 278 ],
   alphaCSR[ 142 ][ 279 ],
   alphaCSR[ 142 ][ 280 ],
   alphaCSR[ 142 ][ 281 ],
   alphaCSR[ 142 ][ 282 ],
   alphaCSR[ 142 ][ 283 ],
   alphaCSR[ 142 ][ 284 ],
   alphaCSR[ 142 ][ 285 ],
   alphaCSR[ 142 ][ 286 ],
   alphaCSR[ 142 ][ 287 ],
   alphaCSR[ 142 ][ 288 ],
   alphaCSR[ 142 ][ 289 ],
   alphaCSR[ 142 ][ 290 ],
   alphaCSR[ 142 ][ 291 ],
   alphaCSR[ 142 ][ 292 ],
   alphaCSR[ 142 ][ 293 ],
   alphaCSR[ 142 ][ 294 ],
   alphaCSR[ 142 ][ 295 ],
   alphaCSR[ 142 ][ 296 ],
   alphaCSR[ 142 ][ 297 ],
   alphaCSR[ 142 ][ 298 ],
   alphaCSR[ 142 ][ 299 ],
   alphaCSR[ 142 ][ 300 ],
   alphaCSR[ 142 ][ 301 ],
   alphaCSR[ 142 ][ 302 ],
   alphaCSR[ 142 ][ 303 ],
   alphaCSR[ 142 ][ 304 ],
   alphaCSR[ 142 ][ 305 ],
   alphaCSR[ 142 ][ 306 ],
   alphaCSR[ 142 ][ 307 ],
   alphaCSR[ 142 ][ 308 ],
   alphaCSR[ 142 ][ 309 ],
   alphaCSR[ 142 ][ 310 ],
   alphaCSR[ 142 ][ 311 ],
   alphaCSR[ 142 ][ 312 ],
   alphaCSR[ 142 ][ 313 ],
   alphaCSR[ 142 ][ 314 ],
   alphaCSR[ 142 ][ 315 ],
   alphaCSR[ 142 ][ 316 ],
   alphaCSR[ 142 ][ 317 ],
   alphaCSR[ 142 ][ 318 ],
   alphaCSR[ 142 ][ 319 ],
   alphaCSR[ 142 ][ 320 ],
   alphaCSR[ 142 ][ 321 ],
   alphaCSR[ 142 ][ 322 ],
   alphaCSR[ 142 ][ 323 ],
   alphaCSR[ 142 ][ 324 ],
   alphaCSR[ 142 ][ 325 ],
   alphaCSR[ 142 ][ 326 ],
   alphaCSR[ 142 ][ 327 ],
   alphaCSR[ 142 ][ 328 ],
   alphaCSR[ 142 ][ 329 ],
   alphaCSR[ 142 ][ 330 ],
   alphaCSR[ 142 ][ 331 ],
   alphaCSR[ 142 ][ 332 ],
   alphaCSR[ 142 ][ 333 ],
   alphaCSR[ 142 ][ 334 ],
   alphaCSR[ 142 ][ 335 ],
   alphaCSR[ 142 ][ 336 ],
   alphaCSR[ 142 ][ 337 ],
   alphaCSR[ 142 ][ 338 ],
   alphaCSR[ 142 ][ 339 ],
   alphaCSR[ 142 ][ 340 ],
   alphaCSR[ 142 ][ 341 ],
   alphaCSR[ 142 ][ 342 ],
   alphaCSR[ 142 ][ 343 ],
   alphaCSR[ 142 ][ 344 ],
   alphaCSR[ 142 ][ 345 ],
   alphaCSR[ 142 ][ 346 ],
   alphaCSR[ 142 ][ 347 ],
   alphaCSR[ 142 ][ 348 ],
   alphaCSR[ 142 ][ 349 ],
   alphaCSR[ 142 ][ 350 ],
   alphaCSR[ 142 ][ 351 ],
   alphaCSR[ 142 ][ 352 ],
   alphaCSR[ 142 ][ 353 ],
   alphaCSR[ 142 ][ 354 ],
   alphaCSR[ 142 ][ 355 ],
   alphaCSR[ 142 ][ 356 ],
   alphaCSR[ 142 ][ 357 ],
   alphaCSR[ 142 ][ 358 ],
   alphaCSR[ 142 ][ 359 ],
   alphaCSR[ 142 ][ 360 ],
   alphaCSR[ 142 ][ 361 ],
   alphaCSR[ 142 ][ 362 ],
   alphaCSR[ 142 ][ 363 ],
   alphaCSR[ 142 ][ 364 ],
   alphaCSR[ 142 ][ 365 ],
   alphaCSR[ 142 ][ 366 ],
   alphaCSR[ 142 ][ 367 ],
   alphaCSR[ 142 ][ 368 ],
   alphaCSR[ 142 ][ 369 ],
   alphaCSR[ 142 ][ 370 ],
   alphaCSR[ 142 ][ 371 ],
   alphaCSR[ 142 ][ 372 ],
   alphaCSR[ 142 ][ 373 ],
   alphaCSR[ 142 ][ 374 ],
   alphaCSR[ 142 ][ 375 ],
   alphaCSR[ 142 ][ 376 ],
   alphaCSR[ 142 ][ 377 ],
   alphaCSR[ 142 ][ 378 ],
   alphaCSR[ 142 ][ 379 ],
   alphaCSR[ 142 ][ 380 ],
   alphaCSR[ 142 ][ 381 ],
   alphaCSR[ 142 ][ 382 ],
   alphaCSR[ 142 ][ 383 ],
   alphaCSR[ 143 ][ 0 ],
   alphaCSR[ 143 ][ 1 ],
   alphaCSR[ 143 ][ 2 ],
   alphaCSR[ 143 ][ 3 ],
   alphaCSR[ 143 ][ 4 ],
   alphaCSR[ 143 ][ 5 ],
   alphaCSR[ 143 ][ 6 ],
   alphaCSR[ 143 ][ 7 ],
   alphaCSR[ 143 ][ 8 ],
   alphaCSR[ 143 ][ 9 ],
   alphaCSR[ 143 ][ 10 ],
   alphaCSR[ 143 ][ 11 ],
   alphaCSR[ 143 ][ 12 ],
   alphaCSR[ 143 ][ 13 ],
   alphaCSR[ 143 ][ 14 ],
   alphaCSR[ 143 ][ 15 ],
   alphaCSR[ 143 ][ 16 ],
   alphaCSR[ 143 ][ 17 ],
   alphaCSR[ 143 ][ 18 ],
   alphaCSR[ 143 ][ 19 ],
   alphaCSR[ 143 ][ 20 ],
   alphaCSR[ 143 ][ 21 ],
   alphaCSR[ 143 ][ 22 ],
   alphaCSR[ 143 ][ 23 ],
   alphaCSR[ 143 ][ 24 ],
   alphaCSR[ 143 ][ 25 ],
   alphaCSR[ 143 ][ 26 ],
   alphaCSR[ 143 ][ 27 ],
   alphaCSR[ 143 ][ 28 ],
   alphaCSR[ 143 ][ 29 ],
   alphaCSR[ 143 ][ 30 ],
   alphaCSR[ 143 ][ 31 ],
   alphaCSR[ 143 ][ 32 ],
   alphaCSR[ 143 ][ 33 ],
   alphaCSR[ 143 ][ 34 ],
   alphaCSR[ 143 ][ 35 ],
   alphaCSR[ 143 ][ 36 ],
   alphaCSR[ 143 ][ 37 ],
   alphaCSR[ 143 ][ 38 ],
   alphaCSR[ 143 ][ 39 ],
   alphaCSR[ 143 ][ 40 ],
   alphaCSR[ 143 ][ 41 ],
   alphaCSR[ 143 ][ 42 ],
   alphaCSR[ 143 ][ 43 ],
   alphaCSR[ 143 ][ 44 ],
   alphaCSR[ 143 ][ 45 ],
   alphaCSR[ 143 ][ 46 ],
   alphaCSR[ 143 ][ 47 ],
   alphaCSR[ 143 ][ 48 ],
   alphaCSR[ 143 ][ 49 ],
   alphaCSR[ 143 ][ 50 ],
   alphaCSR[ 143 ][ 51 ],
   alphaCSR[ 143 ][ 52 ],
   alphaCSR[ 143 ][ 53 ],
   alphaCSR[ 143 ][ 54 ],
   alphaCSR[ 143 ][ 55 ],
   alphaCSR[ 143 ][ 56 ],
   alphaCSR[ 143 ][ 57 ],
   alphaCSR[ 143 ][ 58 ],
   alphaCSR[ 143 ][ 59 ],
   alphaCSR[ 143 ][ 60 ],
   alphaCSR[ 143 ][ 61 ],
   alphaCSR[ 143 ][ 62 ],
   alphaCSR[ 143 ][ 63 ],
   alphaCSR[ 143 ][ 64 ],
   alphaCSR[ 143 ][ 65 ],
   alphaCSR[ 143 ][ 66 ],
   alphaCSR[ 143 ][ 67 ],
   alphaCSR[ 143 ][ 68 ],
   alphaCSR[ 143 ][ 69 ],
   alphaCSR[ 143 ][ 70 ],
   alphaCSR[ 143 ][ 71 ],
   alphaCSR[ 143 ][ 72 ],
   alphaCSR[ 143 ][ 73 ],
   alphaCSR[ 143 ][ 74 ],
   alphaCSR[ 143 ][ 75 ],
   alphaCSR[ 143 ][ 76 ],
   alphaCSR[ 143 ][ 77 ],
   alphaCSR[ 143 ][ 78 ],
   alphaCSR[ 143 ][ 79 ],
   alphaCSR[ 143 ][ 80 ],
   alphaCSR[ 143 ][ 81 ],
   alphaCSR[ 143 ][ 82 ],
   alphaCSR[ 143 ][ 83 ],
   alphaCSR[ 143 ][ 84 ],
   alphaCSR[ 143 ][ 85 ],
   alphaCSR[ 143 ][ 86 ],
   alphaCSR[ 143 ][ 87 ],
   alphaCSR[ 143 ][ 88 ],
   alphaCSR[ 143 ][ 89 ],
   alphaCSR[ 143 ][ 90 ],
   alphaCSR[ 143 ][ 91 ],
   alphaCSR[ 143 ][ 92 ],
   alphaCSR[ 143 ][ 93 ],
   alphaCSR[ 143 ][ 94 ],
   alphaCSR[ 143 ][ 95 ],
   alphaCSR[ 143 ][ 96 ],
   alphaCSR[ 143 ][ 97 ],
   alphaCSR[ 143 ][ 98 ],
   alphaCSR[ 143 ][ 99 ],
   alphaCSR[ 143 ][ 100 ],
   alphaCSR[ 143 ][ 101 ],
   alphaCSR[ 143 ][ 102 ],
   alphaCSR[ 143 ][ 103 ],
   alphaCSR[ 143 ][ 104 ],
   alphaCSR[ 143 ][ 105 ],
   alphaCSR[ 143 ][ 106 ],
   alphaCSR[ 143 ][ 107 ],
   alphaCSR[ 143 ][ 108 ],
   alphaCSR[ 143 ][ 109 ],
   alphaCSR[ 143 ][ 110 ],
   alphaCSR[ 143 ][ 111 ],
   alphaCSR[ 143 ][ 112 ],
   alphaCSR[ 143 ][ 113 ],
   alphaCSR[ 143 ][ 114 ],
   alphaCSR[ 143 ][ 115 ],
   alphaCSR[ 143 ][ 116 ],
   alphaCSR[ 143 ][ 117 ],
   alphaCSR[ 143 ][ 118 ],
   alphaCSR[ 143 ][ 119 ],
   alphaCSR[ 143 ][ 120 ],
   alphaCSR[ 143 ][ 121 ],
   alphaCSR[ 143 ][ 122 ],
   alphaCSR[ 143 ][ 123 ],
   alphaCSR[ 143 ][ 124 ],
   alphaCSR[ 143 ][ 125 ],
   alphaCSR[ 143 ][ 126 ],
   alphaCSR[ 143 ][ 127 ],
   alphaCSR[ 143 ][ 128 ],
   alphaCSR[ 143 ][ 129 ],
   alphaCSR[ 143 ][ 130 ],
   alphaCSR[ 143 ][ 131 ],
   alphaCSR[ 143 ][ 132 ],
   alphaCSR[ 143 ][ 133 ],
   alphaCSR[ 143 ][ 134 ],
   alphaCSR[ 143 ][ 135 ],
   alphaCSR[ 143 ][ 136 ],
   alphaCSR[ 143 ][ 137 ],
   alphaCSR[ 143 ][ 138 ],
   alphaCSR[ 143 ][ 139 ],
   alphaCSR[ 143 ][ 140 ],
   alphaCSR[ 143 ][ 141 ],
   alphaCSR[ 143 ][ 142 ],
   alphaCSR[ 143 ][ 143 ],
   alphaCSR[ 143 ][ 144 ],
   alphaCSR[ 143 ][ 145 ],
   alphaCSR[ 143 ][ 146 ],
   alphaCSR[ 143 ][ 147 ],
   alphaCSR[ 143 ][ 148 ],
   alphaCSR[ 143 ][ 149 ],
   alphaCSR[ 143 ][ 150 ],
   alphaCSR[ 143 ][ 151 ],
   alphaCSR[ 143 ][ 152 ],
   alphaCSR[ 143 ][ 153 ],
   alphaCSR[ 143 ][ 154 ],
   alphaCSR[ 143 ][ 155 ],
   alphaCSR[ 143 ][ 156 ],
   alphaCSR[ 143 ][ 157 ],
   alphaCSR[ 143 ][ 158 ],
   alphaCSR[ 143 ][ 159 ],
   alphaCSR[ 143 ][ 160 ],
   alphaCSR[ 143 ][ 161 ],
   alphaCSR[ 143 ][ 162 ],
   alphaCSR[ 143 ][ 163 ],
   alphaCSR[ 143 ][ 164 ],
   alphaCSR[ 143 ][ 165 ],
   alphaCSR[ 143 ][ 166 ],
   alphaCSR[ 143 ][ 167 ],
   alphaCSR[ 143 ][ 168 ],
   alphaCSR[ 143 ][ 169 ],
   alphaCSR[ 143 ][ 170 ],
   alphaCSR[ 143 ][ 171 ],
   alphaCSR[ 143 ][ 172 ],
   alphaCSR[ 143 ][ 173 ],
   alphaCSR[ 143 ][ 174 ],
   alphaCSR[ 143 ][ 175 ],
   alphaCSR[ 143 ][ 176 ],
   alphaCSR[ 143 ][ 177 ],
   alphaCSR[ 143 ][ 178 ],
   alphaCSR[ 143 ][ 179 ],
   alphaCSR[ 143 ][ 180 ],
   alphaCSR[ 143 ][ 181 ],
   alphaCSR[ 143 ][ 182 ],
   alphaCSR[ 143 ][ 183 ],
   alphaCSR[ 143 ][ 184 ],
   alphaCSR[ 143 ][ 185 ],
   alphaCSR[ 143 ][ 186 ],
   alphaCSR[ 143 ][ 187 ],
   alphaCSR[ 143 ][ 188 ],
   alphaCSR[ 143 ][ 189 ],
   alphaCSR[ 143 ][ 190 ],
   alphaCSR[ 143 ][ 191 ],
   alphaCSR[ 143 ][ 192 ],
   alphaCSR[ 143 ][ 193 ],
   alphaCSR[ 143 ][ 194 ],
   alphaCSR[ 143 ][ 195 ],
   alphaCSR[ 143 ][ 196 ],
   alphaCSR[ 143 ][ 197 ],
   alphaCSR[ 143 ][ 198 ],
   alphaCSR[ 143 ][ 199 ],
   alphaCSR[ 143 ][ 200 ],
   alphaCSR[ 143 ][ 201 ],
   alphaCSR[ 143 ][ 202 ],
   alphaCSR[ 143 ][ 203 ],
   alphaCSR[ 143 ][ 204 ],
   alphaCSR[ 143 ][ 205 ],
   alphaCSR[ 143 ][ 206 ],
   alphaCSR[ 143 ][ 207 ],
   alphaCSR[ 143 ][ 208 ],
   alphaCSR[ 143 ][ 209 ],
   alphaCSR[ 143 ][ 210 ],
   alphaCSR[ 143 ][ 211 ],
   alphaCSR[ 143 ][ 212 ],
   alphaCSR[ 143 ][ 213 ],
   alphaCSR[ 143 ][ 214 ],
   alphaCSR[ 143 ][ 215 ],
   alphaCSR[ 143 ][ 216 ],
   alphaCSR[ 143 ][ 217 ],
   alphaCSR[ 143 ][ 218 ],
   alphaCSR[ 143 ][ 219 ],
   alphaCSR[ 143 ][ 220 ],
   alphaCSR[ 143 ][ 221 ],
   alphaCSR[ 143 ][ 222 ],
   alphaCSR[ 143 ][ 223 ],
   alphaCSR[ 143 ][ 224 ],
   alphaCSR[ 143 ][ 225 ],
   alphaCSR[ 143 ][ 226 ],
   alphaCSR[ 143 ][ 227 ],
   alphaCSR[ 143 ][ 228 ],
   alphaCSR[ 143 ][ 229 ],
   alphaCSR[ 143 ][ 230 ],
   alphaCSR[ 143 ][ 231 ],
   alphaCSR[ 143 ][ 232 ],
   alphaCSR[ 143 ][ 233 ],
   alphaCSR[ 143 ][ 234 ],
   alphaCSR[ 143 ][ 235 ],
   alphaCSR[ 143 ][ 236 ],
   alphaCSR[ 143 ][ 237 ],
   alphaCSR[ 143 ][ 238 ],
   alphaCSR[ 143 ][ 239 ],
   alphaCSR[ 143 ][ 240 ],
   alphaCSR[ 143 ][ 241 ],
   alphaCSR[ 143 ][ 242 ],
   alphaCSR[ 143 ][ 243 ],
   alphaCSR[ 143 ][ 244 ],
   alphaCSR[ 143 ][ 245 ],
   alphaCSR[ 143 ][ 246 ],
   alphaCSR[ 143 ][ 247 ],
   alphaCSR[ 143 ][ 248 ],
   alphaCSR[ 143 ][ 249 ],
   alphaCSR[ 143 ][ 250 ],
   alphaCSR[ 143 ][ 251 ],
   alphaCSR[ 143 ][ 252 ],
   alphaCSR[ 143 ][ 253 ],
   alphaCSR[ 143 ][ 254 ],
   alphaCSR[ 143 ][ 255 ],
   alphaCSR[ 143 ][ 256 ],
   alphaCSR[ 143 ][ 257 ],
   alphaCSR[ 143 ][ 258 ],
   alphaCSR[ 143 ][ 259 ],
   alphaCSR[ 143 ][ 260 ],
   alphaCSR[ 143 ][ 261 ],
   alphaCSR[ 143 ][ 262 ],
   alphaCSR[ 143 ][ 263 ],
   alphaCSR[ 143 ][ 264 ],
   alphaCSR[ 143 ][ 265 ],
   alphaCSR[ 143 ][ 266 ],
   alphaCSR[ 143 ][ 267 ],
   alphaCSR[ 143 ][ 268 ],
   alphaCSR[ 143 ][ 269 ],
   alphaCSR[ 143 ][ 270 ],
   alphaCSR[ 143 ][ 271 ],
   alphaCSR[ 143 ][ 272 ],
   alphaCSR[ 143 ][ 273 ],
   alphaCSR[ 143 ][ 274 ],
   alphaCSR[ 143 ][ 275 ],
   alphaCSR[ 143 ][ 276 ],
   alphaCSR[ 143 ][ 277 ],
   alphaCSR[ 143 ][ 278 ],
   alphaCSR[ 143 ][ 279 ],
   alphaCSR[ 143 ][ 280 ],
   alphaCSR[ 143 ][ 281 ],
   alphaCSR[ 143 ][ 282 ],
   alphaCSR[ 143 ][ 283 ],
   alphaCSR[ 143 ][ 284 ],
   alphaCSR[ 143 ][ 285 ],
   alphaCSR[ 143 ][ 286 ],
   alphaCSR[ 143 ][ 287 ],
   alphaCSR[ 143 ][ 288 ],
   alphaCSR[ 143 ][ 289 ],
   alphaCSR[ 143 ][ 290 ],
   alphaCSR[ 143 ][ 291 ],
   alphaCSR[ 143 ][ 292 ],
   alphaCSR[ 143 ][ 293 ],
   alphaCSR[ 143 ][ 294 ],
   alphaCSR[ 143 ][ 295 ],
   alphaCSR[ 143 ][ 296 ],
   alphaCSR[ 143 ][ 297 ],
   alphaCSR[ 143 ][ 298 ],
   alphaCSR[ 143 ][ 299 ],
   alphaCSR[ 143 ][ 300 ],
   alphaCSR[ 143 ][ 301 ],
   alphaCSR[ 143 ][ 302 ],
   alphaCSR[ 143 ][ 303 ],
   alphaCSR[ 143 ][ 304 ],
   alphaCSR[ 143 ][ 305 ],
   alphaCSR[ 143 ][ 306 ],
   alphaCSR[ 143 ][ 307 ],
   alphaCSR[ 143 ][ 308 ],
   alphaCSR[ 143 ][ 309 ],
   alphaCSR[ 143 ][ 310 ],
   alphaCSR[ 143 ][ 311 ],
   alphaCSR[ 143 ][ 312 ],
   alphaCSR[ 143 ][ 313 ],
   alphaCSR[ 143 ][ 314 ],
   alphaCSR[ 143 ][ 315 ],
   alphaCSR[ 143 ][ 316 ],
   alphaCSR[ 143 ][ 317 ],
   alphaCSR[ 143 ][ 318 ],
   alphaCSR[ 143 ][ 319 ],
   alphaCSR[ 143 ][ 320 ],
   alphaCSR[ 143 ][ 321 ],
   alphaCSR[ 143 ][ 322 ],
   alphaCSR[ 143 ][ 323 ],
   alphaCSR[ 143 ][ 324 ],
   alphaCSR[ 143 ][ 325 ],
   alphaCSR[ 143 ][ 326 ],
   alphaCSR[ 143 ][ 327 ],
   alphaCSR[ 143 ][ 328 ],
   alphaCSR[ 143 ][ 329 ],
   alphaCSR[ 143 ][ 330 ],
   alphaCSR[ 143 ][ 331 ],
   alphaCSR[ 143 ][ 332 ],
   alphaCSR[ 143 ][ 333 ],
   alphaCSR[ 143 ][ 334 ],
   alphaCSR[ 143 ][ 335 ],
   alphaCSR[ 143 ][ 336 ],
   alphaCSR[ 143 ][ 337 ],
   alphaCSR[ 143 ][ 338 ],
   alphaCSR[ 143 ][ 339 ],
   alphaCSR[ 143 ][ 340 ],
   alphaCSR[ 143 ][ 341 ],
   alphaCSR[ 143 ][ 342 ],
   alphaCSR[ 143 ][ 343 ],
   alphaCSR[ 143 ][ 344 ],
   alphaCSR[ 143 ][ 345 ],
   alphaCSR[ 143 ][ 346 ],
   alphaCSR[ 143 ][ 347 ],
   alphaCSR[ 143 ][ 348 ],
   alphaCSR[ 143 ][ 349 ],
   alphaCSR[ 143 ][ 350 ],
   alphaCSR[ 143 ][ 351 ],
   alphaCSR[ 143 ][ 352 ],
   alphaCSR[ 143 ][ 353 ],
   alphaCSR[ 143 ][ 354 ],
   alphaCSR[ 143 ][ 355 ],
   alphaCSR[ 143 ][ 356 ],
   alphaCSR[ 143 ][ 357 ],
   alphaCSR[ 143 ][ 358 ],
   alphaCSR[ 143 ][ 359 ],
   alphaCSR[ 143 ][ 360 ],
   alphaCSR[ 143 ][ 361 ],
   alphaCSR[ 143 ][ 362 ],
   alphaCSR[ 143 ][ 363 ],
   alphaCSR[ 143 ][ 364 ],
   alphaCSR[ 143 ][ 365 ],
   alphaCSR[ 143 ][ 366 ],
   alphaCSR[ 143 ][ 367 ],
   alphaCSR[ 143 ][ 368 ],
   alphaCSR[ 143 ][ 369 ],
   alphaCSR[ 143 ][ 370 ],
   alphaCSR[ 143 ][ 371 ],
   alphaCSR[ 143 ][ 372 ],
   alphaCSR[ 143 ][ 373 ],
   alphaCSR[ 143 ][ 374 ],
   alphaCSR[ 143 ][ 375 ],
   alphaCSR[ 143 ][ 376 ],
   alphaCSR[ 143 ][ 377 ],
   alphaCSR[ 143 ][ 378 ],
   alphaCSR[ 143 ][ 379 ],
   alphaCSR[ 143 ][ 380 ],
   alphaCSR[ 143 ][ 381 ],
   alphaCSR[ 143 ][ 382 ],
   alphaCSR[ 143 ][ 383 ],
   alphaCSR[ 144 ][ 0 ],
   alphaCSR[ 144 ][ 1 ],
   alphaCSR[ 144 ][ 2 ],
   alphaCSR[ 144 ][ 3 ],
   alphaCSR[ 144 ][ 4 ],
   alphaCSR[ 144 ][ 5 ],
   alphaCSR[ 144 ][ 6 ],
   alphaCSR[ 144 ][ 7 ],
   alphaCSR[ 144 ][ 8 ],
   alphaCSR[ 144 ][ 9 ],
   alphaCSR[ 144 ][ 10 ],
   alphaCSR[ 144 ][ 11 ],
   alphaCSR[ 144 ][ 12 ],
   alphaCSR[ 144 ][ 13 ],
   alphaCSR[ 144 ][ 14 ],
   alphaCSR[ 144 ][ 15 ],
   alphaCSR[ 144 ][ 16 ],
   alphaCSR[ 144 ][ 17 ],
   alphaCSR[ 144 ][ 18 ],
   alphaCSR[ 144 ][ 19 ],
   alphaCSR[ 144 ][ 20 ],
   alphaCSR[ 144 ][ 21 ],
   alphaCSR[ 144 ][ 22 ],
   alphaCSR[ 144 ][ 23 ],
   alphaCSR[ 144 ][ 24 ],
   alphaCSR[ 144 ][ 25 ],
   alphaCSR[ 144 ][ 26 ],
   alphaCSR[ 144 ][ 27 ],
   alphaCSR[ 144 ][ 28 ],
   alphaCSR[ 144 ][ 29 ],
   alphaCSR[ 144 ][ 30 ],
   alphaCSR[ 144 ][ 31 ],
   alphaCSR[ 144 ][ 32 ],
   alphaCSR[ 144 ][ 33 ],
   alphaCSR[ 144 ][ 34 ],
   alphaCSR[ 144 ][ 35 ],
   alphaCSR[ 144 ][ 36 ],
   alphaCSR[ 144 ][ 37 ],
   alphaCSR[ 144 ][ 38 ],
   alphaCSR[ 144 ][ 39 ],
   alphaCSR[ 144 ][ 40 ],
   alphaCSR[ 144 ][ 41 ],
   alphaCSR[ 144 ][ 42 ],
   alphaCSR[ 144 ][ 43 ],
   alphaCSR[ 144 ][ 44 ],
   alphaCSR[ 144 ][ 45 ],
   alphaCSR[ 144 ][ 46 ],
   alphaCSR[ 144 ][ 47 ],
   alphaCSR[ 144 ][ 48 ],
   alphaCSR[ 144 ][ 49 ],
   alphaCSR[ 144 ][ 50 ],
   alphaCSR[ 144 ][ 51 ],
   alphaCSR[ 144 ][ 52 ],
   alphaCSR[ 144 ][ 53 ],
   alphaCSR[ 144 ][ 54 ],
   alphaCSR[ 144 ][ 55 ],
   alphaCSR[ 144 ][ 56 ],
   alphaCSR[ 144 ][ 57 ],
   alphaCSR[ 144 ][ 58 ],
   alphaCSR[ 144 ][ 59 ],
   alphaCSR[ 144 ][ 60 ],
   alphaCSR[ 144 ][ 61 ],
   alphaCSR[ 144 ][ 62 ],
   alphaCSR[ 144 ][ 63 ],
   alphaCSR[ 144 ][ 64 ],
   alphaCSR[ 144 ][ 65 ],
   alphaCSR[ 144 ][ 66 ],
   alphaCSR[ 144 ][ 67 ],
   alphaCSR[ 144 ][ 68 ],
   alphaCSR[ 144 ][ 69 ],
   alphaCSR[ 144 ][ 70 ],
   alphaCSR[ 144 ][ 71 ],
   alphaCSR[ 144 ][ 72 ],
   alphaCSR[ 144 ][ 73 ],
   alphaCSR[ 144 ][ 74 ],
   alphaCSR[ 144 ][ 75 ],
   alphaCSR[ 144 ][ 76 ],
   alphaCSR[ 144 ][ 77 ],
   alphaCSR[ 144 ][ 78 ],
   alphaCSR[ 144 ][ 79 ],
   alphaCSR[ 144 ][ 80 ],
   alphaCSR[ 144 ][ 81 ],
   alphaCSR[ 144 ][ 82 ],
   alphaCSR[ 144 ][ 83 ],
   alphaCSR[ 144 ][ 84 ],
   alphaCSR[ 144 ][ 85 ],
   alphaCSR[ 144 ][ 86 ],
   alphaCSR[ 144 ][ 87 ],
   alphaCSR[ 144 ][ 88 ],
   alphaCSR[ 144 ][ 89 ],
   alphaCSR[ 144 ][ 90 ],
   alphaCSR[ 144 ][ 91 ],
   alphaCSR[ 144 ][ 92 ],
   alphaCSR[ 144 ][ 93 ],
   alphaCSR[ 144 ][ 94 ],
   alphaCSR[ 144 ][ 95 ],
   alphaCSR[ 144 ][ 96 ],
   alphaCSR[ 144 ][ 97 ],
   alphaCSR[ 144 ][ 98 ],
   alphaCSR[ 144 ][ 99 ],
   alphaCSR[ 144 ][ 100 ],
   alphaCSR[ 144 ][ 101 ],
   alphaCSR[ 144 ][ 102 ],
   alphaCSR[ 144 ][ 103 ],
   alphaCSR[ 144 ][ 104 ],
   alphaCSR[ 144 ][ 105 ],
   alphaCSR[ 144 ][ 106 ],
   alphaCSR[ 144 ][ 107 ],
   alphaCSR[ 144 ][ 108 ],
   alphaCSR[ 144 ][ 109 ],
   alphaCSR[ 144 ][ 110 ],
   alphaCSR[ 144 ][ 111 ],
   alphaCSR[ 144 ][ 112 ],
   alphaCSR[ 144 ][ 113 ],
   alphaCSR[ 144 ][ 114 ],
   alphaCSR[ 144 ][ 115 ],
   alphaCSR[ 144 ][ 116 ],
   alphaCSR[ 144 ][ 117 ],
   alphaCSR[ 144 ][ 118 ],
   alphaCSR[ 144 ][ 119 ],
   alphaCSR[ 144 ][ 120 ],
   alphaCSR[ 144 ][ 121 ],
   alphaCSR[ 144 ][ 122 ],
   alphaCSR[ 144 ][ 123 ],
   alphaCSR[ 144 ][ 124 ],
   alphaCSR[ 144 ][ 125 ],
   alphaCSR[ 144 ][ 126 ],
   alphaCSR[ 144 ][ 127 ],
   alphaCSR[ 144 ][ 128 ],
   alphaCSR[ 144 ][ 129 ],
   alphaCSR[ 144 ][ 130 ],
   alphaCSR[ 144 ][ 131 ],
   alphaCSR[ 144 ][ 132 ],
   alphaCSR[ 144 ][ 133 ],
   alphaCSR[ 144 ][ 134 ],
   alphaCSR[ 144 ][ 135 ],
   alphaCSR[ 144 ][ 136 ],
   alphaCSR[ 144 ][ 137 ],
   alphaCSR[ 144 ][ 138 ],
   alphaCSR[ 144 ][ 139 ],
   alphaCSR[ 144 ][ 140 ],
   alphaCSR[ 144 ][ 141 ],
   alphaCSR[ 144 ][ 142 ],
   alphaCSR[ 144 ][ 143 ],
   alphaCSR[ 144 ][ 144 ],
   alphaCSR[ 144 ][ 145 ],
   alphaCSR[ 144 ][ 146 ],
   alphaCSR[ 144 ][ 147 ],
   alphaCSR[ 144 ][ 148 ],
   alphaCSR[ 144 ][ 149 ],
   alphaCSR[ 144 ][ 150 ],
   alphaCSR[ 144 ][ 151 ],
   alphaCSR[ 144 ][ 152 ],
   alphaCSR[ 144 ][ 153 ],
   alphaCSR[ 144 ][ 154 ],
   alphaCSR[ 144 ][ 155 ],
   alphaCSR[ 144 ][ 156 ],
   alphaCSR[ 144 ][ 157 ],
   alphaCSR[ 144 ][ 158 ],
   alphaCSR[ 144 ][ 159 ],
   alphaCSR[ 144 ][ 160 ],
   alphaCSR[ 144 ][ 161 ],
   alphaCSR[ 144 ][ 162 ],
   alphaCSR[ 144 ][ 163 ],
   alphaCSR[ 144 ][ 164 ],
   alphaCSR[ 144 ][ 165 ],
   alphaCSR[ 144 ][ 166 ],
   alphaCSR[ 144 ][ 167 ],
   alphaCSR[ 144 ][ 168 ],
   alphaCSR[ 144 ][ 169 ],
   alphaCSR[ 144 ][ 170 ],
   alphaCSR[ 144 ][ 171 ],
   alphaCSR[ 144 ][ 172 ],
   alphaCSR[ 144 ][ 173 ],
   alphaCSR[ 144 ][ 174 ],
   alphaCSR[ 144 ][ 175 ],
   alphaCSR[ 144 ][ 176 ],
   alphaCSR[ 144 ][ 177 ],
   alphaCSR[ 144 ][ 178 ],
   alphaCSR[ 144 ][ 179 ],
   alphaCSR[ 144 ][ 180 ],
   alphaCSR[ 144 ][ 181 ],
   alphaCSR[ 144 ][ 182 ],
   alphaCSR[ 144 ][ 183 ],
   alphaCSR[ 144 ][ 184 ],
   alphaCSR[ 144 ][ 185 ],
   alphaCSR[ 144 ][ 186 ],
   alphaCSR[ 144 ][ 187 ],
   alphaCSR[ 144 ][ 188 ],
   alphaCSR[ 144 ][ 189 ],
   alphaCSR[ 144 ][ 190 ],
   alphaCSR[ 144 ][ 191 ],
   alphaCSR[ 144 ][ 192 ],
   alphaCSR[ 144 ][ 193 ],
   alphaCSR[ 144 ][ 194 ],
   alphaCSR[ 144 ][ 195 ],
   alphaCSR[ 144 ][ 196 ],
   alphaCSR[ 144 ][ 197 ],
   alphaCSR[ 144 ][ 198 ],
   alphaCSR[ 144 ][ 199 ],
   alphaCSR[ 144 ][ 200 ],
   alphaCSR[ 144 ][ 201 ],
   alphaCSR[ 144 ][ 202 ],
   alphaCSR[ 144 ][ 203 ],
   alphaCSR[ 144 ][ 204 ],
   alphaCSR[ 144 ][ 205 ],
   alphaCSR[ 144 ][ 206 ],
   alphaCSR[ 144 ][ 207 ],
   alphaCSR[ 144 ][ 208 ],
   alphaCSR[ 144 ][ 209 ],
   alphaCSR[ 144 ][ 210 ],
   alphaCSR[ 144 ][ 211 ],
   alphaCSR[ 144 ][ 212 ],
   alphaCSR[ 144 ][ 213 ],
   alphaCSR[ 144 ][ 214 ],
   alphaCSR[ 144 ][ 215 ],
   alphaCSR[ 144 ][ 216 ],
   alphaCSR[ 144 ][ 217 ],
   alphaCSR[ 144 ][ 218 ],
   alphaCSR[ 144 ][ 219 ],
   alphaCSR[ 144 ][ 220 ],
   alphaCSR[ 144 ][ 221 ],
   alphaCSR[ 144 ][ 222 ],
   alphaCSR[ 144 ][ 223 ],
   alphaCSR[ 144 ][ 224 ],
   alphaCSR[ 144 ][ 225 ],
   alphaCSR[ 144 ][ 226 ],
   alphaCSR[ 144 ][ 227 ],
   alphaCSR[ 144 ][ 228 ],
   alphaCSR[ 144 ][ 229 ],
   alphaCSR[ 144 ][ 230 ],
   alphaCSR[ 144 ][ 231 ],
   alphaCSR[ 144 ][ 232 ],
   alphaCSR[ 144 ][ 233 ],
   alphaCSR[ 144 ][ 234 ],
   alphaCSR[ 144 ][ 235 ],
   alphaCSR[ 144 ][ 236 ],
   alphaCSR[ 144 ][ 237 ],
   alphaCSR[ 144 ][ 238 ],
   alphaCSR[ 144 ][ 239 ],
   alphaCSR[ 144 ][ 240 ],
   alphaCSR[ 144 ][ 241 ],
   alphaCSR[ 144 ][ 242 ],
   alphaCSR[ 144 ][ 243 ],
   alphaCSR[ 144 ][ 244 ],
   alphaCSR[ 144 ][ 245 ],
   alphaCSR[ 144 ][ 246 ],
   alphaCSR[ 144 ][ 247 ],
   alphaCSR[ 144 ][ 248 ],
   alphaCSR[ 144 ][ 249 ],
   alphaCSR[ 144 ][ 250 ],
   alphaCSR[ 144 ][ 251 ],
   alphaCSR[ 144 ][ 252 ],
   alphaCSR[ 144 ][ 253 ],
   alphaCSR[ 144 ][ 254 ],
   alphaCSR[ 144 ][ 255 ],
   alphaCSR[ 144 ][ 256 ],
   alphaCSR[ 144 ][ 257 ],
   alphaCSR[ 144 ][ 258 ],
   alphaCSR[ 144 ][ 259 ],
   alphaCSR[ 144 ][ 260 ],
   alphaCSR[ 144 ][ 261 ],
   alphaCSR[ 144 ][ 262 ],
   alphaCSR[ 144 ][ 263 ],
   alphaCSR[ 144 ][ 264 ],
   alphaCSR[ 144 ][ 265 ],
   alphaCSR[ 144 ][ 266 ],
   alphaCSR[ 144 ][ 267 ],
   alphaCSR[ 144 ][ 268 ],
   alphaCSR[ 144 ][ 269 ],
   alphaCSR[ 144 ][ 270 ],
   alphaCSR[ 144 ][ 271 ],
   alphaCSR[ 144 ][ 272 ],
   alphaCSR[ 144 ][ 273 ],
   alphaCSR[ 144 ][ 274 ],
   alphaCSR[ 144 ][ 275 ],
   alphaCSR[ 144 ][ 276 ],
   alphaCSR[ 144 ][ 277 ],
   alphaCSR[ 144 ][ 278 ],
   alphaCSR[ 144 ][ 279 ],
   alphaCSR[ 144 ][ 280 ],
   alphaCSR[ 144 ][ 281 ],
   alphaCSR[ 144 ][ 282 ],
   alphaCSR[ 144 ][ 283 ],
   alphaCSR[ 144 ][ 284 ],
   alphaCSR[ 144 ][ 285 ],
   alphaCSR[ 144 ][ 286 ],
   alphaCSR[ 144 ][ 287 ],
   alphaCSR[ 144 ][ 288 ],
   alphaCSR[ 144 ][ 289 ],
   alphaCSR[ 144 ][ 290 ],
   alphaCSR[ 144 ][ 291 ],
   alphaCSR[ 144 ][ 292 ],
   alphaCSR[ 144 ][ 293 ],
   alphaCSR[ 144 ][ 294 ],
   alphaCSR[ 144 ][ 295 ],
   alphaCSR[ 144 ][ 296 ],
   alphaCSR[ 144 ][ 297 ],
   alphaCSR[ 144 ][ 298 ],
   alphaCSR[ 144 ][ 299 ],
   alphaCSR[ 144 ][ 300 ],
   alphaCSR[ 144 ][ 301 ],
   alphaCSR[ 144 ][ 302 ],
   alphaCSR[ 144 ][ 303 ],
   alphaCSR[ 144 ][ 304 ],
   alphaCSR[ 144 ][ 305 ],
   alphaCSR[ 144 ][ 306 ],
   alphaCSR[ 144 ][ 307 ],
   alphaCSR[ 144 ][ 308 ],
   alphaCSR[ 144 ][ 309 ],
   alphaCSR[ 144 ][ 310 ],
   alphaCSR[ 144 ][ 311 ],
   alphaCSR[ 144 ][ 312 ],
   alphaCSR[ 144 ][ 313 ],
   alphaCSR[ 144 ][ 314 ],
   alphaCSR[ 144 ][ 315 ],
   alphaCSR[ 144 ][ 316 ],
   alphaCSR[ 144 ][ 317 ],
   alphaCSR[ 144 ][ 318 ],
   alphaCSR[ 144 ][ 319 ],
   alphaCSR[ 144 ][ 320 ],
   alphaCSR[ 144 ][ 321 ],
   alphaCSR[ 144 ][ 322 ],
   alphaCSR[ 144 ][ 323 ],
   alphaCSR[ 144 ][ 324 ],
   alphaCSR[ 144 ][ 325 ],
   alphaCSR[ 144 ][ 326 ],
   alphaCSR[ 144 ][ 327 ],
   alphaCSR[ 144 ][ 328 ],
   alphaCSR[ 144 ][ 329 ],
   alphaCSR[ 144 ][ 330 ],
   alphaCSR[ 144 ][ 331 ],
   alphaCSR[ 144 ][ 332 ],
   alphaCSR[ 144 ][ 333 ],
   alphaCSR[ 144 ][ 334 ],
   alphaCSR[ 144 ][ 335 ],
   alphaCSR[ 144 ][ 336 ],
   alphaCSR[ 144 ][ 337 ],
   alphaCSR[ 144 ][ 338 ],
   alphaCSR[ 144 ][ 339 ],
   alphaCSR[ 144 ][ 340 ],
   alphaCSR[ 144 ][ 341 ],
   alphaCSR[ 144 ][ 342 ],
   alphaCSR[ 144 ][ 343 ],
   alphaCSR[ 144 ][ 344 ],
   alphaCSR[ 144 ][ 345 ],
   alphaCSR[ 144 ][ 346 ],
   alphaCSR[ 144 ][ 347 ],
   alphaCSR[ 144 ][ 348 ],
   alphaCSR[ 144 ][ 349 ],
   alphaCSR[ 144 ][ 350 ],
   alphaCSR[ 144 ][ 351 ],
   alphaCSR[ 144 ][ 352 ],
   alphaCSR[ 144 ][ 353 ],
   alphaCSR[ 144 ][ 354 ],
   alphaCSR[ 144 ][ 355 ],
   alphaCSR[ 144 ][ 356 ],
   alphaCSR[ 144 ][ 357 ],
   alphaCSR[ 144 ][ 358 ],
   alphaCSR[ 144 ][ 359 ],
   alphaCSR[ 144 ][ 360 ],
   alphaCSR[ 144 ][ 361 ],
   alphaCSR[ 144 ][ 362 ],
   alphaCSR[ 144 ][ 363 ],
   alphaCSR[ 144 ][ 364 ],
   alphaCSR[ 144 ][ 365 ],
   alphaCSR[ 144 ][ 366 ],
   alphaCSR[ 144 ][ 367 ],
   alphaCSR[ 144 ][ 368 ],
   alphaCSR[ 144 ][ 369 ],
   alphaCSR[ 144 ][ 370 ],
   alphaCSR[ 144 ][ 371 ],
   alphaCSR[ 144 ][ 372 ],
   alphaCSR[ 144 ][ 373 ],
   alphaCSR[ 144 ][ 374 ],
   alphaCSR[ 144 ][ 375 ],
   alphaCSR[ 144 ][ 376 ],
   alphaCSR[ 144 ][ 377 ],
   alphaCSR[ 144 ][ 378 ],
   alphaCSR[ 144 ][ 379 ],
   alphaCSR[ 144 ][ 380 ],
   alphaCSR[ 144 ][ 381 ],
   alphaCSR[ 144 ][ 382 ],
   alphaCSR[ 144 ][ 383 ],
   alphaCSR[ 145 ][ 0 ],
   alphaCSR[ 145 ][ 1 ],
   alphaCSR[ 145 ][ 2 ],
   alphaCSR[ 145 ][ 3 ],
   alphaCSR[ 145 ][ 4 ],
   alphaCSR[ 145 ][ 5 ],
   alphaCSR[ 145 ][ 6 ],
   alphaCSR[ 145 ][ 7 ],
   alphaCSR[ 145 ][ 8 ],
   alphaCSR[ 145 ][ 9 ],
   alphaCSR[ 145 ][ 10 ],
   alphaCSR[ 145 ][ 11 ],
   alphaCSR[ 145 ][ 12 ],
   alphaCSR[ 145 ][ 13 ],
   alphaCSR[ 145 ][ 14 ],
   alphaCSR[ 145 ][ 15 ],
   alphaCSR[ 145 ][ 16 ],
   alphaCSR[ 145 ][ 17 ],
   alphaCSR[ 145 ][ 18 ],
   alphaCSR[ 145 ][ 19 ],
   alphaCSR[ 145 ][ 20 ],
   alphaCSR[ 145 ][ 21 ],
   alphaCSR[ 145 ][ 22 ],
   alphaCSR[ 145 ][ 23 ],
   alphaCSR[ 145 ][ 24 ],
   alphaCSR[ 145 ][ 25 ],
   alphaCSR[ 145 ][ 26 ],
   alphaCSR[ 145 ][ 27 ],
   alphaCSR[ 145 ][ 28 ],
   alphaCSR[ 145 ][ 29 ],
   alphaCSR[ 145 ][ 30 ],
   alphaCSR[ 145 ][ 31 ],
   alphaCSR[ 145 ][ 32 ],
   alphaCSR[ 145 ][ 33 ],
   alphaCSR[ 145 ][ 34 ],
   alphaCSR[ 145 ][ 35 ],
   alphaCSR[ 145 ][ 36 ],
   alphaCSR[ 145 ][ 37 ],
   alphaCSR[ 145 ][ 38 ],
   alphaCSR[ 145 ][ 39 ],
   alphaCSR[ 145 ][ 40 ],
   alphaCSR[ 145 ][ 41 ],
   alphaCSR[ 145 ][ 42 ],
   alphaCSR[ 145 ][ 43 ],
   alphaCSR[ 145 ][ 44 ],
   alphaCSR[ 145 ][ 45 ],
   alphaCSR[ 145 ][ 46 ],
   alphaCSR[ 145 ][ 47 ],
   alphaCSR[ 145 ][ 48 ],
   alphaCSR[ 145 ][ 49 ],
   alphaCSR[ 145 ][ 50 ],
   alphaCSR[ 145 ][ 51 ],
   alphaCSR[ 145 ][ 52 ],
   alphaCSR[ 145 ][ 53 ],
   alphaCSR[ 145 ][ 54 ],
   alphaCSR[ 145 ][ 55 ],
   alphaCSR[ 145 ][ 56 ],
   alphaCSR[ 145 ][ 57 ],
   alphaCSR[ 145 ][ 58 ],
   alphaCSR[ 145 ][ 59 ],
   alphaCSR[ 145 ][ 60 ],
   alphaCSR[ 145 ][ 61 ],
   alphaCSR[ 145 ][ 62 ],
   alphaCSR[ 145 ][ 63 ],
   alphaCSR[ 145 ][ 64 ],
   alphaCSR[ 145 ][ 65 ],
   alphaCSR[ 145 ][ 66 ],
   alphaCSR[ 145 ][ 67 ],
   alphaCSR[ 145 ][ 68 ],
   alphaCSR[ 145 ][ 69 ],
   alphaCSR[ 145 ][ 70 ],
   alphaCSR[ 145 ][ 71 ],
   alphaCSR[ 145 ][ 72 ],
   alphaCSR[ 145 ][ 73 ],
   alphaCSR[ 145 ][ 74 ],
   alphaCSR[ 145 ][ 75 ],
   alphaCSR[ 145 ][ 76 ],
   alphaCSR[ 145 ][ 77 ],
   alphaCSR[ 145 ][ 78 ],
   alphaCSR[ 145 ][ 79 ],
   alphaCSR[ 145 ][ 80 ],
   alphaCSR[ 145 ][ 81 ],
   alphaCSR[ 145 ][ 82 ],
   alphaCSR[ 145 ][ 83 ],
   alphaCSR[ 145 ][ 84 ],
   alphaCSR[ 145 ][ 85 ],
   alphaCSR[ 145 ][ 86 ],
   alphaCSR[ 145 ][ 87 ],
   alphaCSR[ 145 ][ 88 ],
   alphaCSR[ 145 ][ 89 ],
   alphaCSR[ 145 ][ 90 ],
   alphaCSR[ 145 ][ 91 ],
   alphaCSR[ 145 ][ 92 ],
   alphaCSR[ 145 ][ 93 ],
   alphaCSR[ 145 ][ 94 ],
   alphaCSR[ 145 ][ 95 ],
   alphaCSR[ 145 ][ 96 ],
   alphaCSR[ 145 ][ 97 ],
   alphaCSR[ 145 ][ 98 ],
   alphaCSR[ 145 ][ 99 ],
   alphaCSR[ 145 ][ 100 ],
   alphaCSR[ 145 ][ 101 ],
   alphaCSR[ 145 ][ 102 ],
   alphaCSR[ 145 ][ 103 ],
   alphaCSR[ 145 ][ 104 ],
   alphaCSR[ 145 ][ 105 ],
   alphaCSR[ 145 ][ 106 ],
   alphaCSR[ 145 ][ 107 ],
   alphaCSR[ 145 ][ 108 ],
   alphaCSR[ 145 ][ 109 ],
   alphaCSR[ 145 ][ 110 ],
   alphaCSR[ 145 ][ 111 ],
   alphaCSR[ 145 ][ 112 ],
   alphaCSR[ 145 ][ 113 ],
   alphaCSR[ 145 ][ 114 ],
   alphaCSR[ 145 ][ 115 ],
   alphaCSR[ 145 ][ 116 ],
   alphaCSR[ 145 ][ 117 ],
   alphaCSR[ 145 ][ 118 ],
   alphaCSR[ 145 ][ 119 ],
   alphaCSR[ 145 ][ 120 ],
   alphaCSR[ 145 ][ 121 ],
   alphaCSR[ 145 ][ 122 ],
   alphaCSR[ 145 ][ 123 ],
   alphaCSR[ 145 ][ 124 ],
   alphaCSR[ 145 ][ 125 ],
   alphaCSR[ 145 ][ 126 ],
   alphaCSR[ 145 ][ 127 ],
   alphaCSR[ 145 ][ 128 ],
   alphaCSR[ 145 ][ 129 ],
   alphaCSR[ 145 ][ 130 ],
   alphaCSR[ 145 ][ 131 ],
   alphaCSR[ 145 ][ 132 ],
   alphaCSR[ 145 ][ 133 ],
   alphaCSR[ 145 ][ 134 ],
   alphaCSR[ 145 ][ 135 ],
   alphaCSR[ 145 ][ 136 ],
   alphaCSR[ 145 ][ 137 ],
   alphaCSR[ 145 ][ 138 ],
   alphaCSR[ 145 ][ 139 ],
   alphaCSR[ 145 ][ 140 ],
   alphaCSR[ 145 ][ 141 ],
   alphaCSR[ 145 ][ 142 ],
   alphaCSR[ 145 ][ 143 ],
   alphaCSR[ 145 ][ 144 ],
   alphaCSR[ 145 ][ 145 ],
   alphaCSR[ 145 ][ 146 ],
   alphaCSR[ 145 ][ 147 ],
   alphaCSR[ 145 ][ 148 ],
   alphaCSR[ 145 ][ 149 ],
   alphaCSR[ 145 ][ 150 ],
   alphaCSR[ 145 ][ 151 ],
   alphaCSR[ 145 ][ 152 ],
   alphaCSR[ 145 ][ 153 ],
   alphaCSR[ 145 ][ 154 ],
   alphaCSR[ 145 ][ 155 ],
   alphaCSR[ 145 ][ 156 ],
   alphaCSR[ 145 ][ 157 ],
   alphaCSR[ 145 ][ 158 ],
   alphaCSR[ 145 ][ 159 ],
   alphaCSR[ 145 ][ 160 ],
   alphaCSR[ 145 ][ 161 ],
   alphaCSR[ 145 ][ 162 ],
   alphaCSR[ 145 ][ 163 ],
   alphaCSR[ 145 ][ 164 ],
   alphaCSR[ 145 ][ 165 ],
   alphaCSR[ 145 ][ 166 ],
   alphaCSR[ 145 ][ 167 ],
   alphaCSR[ 145 ][ 168 ],
   alphaCSR[ 145 ][ 169 ],
   alphaCSR[ 145 ][ 170 ],
   alphaCSR[ 145 ][ 171 ],
   alphaCSR[ 145 ][ 172 ],
   alphaCSR[ 145 ][ 173 ],
   alphaCSR[ 145 ][ 174 ],
   alphaCSR[ 145 ][ 175 ],
   alphaCSR[ 145 ][ 176 ],
   alphaCSR[ 145 ][ 177 ],
   alphaCSR[ 145 ][ 178 ],
   alphaCSR[ 145 ][ 179 ],
   alphaCSR[ 145 ][ 180 ],
   alphaCSR[ 145 ][ 181 ],
   alphaCSR[ 145 ][ 182 ],
   alphaCSR[ 145 ][ 183 ],
   alphaCSR[ 145 ][ 184 ],
   alphaCSR[ 145 ][ 185 ],
   alphaCSR[ 145 ][ 186 ],
   alphaCSR[ 145 ][ 187 ],
   alphaCSR[ 145 ][ 188 ],
   alphaCSR[ 145 ][ 189 ],
   alphaCSR[ 145 ][ 190 ],
   alphaCSR[ 145 ][ 191 ],
   alphaCSR[ 145 ][ 192 ],
   alphaCSR[ 145 ][ 193 ],
   alphaCSR[ 145 ][ 194 ],
   alphaCSR[ 145 ][ 195 ],
   alphaCSR[ 145 ][ 196 ],
   alphaCSR[ 145 ][ 197 ],
   alphaCSR[ 145 ][ 198 ],
   alphaCSR[ 145 ][ 199 ],
   alphaCSR[ 145 ][ 200 ],
   alphaCSR[ 145 ][ 201 ],
   alphaCSR[ 145 ][ 202 ],
   alphaCSR[ 145 ][ 203 ],
   alphaCSR[ 145 ][ 204 ],
   alphaCSR[ 145 ][ 205 ],
   alphaCSR[ 145 ][ 206 ],
   alphaCSR[ 145 ][ 207 ],
   alphaCSR[ 145 ][ 208 ],
   alphaCSR[ 145 ][ 209 ],
   alphaCSR[ 145 ][ 210 ],
   alphaCSR[ 145 ][ 211 ],
   alphaCSR[ 145 ][ 212 ],
   alphaCSR[ 145 ][ 213 ],
   alphaCSR[ 145 ][ 214 ],
   alphaCSR[ 145 ][ 215 ],
   alphaCSR[ 145 ][ 216 ],
   alphaCSR[ 145 ][ 217 ],
   alphaCSR[ 145 ][ 218 ],
   alphaCSR[ 145 ][ 219 ],
   alphaCSR[ 145 ][ 220 ],
   alphaCSR[ 145 ][ 221 ],
   alphaCSR[ 145 ][ 222 ],
   alphaCSR[ 145 ][ 223 ],
   alphaCSR[ 145 ][ 224 ],
   alphaCSR[ 145 ][ 225 ],
   alphaCSR[ 145 ][ 226 ],
   alphaCSR[ 145 ][ 227 ],
   alphaCSR[ 145 ][ 228 ],
   alphaCSR[ 145 ][ 229 ],
   alphaCSR[ 145 ][ 230 ],
   alphaCSR[ 145 ][ 231 ],
   alphaCSR[ 145 ][ 232 ],
   alphaCSR[ 145 ][ 233 ],
   alphaCSR[ 145 ][ 234 ],
   alphaCSR[ 145 ][ 235 ],
   alphaCSR[ 145 ][ 236 ],
   alphaCSR[ 145 ][ 237 ],
   alphaCSR[ 145 ][ 238 ],
   alphaCSR[ 145 ][ 239 ],
   alphaCSR[ 145 ][ 240 ],
   alphaCSR[ 145 ][ 241 ],
   alphaCSR[ 145 ][ 242 ],
   alphaCSR[ 145 ][ 243 ],
   alphaCSR[ 145 ][ 244 ],
   alphaCSR[ 145 ][ 245 ],
   alphaCSR[ 145 ][ 246 ],
   alphaCSR[ 145 ][ 247 ],
   alphaCSR[ 145 ][ 248 ],
   alphaCSR[ 145 ][ 249 ],
   alphaCSR[ 145 ][ 250 ],
   alphaCSR[ 145 ][ 251 ],
   alphaCSR[ 145 ][ 252 ],
   alphaCSR[ 145 ][ 253 ],
   alphaCSR[ 145 ][ 254 ],
   alphaCSR[ 145 ][ 255 ],
   alphaCSR[ 145 ][ 256 ],
   alphaCSR[ 145 ][ 257 ],
   alphaCSR[ 145 ][ 258 ],
   alphaCSR[ 145 ][ 259 ],
   alphaCSR[ 145 ][ 260 ],
   alphaCSR[ 145 ][ 261 ],
   alphaCSR[ 145 ][ 262 ],
   alphaCSR[ 145 ][ 263 ],
   alphaCSR[ 145 ][ 264 ],
   alphaCSR[ 145 ][ 265 ],
   alphaCSR[ 145 ][ 266 ],
   alphaCSR[ 145 ][ 267 ],
   alphaCSR[ 145 ][ 268 ],
   alphaCSR[ 145 ][ 269 ],
   alphaCSR[ 145 ][ 270 ],
   alphaCSR[ 145 ][ 271 ],
   alphaCSR[ 145 ][ 272 ],
   alphaCSR[ 145 ][ 273 ],
   alphaCSR[ 145 ][ 274 ],
   alphaCSR[ 145 ][ 275 ],
   alphaCSR[ 145 ][ 276 ],
   alphaCSR[ 145 ][ 277 ],
   alphaCSR[ 145 ][ 278 ],
   alphaCSR[ 145 ][ 279 ],
   alphaCSR[ 145 ][ 280 ],
   alphaCSR[ 145 ][ 281 ],
   alphaCSR[ 145 ][ 282 ],
   alphaCSR[ 145 ][ 283 ],
   alphaCSR[ 145 ][ 284 ],
   alphaCSR[ 145 ][ 285 ],
   alphaCSR[ 145 ][ 286 ],
   alphaCSR[ 145 ][ 287 ],
   alphaCSR[ 145 ][ 288 ],
   alphaCSR[ 145 ][ 289 ],
   alphaCSR[ 145 ][ 290 ],
   alphaCSR[ 145 ][ 291 ],
   alphaCSR[ 145 ][ 292 ],
   alphaCSR[ 145 ][ 293 ],
   alphaCSR[ 145 ][ 294 ],
   alphaCSR[ 145 ][ 295 ],
   alphaCSR[ 145 ][ 296 ],
   alphaCSR[ 145 ][ 297 ],
   alphaCSR[ 145 ][ 298 ],
   alphaCSR[ 145 ][ 299 ],
   alphaCSR[ 145 ][ 300 ],
   alphaCSR[ 145 ][ 301 ],
   alphaCSR[ 145 ][ 302 ],
   alphaCSR[ 145 ][ 303 ],
   alphaCSR[ 145 ][ 304 ],
   alphaCSR[ 145 ][ 305 ],
   alphaCSR[ 145 ][ 306 ],
   alphaCSR[ 145 ][ 307 ],
   alphaCSR[ 145 ][ 308 ],
   alphaCSR[ 145 ][ 309 ],
   alphaCSR[ 145 ][ 310 ],
   alphaCSR[ 145 ][ 311 ],
   alphaCSR[ 145 ][ 312 ],
   alphaCSR[ 145 ][ 313 ],
   alphaCSR[ 145 ][ 314 ],
   alphaCSR[ 145 ][ 315 ],
   alphaCSR[ 145 ][ 316 ],
   alphaCSR[ 145 ][ 317 ],
   alphaCSR[ 145 ][ 318 ],
   alphaCSR[ 145 ][ 319 ],
   alphaCSR[ 145 ][ 320 ],
   alphaCSR[ 145 ][ 321 ],
   alphaCSR[ 145 ][ 322 ],
   alphaCSR[ 145 ][ 323 ],
   alphaCSR[ 145 ][ 324 ],
   alphaCSR[ 145 ][ 325 ],
   alphaCSR[ 145 ][ 326 ],
   alphaCSR[ 145 ][ 327 ],
   alphaCSR[ 145 ][ 328 ],
   alphaCSR[ 145 ][ 329 ],
   alphaCSR[ 145 ][ 330 ],
   alphaCSR[ 145 ][ 331 ],
   alphaCSR[ 145 ][ 332 ],
   alphaCSR[ 145 ][ 333 ],
   alphaCSR[ 145 ][ 334 ],
   alphaCSR[ 145 ][ 335 ],
   alphaCSR[ 145 ][ 336 ],
   alphaCSR[ 145 ][ 337 ],
   alphaCSR[ 145 ][ 338 ],
   alphaCSR[ 145 ][ 339 ],
   alphaCSR[ 145 ][ 340 ],
   alphaCSR[ 145 ][ 341 ],
   alphaCSR[ 145 ][ 342 ],
   alphaCSR[ 145 ][ 343 ],
   alphaCSR[ 145 ][ 344 ],
   alphaCSR[ 145 ][ 345 ],
   alphaCSR[ 145 ][ 346 ],
   alphaCSR[ 145 ][ 347 ],
   alphaCSR[ 145 ][ 348 ],
   alphaCSR[ 145 ][ 349 ],
   alphaCSR[ 145 ][ 350 ],
   alphaCSR[ 145 ][ 351 ],
   alphaCSR[ 145 ][ 352 ],
   alphaCSR[ 145 ][ 353 ],
   alphaCSR[ 145 ][ 354 ],
   alphaCSR[ 145 ][ 355 ],
   alphaCSR[ 145 ][ 356 ],
   alphaCSR[ 145 ][ 357 ],
   alphaCSR[ 145 ][ 358 ],
   alphaCSR[ 145 ][ 359 ],
   alphaCSR[ 145 ][ 360 ],
   alphaCSR[ 145 ][ 361 ],
   alphaCSR[ 145 ][ 362 ],
   alphaCSR[ 145 ][ 363 ],
   alphaCSR[ 145 ][ 364 ],
   alphaCSR[ 145 ][ 365 ],
   alphaCSR[ 145 ][ 366 ],
   alphaCSR[ 145 ][ 367 ],
   alphaCSR[ 145 ][ 368 ],
   alphaCSR[ 145 ][ 369 ],
   alphaCSR[ 145 ][ 370 ],
   alphaCSR[ 145 ][ 371 ],
   alphaCSR[ 145 ][ 372 ],
   alphaCSR[ 145 ][ 373 ],
   alphaCSR[ 145 ][ 374 ],
   alphaCSR[ 145 ][ 375 ],
   alphaCSR[ 145 ][ 376 ],
   alphaCSR[ 145 ][ 377 ],
   alphaCSR[ 145 ][ 378 ],
   alphaCSR[ 145 ][ 379 ],
   alphaCSR[ 145 ][ 380 ],
   alphaCSR[ 145 ][ 381 ],
   alphaCSR[ 145 ][ 382 ],
   alphaCSR[ 145 ][ 383 ],
   alphaCSR[ 146 ][ 0 ],
   alphaCSR[ 146 ][ 1 ],
   alphaCSR[ 146 ][ 2 ],
   alphaCSR[ 146 ][ 3 ],
   alphaCSR[ 146 ][ 4 ],
   alphaCSR[ 146 ][ 5 ],
   alphaCSR[ 146 ][ 6 ],
   alphaCSR[ 146 ][ 7 ],
   alphaCSR[ 146 ][ 8 ],
   alphaCSR[ 146 ][ 9 ],
   alphaCSR[ 146 ][ 10 ],
   alphaCSR[ 146 ][ 11 ],
   alphaCSR[ 146 ][ 12 ],
   alphaCSR[ 146 ][ 13 ],
   alphaCSR[ 146 ][ 14 ],
   alphaCSR[ 146 ][ 15 ],
   alphaCSR[ 146 ][ 16 ],
   alphaCSR[ 146 ][ 17 ],
   alphaCSR[ 146 ][ 18 ],
   alphaCSR[ 146 ][ 19 ],
   alphaCSR[ 146 ][ 20 ],
   alphaCSR[ 146 ][ 21 ],
   alphaCSR[ 146 ][ 22 ],
   alphaCSR[ 146 ][ 23 ],
   alphaCSR[ 146 ][ 24 ],
   alphaCSR[ 146 ][ 25 ],
   alphaCSR[ 146 ][ 26 ],
   alphaCSR[ 146 ][ 27 ],
   alphaCSR[ 146 ][ 28 ],
   alphaCSR[ 146 ][ 29 ],
   alphaCSR[ 146 ][ 30 ],
   alphaCSR[ 146 ][ 31 ],
   alphaCSR[ 146 ][ 32 ],
   alphaCSR[ 146 ][ 33 ],
   alphaCSR[ 146 ][ 34 ],
   alphaCSR[ 146 ][ 35 ],
   alphaCSR[ 146 ][ 36 ],
   alphaCSR[ 146 ][ 37 ],
   alphaCSR[ 146 ][ 38 ],
   alphaCSR[ 146 ][ 39 ],
   alphaCSR[ 146 ][ 40 ],
   alphaCSR[ 146 ][ 41 ],
   alphaCSR[ 146 ][ 42 ],
   alphaCSR[ 146 ][ 43 ],
   alphaCSR[ 146 ][ 44 ],
   alphaCSR[ 146 ][ 45 ],
   alphaCSR[ 146 ][ 46 ],
   alphaCSR[ 146 ][ 47 ],
   alphaCSR[ 146 ][ 48 ],
   alphaCSR[ 146 ][ 49 ],
   alphaCSR[ 146 ][ 50 ],
   alphaCSR[ 146 ][ 51 ],
   alphaCSR[ 146 ][ 52 ],
   alphaCSR[ 146 ][ 53 ],
   alphaCSR[ 146 ][ 54 ],
   alphaCSR[ 146 ][ 55 ],
   alphaCSR[ 146 ][ 56 ],
   alphaCSR[ 146 ][ 57 ],
   alphaCSR[ 146 ][ 58 ],
   alphaCSR[ 146 ][ 59 ],
   alphaCSR[ 146 ][ 60 ],
   alphaCSR[ 146 ][ 61 ],
   alphaCSR[ 146 ][ 62 ],
   alphaCSR[ 146 ][ 63 ],
   alphaCSR[ 146 ][ 64 ],
   alphaCSR[ 146 ][ 65 ],
   alphaCSR[ 146 ][ 66 ],
   alphaCSR[ 146 ][ 67 ],
   alphaCSR[ 146 ][ 68 ],
   alphaCSR[ 146 ][ 69 ],
   alphaCSR[ 146 ][ 70 ],
   alphaCSR[ 146 ][ 71 ],
   alphaCSR[ 146 ][ 72 ],
   alphaCSR[ 146 ][ 73 ],
   alphaCSR[ 146 ][ 74 ],
   alphaCSR[ 146 ][ 75 ],
   alphaCSR[ 146 ][ 76 ],
   alphaCSR[ 146 ][ 77 ],
   alphaCSR[ 146 ][ 78 ],
   alphaCSR[ 146 ][ 79 ],
   alphaCSR[ 146 ][ 80 ],
   alphaCSR[ 146 ][ 81 ],
   alphaCSR[ 146 ][ 82 ],
   alphaCSR[ 146 ][ 83 ],
   alphaCSR[ 146 ][ 84 ],
   alphaCSR[ 146 ][ 85 ],
   alphaCSR[ 146 ][ 86 ],
   alphaCSR[ 146 ][ 87 ],
   alphaCSR[ 146 ][ 88 ],
   alphaCSR[ 146 ][ 89 ],
   alphaCSR[ 146 ][ 90 ],
   alphaCSR[ 146 ][ 91 ],
   alphaCSR[ 146 ][ 92 ],
   alphaCSR[ 146 ][ 93 ],
   alphaCSR[ 146 ][ 94 ],
   alphaCSR[ 146 ][ 95 ],
   alphaCSR[ 146 ][ 96 ],
   alphaCSR[ 146 ][ 97 ],
   alphaCSR[ 146 ][ 98 ],
   alphaCSR[ 146 ][ 99 ],
   alphaCSR[ 146 ][ 100 ],
   alphaCSR[ 146 ][ 101 ],
   alphaCSR[ 146 ][ 102 ],
   alphaCSR[ 146 ][ 103 ],
   alphaCSR[ 146 ][ 104 ],
   alphaCSR[ 146 ][ 105 ],
   alphaCSR[ 146 ][ 106 ],
   alphaCSR[ 146 ][ 107 ],
   alphaCSR[ 146 ][ 108 ],
   alphaCSR[ 146 ][ 109 ],
   alphaCSR[ 146 ][ 110 ],
   alphaCSR[ 146 ][ 111 ],
   alphaCSR[ 146 ][ 112 ],
   alphaCSR[ 146 ][ 113 ],
   alphaCSR[ 146 ][ 114 ],
   alphaCSR[ 146 ][ 115 ],
   alphaCSR[ 146 ][ 116 ],
   alphaCSR[ 146 ][ 117 ],
   alphaCSR[ 146 ][ 118 ],
   alphaCSR[ 146 ][ 119 ],
   alphaCSR[ 146 ][ 120 ],
   alphaCSR[ 146 ][ 121 ],
   alphaCSR[ 146 ][ 122 ],
   alphaCSR[ 146 ][ 123 ],
   alphaCSR[ 146 ][ 124 ],
   alphaCSR[ 146 ][ 125 ],
   alphaCSR[ 146 ][ 126 ],
   alphaCSR[ 146 ][ 127 ],
   alphaCSR[ 146 ][ 128 ],
   alphaCSR[ 146 ][ 129 ],
   alphaCSR[ 146 ][ 130 ],
   alphaCSR[ 146 ][ 131 ],
   alphaCSR[ 146 ][ 132 ],
   alphaCSR[ 146 ][ 133 ],
   alphaCSR[ 146 ][ 134 ],
   alphaCSR[ 146 ][ 135 ],
   alphaCSR[ 146 ][ 136 ],
   alphaCSR[ 146 ][ 137 ],
   alphaCSR[ 146 ][ 138 ],
   alphaCSR[ 146 ][ 139 ],
   alphaCSR[ 146 ][ 140 ],
   alphaCSR[ 146 ][ 141 ],
   alphaCSR[ 146 ][ 142 ],
   alphaCSR[ 146 ][ 143 ],
   alphaCSR[ 146 ][ 144 ],
   alphaCSR[ 146 ][ 145 ],
   alphaCSR[ 146 ][ 146 ],
   alphaCSR[ 146 ][ 147 ],
   alphaCSR[ 146 ][ 148 ],
   alphaCSR[ 146 ][ 149 ],
   alphaCSR[ 146 ][ 150 ],
   alphaCSR[ 146 ][ 151 ],
   alphaCSR[ 146 ][ 152 ],
   alphaCSR[ 146 ][ 153 ],
   alphaCSR[ 146 ][ 154 ],
   alphaCSR[ 146 ][ 155 ],
   alphaCSR[ 146 ][ 156 ],
   alphaCSR[ 146 ][ 157 ],
   alphaCSR[ 146 ][ 158 ],
   alphaCSR[ 146 ][ 159 ],
   alphaCSR[ 146 ][ 160 ],
   alphaCSR[ 146 ][ 161 ],
   alphaCSR[ 146 ][ 162 ],
   alphaCSR[ 146 ][ 163 ],
   alphaCSR[ 146 ][ 164 ],
   alphaCSR[ 146 ][ 165 ],
   alphaCSR[ 146 ][ 166 ],
   alphaCSR[ 146 ][ 167 ],
   alphaCSR[ 146 ][ 168 ],
   alphaCSR[ 146 ][ 169 ],
   alphaCSR[ 146 ][ 170 ],
   alphaCSR[ 146 ][ 171 ],
   alphaCSR[ 146 ][ 172 ],
   alphaCSR[ 146 ][ 173 ],
   alphaCSR[ 146 ][ 174 ],
   alphaCSR[ 146 ][ 175 ],
   alphaCSR[ 146 ][ 176 ],
   alphaCSR[ 146 ][ 177 ],
   alphaCSR[ 146 ][ 178 ],
   alphaCSR[ 146 ][ 179 ],
   alphaCSR[ 146 ][ 180 ],
   alphaCSR[ 146 ][ 181 ],
   alphaCSR[ 146 ][ 182 ],
   alphaCSR[ 146 ][ 183 ],
   alphaCSR[ 146 ][ 184 ],
   alphaCSR[ 146 ][ 185 ],
   alphaCSR[ 146 ][ 186 ],
   alphaCSR[ 146 ][ 187 ],
   alphaCSR[ 146 ][ 188 ],
   alphaCSR[ 146 ][ 189 ],
   alphaCSR[ 146 ][ 190 ],
   alphaCSR[ 146 ][ 191 ],
   alphaCSR[ 146 ][ 192 ],
   alphaCSR[ 146 ][ 193 ],
   alphaCSR[ 146 ][ 194 ],
   alphaCSR[ 146 ][ 195 ],
   alphaCSR[ 146 ][ 196 ],
   alphaCSR[ 146 ][ 197 ],
   alphaCSR[ 146 ][ 198 ],
   alphaCSR[ 146 ][ 199 ],
   alphaCSR[ 146 ][ 200 ],
   alphaCSR[ 146 ][ 201 ],
   alphaCSR[ 146 ][ 202 ],
   alphaCSR[ 146 ][ 203 ],
   alphaCSR[ 146 ][ 204 ],
   alphaCSR[ 146 ][ 205 ],
   alphaCSR[ 146 ][ 206 ],
   alphaCSR[ 146 ][ 207 ],
   alphaCSR[ 146 ][ 208 ],
   alphaCSR[ 146 ][ 209 ],
   alphaCSR[ 146 ][ 210 ],
   alphaCSR[ 146 ][ 211 ],
   alphaCSR[ 146 ][ 212 ],
   alphaCSR[ 146 ][ 213 ],
   alphaCSR[ 146 ][ 214 ],
   alphaCSR[ 146 ][ 215 ],
   alphaCSR[ 146 ][ 216 ],
   alphaCSR[ 146 ][ 217 ],
   alphaCSR[ 146 ][ 218 ],
   alphaCSR[ 146 ][ 219 ],
   alphaCSR[ 146 ][ 220 ],
   alphaCSR[ 146 ][ 221 ],
   alphaCSR[ 146 ][ 222 ],
   alphaCSR[ 146 ][ 223 ],
   alphaCSR[ 146 ][ 224 ],
   alphaCSR[ 146 ][ 225 ],
   alphaCSR[ 146 ][ 226 ],
   alphaCSR[ 146 ][ 227 ],
   alphaCSR[ 146 ][ 228 ],
   alphaCSR[ 146 ][ 229 ],
   alphaCSR[ 146 ][ 230 ],
   alphaCSR[ 146 ][ 231 ],
   alphaCSR[ 146 ][ 232 ],
   alphaCSR[ 146 ][ 233 ],
   alphaCSR[ 146 ][ 234 ],
   alphaCSR[ 146 ][ 235 ],
   alphaCSR[ 146 ][ 236 ],
   alphaCSR[ 146 ][ 237 ],
   alphaCSR[ 146 ][ 238 ],
   alphaCSR[ 146 ][ 239 ],
   alphaCSR[ 146 ][ 240 ],
   alphaCSR[ 146 ][ 241 ],
   alphaCSR[ 146 ][ 242 ],
   alphaCSR[ 146 ][ 243 ],
   alphaCSR[ 146 ][ 244 ],
   alphaCSR[ 146 ][ 245 ],
   alphaCSR[ 146 ][ 246 ],
   alphaCSR[ 146 ][ 247 ],
   alphaCSR[ 146 ][ 248 ],
   alphaCSR[ 146 ][ 249 ],
   alphaCSR[ 146 ][ 250 ],
   alphaCSR[ 146 ][ 251 ],
   alphaCSR[ 146 ][ 252 ],
   alphaCSR[ 146 ][ 253 ],
   alphaCSR[ 146 ][ 254 ],
   alphaCSR[ 146 ][ 255 ],
   alphaCSR[ 146 ][ 256 ],
   alphaCSR[ 146 ][ 257 ],
   alphaCSR[ 146 ][ 258 ],
   alphaCSR[ 146 ][ 259 ],
   alphaCSR[ 146 ][ 260 ],
   alphaCSR[ 146 ][ 261 ],
   alphaCSR[ 146 ][ 262 ],
   alphaCSR[ 146 ][ 263 ],
   alphaCSR[ 146 ][ 264 ],
   alphaCSR[ 146 ][ 265 ],
   alphaCSR[ 146 ][ 266 ],
   alphaCSR[ 146 ][ 267 ],
   alphaCSR[ 146 ][ 268 ],
   alphaCSR[ 146 ][ 269 ],
   alphaCSR[ 146 ][ 270 ],
   alphaCSR[ 146 ][ 271 ],
   alphaCSR[ 146 ][ 272 ],
   alphaCSR[ 146 ][ 273 ],
   alphaCSR[ 146 ][ 274 ],
   alphaCSR[ 146 ][ 275 ],
   alphaCSR[ 146 ][ 276 ],
   alphaCSR[ 146 ][ 277 ],
   alphaCSR[ 146 ][ 278 ],
   alphaCSR[ 146 ][ 279 ],
   alphaCSR[ 146 ][ 280 ],
   alphaCSR[ 146 ][ 281 ],
   alphaCSR[ 146 ][ 282 ],
   alphaCSR[ 146 ][ 283 ],
   alphaCSR[ 146 ][ 284 ],
   alphaCSR[ 146 ][ 285 ],
   alphaCSR[ 146 ][ 286 ],
   alphaCSR[ 146 ][ 287 ],
   alphaCSR[ 146 ][ 288 ],
   alphaCSR[ 146 ][ 289 ],
   alphaCSR[ 146 ][ 290 ],
   alphaCSR[ 146 ][ 291 ],
   alphaCSR[ 146 ][ 292 ],
   alphaCSR[ 146 ][ 293 ],
   alphaCSR[ 146 ][ 294 ],
   alphaCSR[ 146 ][ 295 ],
   alphaCSR[ 146 ][ 296 ],
   alphaCSR[ 146 ][ 297 ],
   alphaCSR[ 146 ][ 298 ],
   alphaCSR[ 146 ][ 299 ],
   alphaCSR[ 146 ][ 300 ],
   alphaCSR[ 146 ][ 301 ],
   alphaCSR[ 146 ][ 302 ],
   alphaCSR[ 146 ][ 303 ],
   alphaCSR[ 146 ][ 304 ],
   alphaCSR[ 146 ][ 305 ],
   alphaCSR[ 146 ][ 306 ],
   alphaCSR[ 146 ][ 307 ],
   alphaCSR[ 146 ][ 308 ],
   alphaCSR[ 146 ][ 309 ],
   alphaCSR[ 146 ][ 310 ],
   alphaCSR[ 146 ][ 311 ],
   alphaCSR[ 146 ][ 312 ],
   alphaCSR[ 146 ][ 313 ],
   alphaCSR[ 146 ][ 314 ],
   alphaCSR[ 146 ][ 315 ],
   alphaCSR[ 146 ][ 316 ],
   alphaCSR[ 146 ][ 317 ],
   alphaCSR[ 146 ][ 318 ],
   alphaCSR[ 146 ][ 319 ],
   alphaCSR[ 146 ][ 320 ],
   alphaCSR[ 146 ][ 321 ],
   alphaCSR[ 146 ][ 322 ],
   alphaCSR[ 146 ][ 323 ],
   alphaCSR[ 146 ][ 324 ],
   alphaCSR[ 146 ][ 325 ],
   alphaCSR[ 146 ][ 326 ],
   alphaCSR[ 146 ][ 327 ],
   alphaCSR[ 146 ][ 328 ],
   alphaCSR[ 146 ][ 329 ],
   alphaCSR[ 146 ][ 330 ],
   alphaCSR[ 146 ][ 331 ],
   alphaCSR[ 146 ][ 332 ],
   alphaCSR[ 146 ][ 333 ],
   alphaCSR[ 146 ][ 334 ],
   alphaCSR[ 146 ][ 335 ],
   alphaCSR[ 146 ][ 336 ],
   alphaCSR[ 146 ][ 337 ],
   alphaCSR[ 146 ][ 338 ],
   alphaCSR[ 146 ][ 339 ],
   alphaCSR[ 146 ][ 340 ],
   alphaCSR[ 146 ][ 341 ],
   alphaCSR[ 146 ][ 342 ],
   alphaCSR[ 146 ][ 343 ],
   alphaCSR[ 146 ][ 344 ],
   alphaCSR[ 146 ][ 345 ],
   alphaCSR[ 146 ][ 346 ],
   alphaCSR[ 146 ][ 347 ],
   alphaCSR[ 146 ][ 348 ],
   alphaCSR[ 146 ][ 349 ],
   alphaCSR[ 146 ][ 350 ],
   alphaCSR[ 146 ][ 351 ],
   alphaCSR[ 146 ][ 352 ],
   alphaCSR[ 146 ][ 353 ],
   alphaCSR[ 146 ][ 354 ],
   alphaCSR[ 146 ][ 355 ],
   alphaCSR[ 146 ][ 356 ],
   alphaCSR[ 146 ][ 357 ],
   alphaCSR[ 146 ][ 358 ],
   alphaCSR[ 146 ][ 359 ],
   alphaCSR[ 146 ][ 360 ],
   alphaCSR[ 146 ][ 361 ],
   alphaCSR[ 146 ][ 362 ],
   alphaCSR[ 146 ][ 363 ],
   alphaCSR[ 146 ][ 364 ],
   alphaCSR[ 146 ][ 365 ],
   alphaCSR[ 146 ][ 366 ],
   alphaCSR[ 146 ][ 367 ],
   alphaCSR[ 146 ][ 368 ],
   alphaCSR[ 146 ][ 369 ],
   alphaCSR[ 146 ][ 370 ],
   alphaCSR[ 146 ][ 371 ],
   alphaCSR[ 146 ][ 372 ],
   alphaCSR[ 146 ][ 373 ],
   alphaCSR[ 146 ][ 374 ],
   alphaCSR[ 146 ][ 375 ],
   alphaCSR[ 146 ][ 376 ],
   alphaCSR[ 146 ][ 377 ],
   alphaCSR[ 146 ][ 378 ],
   alphaCSR[ 146 ][ 379 ],
   alphaCSR[ 146 ][ 380 ],
   alphaCSR[ 146 ][ 381 ],
   alphaCSR[ 146 ][ 382 ],
   alphaCSR[ 146 ][ 383 ],
   alphaCSR[ 147 ][ 0 ],
   alphaCSR[ 147 ][ 1 ],
   alphaCSR[ 147 ][ 2 ],
   alphaCSR[ 147 ][ 3 ],
   alphaCSR[ 147 ][ 4 ],
   alphaCSR[ 147 ][ 5 ],
   alphaCSR[ 147 ][ 6 ],
   alphaCSR[ 147 ][ 7 ],
   alphaCSR[ 147 ][ 8 ],
   alphaCSR[ 147 ][ 9 ],
   alphaCSR[ 147 ][ 10 ],
   alphaCSR[ 147 ][ 11 ],
   alphaCSR[ 147 ][ 12 ],
   alphaCSR[ 147 ][ 13 ],
   alphaCSR[ 147 ][ 14 ],
   alphaCSR[ 147 ][ 15 ],
   alphaCSR[ 147 ][ 16 ],
   alphaCSR[ 147 ][ 17 ],
   alphaCSR[ 147 ][ 18 ],
   alphaCSR[ 147 ][ 19 ],
   alphaCSR[ 147 ][ 20 ],
   alphaCSR[ 147 ][ 21 ],
   alphaCSR[ 147 ][ 22 ],
   alphaCSR[ 147 ][ 23 ],
   alphaCSR[ 147 ][ 24 ],
   alphaCSR[ 147 ][ 25 ],
   alphaCSR[ 147 ][ 26 ],
   alphaCSR[ 147 ][ 27 ],
   alphaCSR[ 147 ][ 28 ],
   alphaCSR[ 147 ][ 29 ],
   alphaCSR[ 147 ][ 30 ],
   alphaCSR[ 147 ][ 31 ],
   alphaCSR[ 147 ][ 32 ],
   alphaCSR[ 147 ][ 33 ],
   alphaCSR[ 147 ][ 34 ],
   alphaCSR[ 147 ][ 35 ],
   alphaCSR[ 147 ][ 36 ],
   alphaCSR[ 147 ][ 37 ],
   alphaCSR[ 147 ][ 38 ],
   alphaCSR[ 147 ][ 39 ],
   alphaCSR[ 147 ][ 40 ],
   alphaCSR[ 147 ][ 41 ],
   alphaCSR[ 147 ][ 42 ],
   alphaCSR[ 147 ][ 43 ],
   alphaCSR[ 147 ][ 44 ],
   alphaCSR[ 147 ][ 45 ],
   alphaCSR[ 147 ][ 46 ],
   alphaCSR[ 147 ][ 47 ],
   alphaCSR[ 147 ][ 48 ],
   alphaCSR[ 147 ][ 49 ],
   alphaCSR[ 147 ][ 50 ],
   alphaCSR[ 147 ][ 51 ],
   alphaCSR[ 147 ][ 52 ],
   alphaCSR[ 147 ][ 53 ],
   alphaCSR[ 147 ][ 54 ],
   alphaCSR[ 147 ][ 55 ],
   alphaCSR[ 147 ][ 56 ],
   alphaCSR[ 147 ][ 57 ],
   alphaCSR[ 147 ][ 58 ],
   alphaCSR[ 147 ][ 59 ],
   alphaCSR[ 147 ][ 60 ],
   alphaCSR[ 147 ][ 61 ],
   alphaCSR[ 147 ][ 62 ],
   alphaCSR[ 147 ][ 63 ],
   alphaCSR[ 147 ][ 64 ],
   alphaCSR[ 147 ][ 65 ],
   alphaCSR[ 147 ][ 66 ],
   alphaCSR[ 147 ][ 67 ],
   alphaCSR[ 147 ][ 68 ],
   alphaCSR[ 147 ][ 69 ],
   alphaCSR[ 147 ][ 70 ],
   alphaCSR[ 147 ][ 71 ],
   alphaCSR[ 147 ][ 72 ],
   alphaCSR[ 147 ][ 73 ],
   alphaCSR[ 147 ][ 74 ],
   alphaCSR[ 147 ][ 75 ],
   alphaCSR[ 147 ][ 76 ],
   alphaCSR[ 147 ][ 77 ],
   alphaCSR[ 147 ][ 78 ],
   alphaCSR[ 147 ][ 79 ],
   alphaCSR[ 147 ][ 80 ],
   alphaCSR[ 147 ][ 81 ],
   alphaCSR[ 147 ][ 82 ],
   alphaCSR[ 147 ][ 83 ],
   alphaCSR[ 147 ][ 84 ],
   alphaCSR[ 147 ][ 85 ],
   alphaCSR[ 147 ][ 86 ],
   alphaCSR[ 147 ][ 87 ],
   alphaCSR[ 147 ][ 88 ],
   alphaCSR[ 147 ][ 89 ],
   alphaCSR[ 147 ][ 90 ],
   alphaCSR[ 147 ][ 91 ],
   alphaCSR[ 147 ][ 92 ],
   alphaCSR[ 147 ][ 93 ],
   alphaCSR[ 147 ][ 94 ],
   alphaCSR[ 147 ][ 95 ],
   alphaCSR[ 147 ][ 96 ],
   alphaCSR[ 147 ][ 97 ],
   alphaCSR[ 147 ][ 98 ],
   alphaCSR[ 147 ][ 99 ],
   alphaCSR[ 147 ][ 100 ],
   alphaCSR[ 147 ][ 101 ],
   alphaCSR[ 147 ][ 102 ],
   alphaCSR[ 147 ][ 103 ],
   alphaCSR[ 147 ][ 104 ],
   alphaCSR[ 147 ][ 105 ],
   alphaCSR[ 147 ][ 106 ],
   alphaCSR[ 147 ][ 107 ],
   alphaCSR[ 147 ][ 108 ],
   alphaCSR[ 147 ][ 109 ],
   alphaCSR[ 147 ][ 110 ],
   alphaCSR[ 147 ][ 111 ],
   alphaCSR[ 147 ][ 112 ],
   alphaCSR[ 147 ][ 113 ],
   alphaCSR[ 147 ][ 114 ],
   alphaCSR[ 147 ][ 115 ],
   alphaCSR[ 147 ][ 116 ],
   alphaCSR[ 147 ][ 117 ],
   alphaCSR[ 147 ][ 118 ],
   alphaCSR[ 147 ][ 119 ],
   alphaCSR[ 147 ][ 120 ],
   alphaCSR[ 147 ][ 121 ],
   alphaCSR[ 147 ][ 122 ],
   alphaCSR[ 147 ][ 123 ],
   alphaCSR[ 147 ][ 124 ],
   alphaCSR[ 147 ][ 125 ],
   alphaCSR[ 147 ][ 126 ],
   alphaCSR[ 147 ][ 127 ],
   alphaCSR[ 147 ][ 128 ],
   alphaCSR[ 147 ][ 129 ],
   alphaCSR[ 147 ][ 130 ],
   alphaCSR[ 147 ][ 131 ],
   alphaCSR[ 147 ][ 132 ],
   alphaCSR[ 147 ][ 133 ],
   alphaCSR[ 147 ][ 134 ],
   alphaCSR[ 147 ][ 135 ],
   alphaCSR[ 147 ][ 136 ],
   alphaCSR[ 147 ][ 137 ],
   alphaCSR[ 147 ][ 138 ],
   alphaCSR[ 147 ][ 139 ],
   alphaCSR[ 147 ][ 140 ],
   alphaCSR[ 147 ][ 141 ],
   alphaCSR[ 147 ][ 142 ],
   alphaCSR[ 147 ][ 143 ],
   alphaCSR[ 147 ][ 144 ],
   alphaCSR[ 147 ][ 145 ],
   alphaCSR[ 147 ][ 146 ],
   alphaCSR[ 147 ][ 147 ],
   alphaCSR[ 147 ][ 148 ],
   alphaCSR[ 147 ][ 149 ],
   alphaCSR[ 147 ][ 150 ],
   alphaCSR[ 147 ][ 151 ],
   alphaCSR[ 147 ][ 152 ],
   alphaCSR[ 147 ][ 153 ],
   alphaCSR[ 147 ][ 154 ],
   alphaCSR[ 147 ][ 155 ],
   alphaCSR[ 147 ][ 156 ],
   alphaCSR[ 147 ][ 157 ],
   alphaCSR[ 147 ][ 158 ],
   alphaCSR[ 147 ][ 159 ],
   alphaCSR[ 147 ][ 160 ],
   alphaCSR[ 147 ][ 161 ],
   alphaCSR[ 147 ][ 162 ],
   alphaCSR[ 147 ][ 163 ],
   alphaCSR[ 147 ][ 164 ],
   alphaCSR[ 147 ][ 165 ],
   alphaCSR[ 147 ][ 166 ],
   alphaCSR[ 147 ][ 167 ],
   alphaCSR[ 147 ][ 168 ],
   alphaCSR[ 147 ][ 169 ],
   alphaCSR[ 147 ][ 170 ],
   alphaCSR[ 147 ][ 171 ],
   alphaCSR[ 147 ][ 172 ],
   alphaCSR[ 147 ][ 173 ],
   alphaCSR[ 147 ][ 174 ],
   alphaCSR[ 147 ][ 175 ],
   alphaCSR[ 147 ][ 176 ],
   alphaCSR[ 147 ][ 177 ],
   alphaCSR[ 147 ][ 178 ],
   alphaCSR[ 147 ][ 179 ],
   alphaCSR[ 147 ][ 180 ],
   alphaCSR[ 147 ][ 181 ],
   alphaCSR[ 147 ][ 182 ],
   alphaCSR[ 147 ][ 183 ],
   alphaCSR[ 147 ][ 184 ],
   alphaCSR[ 147 ][ 185 ],
   alphaCSR[ 147 ][ 186 ],
   alphaCSR[ 147 ][ 187 ],
   alphaCSR[ 147 ][ 188 ],
   alphaCSR[ 147 ][ 189 ],
   alphaCSR[ 147 ][ 190 ],
   alphaCSR[ 147 ][ 191 ],
   alphaCSR[ 147 ][ 192 ],
   alphaCSR[ 147 ][ 193 ],
   alphaCSR[ 147 ][ 194 ],
   alphaCSR[ 147 ][ 195 ],
   alphaCSR[ 147 ][ 196 ],
   alphaCSR[ 147 ][ 197 ],
   alphaCSR[ 147 ][ 198 ],
   alphaCSR[ 147 ][ 199 ],
   alphaCSR[ 147 ][ 200 ],
   alphaCSR[ 147 ][ 201 ],
   alphaCSR[ 147 ][ 202 ],
   alphaCSR[ 147 ][ 203 ],
   alphaCSR[ 147 ][ 204 ],
   alphaCSR[ 147 ][ 205 ],
   alphaCSR[ 147 ][ 206 ],
   alphaCSR[ 147 ][ 207 ],
   alphaCSR[ 147 ][ 208 ],
   alphaCSR[ 147 ][ 209 ],
   alphaCSR[ 147 ][ 210 ],
   alphaCSR[ 147 ][ 211 ],
   alphaCSR[ 147 ][ 212 ],
   alphaCSR[ 147 ][ 213 ],
   alphaCSR[ 147 ][ 214 ],
   alphaCSR[ 147 ][ 215 ],
   alphaCSR[ 147 ][ 216 ],
   alphaCSR[ 147 ][ 217 ],
   alphaCSR[ 147 ][ 218 ],
   alphaCSR[ 147 ][ 219 ],
   alphaCSR[ 147 ][ 220 ],
   alphaCSR[ 147 ][ 221 ],
   alphaCSR[ 147 ][ 222 ],
   alphaCSR[ 147 ][ 223 ],
   alphaCSR[ 147 ][ 224 ],
   alphaCSR[ 147 ][ 225 ],
   alphaCSR[ 147 ][ 226 ],
   alphaCSR[ 147 ][ 227 ],
   alphaCSR[ 147 ][ 228 ],
   alphaCSR[ 147 ][ 229 ],
   alphaCSR[ 147 ][ 230 ],
   alphaCSR[ 147 ][ 231 ],
   alphaCSR[ 147 ][ 232 ],
   alphaCSR[ 147 ][ 233 ],
   alphaCSR[ 147 ][ 234 ],
   alphaCSR[ 147 ][ 235 ],
   alphaCSR[ 147 ][ 236 ],
   alphaCSR[ 147 ][ 237 ],
   alphaCSR[ 147 ][ 238 ],
   alphaCSR[ 147 ][ 239 ],
   alphaCSR[ 147 ][ 240 ],
   alphaCSR[ 147 ][ 241 ],
   alphaCSR[ 147 ][ 242 ],
   alphaCSR[ 147 ][ 243 ],
   alphaCSR[ 147 ][ 244 ],
   alphaCSR[ 147 ][ 245 ],
   alphaCSR[ 147 ][ 246 ],
   alphaCSR[ 147 ][ 247 ],
   alphaCSR[ 147 ][ 248 ],
   alphaCSR[ 147 ][ 249 ],
   alphaCSR[ 147 ][ 250 ],
   alphaCSR[ 147 ][ 251 ],
   alphaCSR[ 147 ][ 252 ],
   alphaCSR[ 147 ][ 253 ],
   alphaCSR[ 147 ][ 254 ],
   alphaCSR[ 147 ][ 255 ],
   alphaCSR[ 147 ][ 256 ],
   alphaCSR[ 147 ][ 257 ],
   alphaCSR[ 147 ][ 258 ],
   alphaCSR[ 147 ][ 259 ],
   alphaCSR[ 147 ][ 260 ],
   alphaCSR[ 147 ][ 261 ],
   alphaCSR[ 147 ][ 262 ],
   alphaCSR[ 147 ][ 263 ],
   alphaCSR[ 147 ][ 264 ],
   alphaCSR[ 147 ][ 265 ],
   alphaCSR[ 147 ][ 266 ],
   alphaCSR[ 147 ][ 267 ],
   alphaCSR[ 147 ][ 268 ],
   alphaCSR[ 147 ][ 269 ],
   alphaCSR[ 147 ][ 270 ],
   alphaCSR[ 147 ][ 271 ],
   alphaCSR[ 147 ][ 272 ],
   alphaCSR[ 147 ][ 273 ],
   alphaCSR[ 147 ][ 274 ],
   alphaCSR[ 147 ][ 275 ],
   alphaCSR[ 147 ][ 276 ],
   alphaCSR[ 147 ][ 277 ],
   alphaCSR[ 147 ][ 278 ],
   alphaCSR[ 147 ][ 279 ],
   alphaCSR[ 147 ][ 280 ],
   alphaCSR[ 147 ][ 281 ],
   alphaCSR[ 147 ][ 282 ],
   alphaCSR[ 147 ][ 283 ],
   alphaCSR[ 147 ][ 284 ],
   alphaCSR[ 147 ][ 285 ],
   alphaCSR[ 147 ][ 286 ],
   alphaCSR[ 147 ][ 287 ],
   alphaCSR[ 147 ][ 288 ],
   alphaCSR[ 147 ][ 289 ],
   alphaCSR[ 147 ][ 290 ],
   alphaCSR[ 147 ][ 291 ],
   alphaCSR[ 147 ][ 292 ],
   alphaCSR[ 147 ][ 293 ],
   alphaCSR[ 147 ][ 294 ],
   alphaCSR[ 147 ][ 295 ],
   alphaCSR[ 147 ][ 296 ],
   alphaCSR[ 147 ][ 297 ],
   alphaCSR[ 147 ][ 298 ],
   alphaCSR[ 147 ][ 299 ],
   alphaCSR[ 147 ][ 300 ],
   alphaCSR[ 147 ][ 301 ],
   alphaCSR[ 147 ][ 302 ],
   alphaCSR[ 147 ][ 303 ],
   alphaCSR[ 147 ][ 304 ],
   alphaCSR[ 147 ][ 305 ],
   alphaCSR[ 147 ][ 306 ],
   alphaCSR[ 147 ][ 307 ],
   alphaCSR[ 147 ][ 308 ],
   alphaCSR[ 147 ][ 309 ],
   alphaCSR[ 147 ][ 310 ],
   alphaCSR[ 147 ][ 311 ],
   alphaCSR[ 147 ][ 312 ],
   alphaCSR[ 147 ][ 313 ],
   alphaCSR[ 147 ][ 314 ],
   alphaCSR[ 147 ][ 315 ],
   alphaCSR[ 147 ][ 316 ],
   alphaCSR[ 147 ][ 317 ],
   alphaCSR[ 147 ][ 318 ],
   alphaCSR[ 147 ][ 319 ],
   alphaCSR[ 147 ][ 320 ],
   alphaCSR[ 147 ][ 321 ],
   alphaCSR[ 147 ][ 322 ],
   alphaCSR[ 147 ][ 323 ],
   alphaCSR[ 147 ][ 324 ],
   alphaCSR[ 147 ][ 325 ],
   alphaCSR[ 147 ][ 326 ],
   alphaCSR[ 147 ][ 327 ],
   alphaCSR[ 147 ][ 328 ],
   alphaCSR[ 147 ][ 329 ],
   alphaCSR[ 147 ][ 330 ],
   alphaCSR[ 147 ][ 331 ],
   alphaCSR[ 147 ][ 332 ],
   alphaCSR[ 147 ][ 333 ],
   alphaCSR[ 147 ][ 334 ],
   alphaCSR[ 147 ][ 335 ],
   alphaCSR[ 147 ][ 336 ],
   alphaCSR[ 147 ][ 337 ],
   alphaCSR[ 147 ][ 338 ],
   alphaCSR[ 147 ][ 339 ],
   alphaCSR[ 147 ][ 340 ],
   alphaCSR[ 147 ][ 341 ],
   alphaCSR[ 147 ][ 342 ],
   alphaCSR[ 147 ][ 343 ],
   alphaCSR[ 147 ][ 344 ],
   alphaCSR[ 147 ][ 345 ],
   alphaCSR[ 147 ][ 346 ],
   alphaCSR[ 147 ][ 347 ],
   alphaCSR[ 147 ][ 348 ],
   alphaCSR[ 147 ][ 349 ],
   alphaCSR[ 147 ][ 350 ],
   alphaCSR[ 147 ][ 351 ],
   alphaCSR[ 147 ][ 352 ],
   alphaCSR[ 147 ][ 353 ],
   alphaCSR[ 147 ][ 354 ],
   alphaCSR[ 147 ][ 355 ],
   alphaCSR[ 147 ][ 356 ],
   alphaCSR[ 147 ][ 357 ],
   alphaCSR[ 147 ][ 358 ],
   alphaCSR[ 147 ][ 359 ],
   alphaCSR[ 147 ][ 360 ],
   alphaCSR[ 147 ][ 361 ],
   alphaCSR[ 147 ][ 362 ],
   alphaCSR[ 147 ][ 363 ],
   alphaCSR[ 147 ][ 364 ],
   alphaCSR[ 147 ][ 365 ],
   alphaCSR[ 147 ][ 366 ],
   alphaCSR[ 147 ][ 367 ],
   alphaCSR[ 147 ][ 368 ],
   alphaCSR[ 147 ][ 369 ],
   alphaCSR[ 147 ][ 370 ],
   alphaCSR[ 147 ][ 371 ],
   alphaCSR[ 147 ][ 372 ],
   alphaCSR[ 147 ][ 373 ],
   alphaCSR[ 147 ][ 374 ],
   alphaCSR[ 147 ][ 375 ],
   alphaCSR[ 147 ][ 376 ],
   alphaCSR[ 147 ][ 377 ],
   alphaCSR[ 147 ][ 378 ],
   alphaCSR[ 147 ][ 379 ],
   alphaCSR[ 147 ][ 380 ],
   alphaCSR[ 147 ][ 381 ],
   alphaCSR[ 147 ][ 382 ],
   alphaCSR[ 147 ][ 383 ],
   alphaCSR[ 148 ][ 0 ],
   alphaCSR[ 148 ][ 1 ],
   alphaCSR[ 148 ][ 2 ],
   alphaCSR[ 148 ][ 3 ],
   alphaCSR[ 148 ][ 4 ],
   alphaCSR[ 148 ][ 5 ],
   alphaCSR[ 148 ][ 6 ],
   alphaCSR[ 148 ][ 7 ],
   alphaCSR[ 148 ][ 8 ],
   alphaCSR[ 148 ][ 9 ],
   alphaCSR[ 148 ][ 10 ],
   alphaCSR[ 148 ][ 11 ],
   alphaCSR[ 148 ][ 12 ],
   alphaCSR[ 148 ][ 13 ],
   alphaCSR[ 148 ][ 14 ],
   alphaCSR[ 148 ][ 15 ],
   alphaCSR[ 148 ][ 16 ],
   alphaCSR[ 148 ][ 17 ],
   alphaCSR[ 148 ][ 18 ],
   alphaCSR[ 148 ][ 19 ],
   alphaCSR[ 148 ][ 20 ],
   alphaCSR[ 148 ][ 21 ],
   alphaCSR[ 148 ][ 22 ],
   alphaCSR[ 148 ][ 23 ],
   alphaCSR[ 148 ][ 24 ],
   alphaCSR[ 148 ][ 25 ],
   alphaCSR[ 148 ][ 26 ],
   alphaCSR[ 148 ][ 27 ],
   alphaCSR[ 148 ][ 28 ],
   alphaCSR[ 148 ][ 29 ],
   alphaCSR[ 148 ][ 30 ],
   alphaCSR[ 148 ][ 31 ],
   alphaCSR[ 148 ][ 32 ],
   alphaCSR[ 148 ][ 33 ],
   alphaCSR[ 148 ][ 34 ],
   alphaCSR[ 148 ][ 35 ],
   alphaCSR[ 148 ][ 36 ],
   alphaCSR[ 148 ][ 37 ],
   alphaCSR[ 148 ][ 38 ],
   alphaCSR[ 148 ][ 39 ],
   alphaCSR[ 148 ][ 40 ],
   alphaCSR[ 148 ][ 41 ],
   alphaCSR[ 148 ][ 42 ],
   alphaCSR[ 148 ][ 43 ],
   alphaCSR[ 148 ][ 44 ],
   alphaCSR[ 148 ][ 45 ],
   alphaCSR[ 148 ][ 46 ],
   alphaCSR[ 148 ][ 47 ],
   alphaCSR[ 148 ][ 48 ],
   alphaCSR[ 148 ][ 49 ],
   alphaCSR[ 148 ][ 50 ],
   alphaCSR[ 148 ][ 51 ],
   alphaCSR[ 148 ][ 52 ],
   alphaCSR[ 148 ][ 53 ],
   alphaCSR[ 148 ][ 54 ],
   alphaCSR[ 148 ][ 55 ],
   alphaCSR[ 148 ][ 56 ],
   alphaCSR[ 148 ][ 57 ],
   alphaCSR[ 148 ][ 58 ],
   alphaCSR[ 148 ][ 59 ],
   alphaCSR[ 148 ][ 60 ],
   alphaCSR[ 148 ][ 61 ],
   alphaCSR[ 148 ][ 62 ],
   alphaCSR[ 148 ][ 63 ],
   alphaCSR[ 148 ][ 64 ],
   alphaCSR[ 148 ][ 65 ],
   alphaCSR[ 148 ][ 66 ],
   alphaCSR[ 148 ][ 67 ],
   alphaCSR[ 148 ][ 68 ],
   alphaCSR[ 148 ][ 69 ],
   alphaCSR[ 148 ][ 70 ],
   alphaCSR[ 148 ][ 71 ],
   alphaCSR[ 148 ][ 72 ],
   alphaCSR[ 148 ][ 73 ],
   alphaCSR[ 148 ][ 74 ],
   alphaCSR[ 148 ][ 75 ],
   alphaCSR[ 148 ][ 76 ],
   alphaCSR[ 148 ][ 77 ],
   alphaCSR[ 148 ][ 78 ],
   alphaCSR[ 148 ][ 79 ],
   alphaCSR[ 148 ][ 80 ],
   alphaCSR[ 148 ][ 81 ],
   alphaCSR[ 148 ][ 82 ],
   alphaCSR[ 148 ][ 83 ],
   alphaCSR[ 148 ][ 84 ],
   alphaCSR[ 148 ][ 85 ],
   alphaCSR[ 148 ][ 86 ],
   alphaCSR[ 148 ][ 87 ],
   alphaCSR[ 148 ][ 88 ],
   alphaCSR[ 148 ][ 89 ],
   alphaCSR[ 148 ][ 90 ],
   alphaCSR[ 148 ][ 91 ],
   alphaCSR[ 148 ][ 92 ],
   alphaCSR[ 148 ][ 93 ],
   alphaCSR[ 148 ][ 94 ],
   alphaCSR[ 148 ][ 95 ],
   alphaCSR[ 148 ][ 96 ],
   alphaCSR[ 148 ][ 97 ],
   alphaCSR[ 148 ][ 98 ],
   alphaCSR[ 148 ][ 99 ],
   alphaCSR[ 148 ][ 100 ],
   alphaCSR[ 148 ][ 101 ],
   alphaCSR[ 148 ][ 102 ],
   alphaCSR[ 148 ][ 103 ],
   alphaCSR[ 148 ][ 104 ],
   alphaCSR[ 148 ][ 105 ],
   alphaCSR[ 148 ][ 106 ],
   alphaCSR[ 148 ][ 107 ],
   alphaCSR[ 148 ][ 108 ],
   alphaCSR[ 148 ][ 109 ],
   alphaCSR[ 148 ][ 110 ],
   alphaCSR[ 148 ][ 111 ],
   alphaCSR[ 148 ][ 112 ],
   alphaCSR[ 148 ][ 113 ],
   alphaCSR[ 148 ][ 114 ],
   alphaCSR[ 148 ][ 115 ],
   alphaCSR[ 148 ][ 116 ],
   alphaCSR[ 148 ][ 117 ],
   alphaCSR[ 148 ][ 118 ],
   alphaCSR[ 148 ][ 119 ],
   alphaCSR[ 148 ][ 120 ],
   alphaCSR[ 148 ][ 121 ],
   alphaCSR[ 148 ][ 122 ],
   alphaCSR[ 148 ][ 123 ],
   alphaCSR[ 148 ][ 124 ],
   alphaCSR[ 148 ][ 125 ],
   alphaCSR[ 148 ][ 126 ],
   alphaCSR[ 148 ][ 127 ],
   alphaCSR[ 148 ][ 128 ],
   alphaCSR[ 148 ][ 129 ],
   alphaCSR[ 148 ][ 130 ],
   alphaCSR[ 148 ][ 131 ],
   alphaCSR[ 148 ][ 132 ],
   alphaCSR[ 148 ][ 133 ],
   alphaCSR[ 148 ][ 134 ],
   alphaCSR[ 148 ][ 135 ],
   alphaCSR[ 148 ][ 136 ],
   alphaCSR[ 148 ][ 137 ],
   alphaCSR[ 148 ][ 138 ],
   alphaCSR[ 148 ][ 139 ],
   alphaCSR[ 148 ][ 140 ],
   alphaCSR[ 148 ][ 141 ],
   alphaCSR[ 148 ][ 142 ],
   alphaCSR[ 148 ][ 143 ],
   alphaCSR[ 148 ][ 144 ],
   alphaCSR[ 148 ][ 145 ],
   alphaCSR[ 148 ][ 146 ],
   alphaCSR[ 148 ][ 147 ],
   alphaCSR[ 148 ][ 148 ],
   alphaCSR[ 148 ][ 149 ],
   alphaCSR[ 148 ][ 150 ],
   alphaCSR[ 148 ][ 151 ],
   alphaCSR[ 148 ][ 152 ],
   alphaCSR[ 148 ][ 153 ],
   alphaCSR[ 148 ][ 154 ],
   alphaCSR[ 148 ][ 155 ],
   alphaCSR[ 148 ][ 156 ],
   alphaCSR[ 148 ][ 157 ],
   alphaCSR[ 148 ][ 158 ],
   alphaCSR[ 148 ][ 159 ],
   alphaCSR[ 148 ][ 160 ],
   alphaCSR[ 148 ][ 161 ],
   alphaCSR[ 148 ][ 162 ],
   alphaCSR[ 148 ][ 163 ],
   alphaCSR[ 148 ][ 164 ],
   alphaCSR[ 148 ][ 165 ],
   alphaCSR[ 148 ][ 166 ],
   alphaCSR[ 148 ][ 167 ],
   alphaCSR[ 148 ][ 168 ],
   alphaCSR[ 148 ][ 169 ],
   alphaCSR[ 148 ][ 170 ],
   alphaCSR[ 148 ][ 171 ],
   alphaCSR[ 148 ][ 172 ],
   alphaCSR[ 148 ][ 173 ],
   alphaCSR[ 148 ][ 174 ],
   alphaCSR[ 148 ][ 175 ],
   alphaCSR[ 148 ][ 176 ],
   alphaCSR[ 148 ][ 177 ],
   alphaCSR[ 148 ][ 178 ],
   alphaCSR[ 148 ][ 179 ],
   alphaCSR[ 148 ][ 180 ],
   alphaCSR[ 148 ][ 181 ],
   alphaCSR[ 148 ][ 182 ],
   alphaCSR[ 148 ][ 183 ],
   alphaCSR[ 148 ][ 184 ],
   alphaCSR[ 148 ][ 185 ],
   alphaCSR[ 148 ][ 186 ],
   alphaCSR[ 148 ][ 187 ],
   alphaCSR[ 148 ][ 188 ],
   alphaCSR[ 148 ][ 189 ],
   alphaCSR[ 148 ][ 190 ],
   alphaCSR[ 148 ][ 191 ],
   alphaCSR[ 148 ][ 192 ],
   alphaCSR[ 148 ][ 193 ],
   alphaCSR[ 148 ][ 194 ],
   alphaCSR[ 148 ][ 195 ],
   alphaCSR[ 148 ][ 196 ],
   alphaCSR[ 148 ][ 197 ],
   alphaCSR[ 148 ][ 198 ],
   alphaCSR[ 148 ][ 199 ],
   alphaCSR[ 148 ][ 200 ],
   alphaCSR[ 148 ][ 201 ],
   alphaCSR[ 148 ][ 202 ],
   alphaCSR[ 148 ][ 203 ],
   alphaCSR[ 148 ][ 204 ],
   alphaCSR[ 148 ][ 205 ],
   alphaCSR[ 148 ][ 206 ],
   alphaCSR[ 148 ][ 207 ],
   alphaCSR[ 148 ][ 208 ],
   alphaCSR[ 148 ][ 209 ],
   alphaCSR[ 148 ][ 210 ],
   alphaCSR[ 148 ][ 211 ],
   alphaCSR[ 148 ][ 212 ],
   alphaCSR[ 148 ][ 213 ],
   alphaCSR[ 148 ][ 214 ],
   alphaCSR[ 148 ][ 215 ],
   alphaCSR[ 148 ][ 216 ],
   alphaCSR[ 148 ][ 217 ],
   alphaCSR[ 148 ][ 218 ],
   alphaCSR[ 148 ][ 219 ],
   alphaCSR[ 148 ][ 220 ],
   alphaCSR[ 148 ][ 221 ],
   alphaCSR[ 148 ][ 222 ],
   alphaCSR[ 148 ][ 223 ],
   alphaCSR[ 148 ][ 224 ],
   alphaCSR[ 148 ][ 225 ],
   alphaCSR[ 148 ][ 226 ],
   alphaCSR[ 148 ][ 227 ],
   alphaCSR[ 148 ][ 228 ],
   alphaCSR[ 148 ][ 229 ],
   alphaCSR[ 148 ][ 230 ],
   alphaCSR[ 148 ][ 231 ],
   alphaCSR[ 148 ][ 232 ],
   alphaCSR[ 148 ][ 233 ],
   alphaCSR[ 148 ][ 234 ],
   alphaCSR[ 148 ][ 235 ],
   alphaCSR[ 148 ][ 236 ],
   alphaCSR[ 148 ][ 237 ],
   alphaCSR[ 148 ][ 238 ],
   alphaCSR[ 148 ][ 239 ],
   alphaCSR[ 148 ][ 240 ],
   alphaCSR[ 148 ][ 241 ],
   alphaCSR[ 148 ][ 242 ],
   alphaCSR[ 148 ][ 243 ],
   alphaCSR[ 148 ][ 244 ],
   alphaCSR[ 148 ][ 245 ],
   alphaCSR[ 148 ][ 246 ],
   alphaCSR[ 148 ][ 247 ],
   alphaCSR[ 148 ][ 248 ],
   alphaCSR[ 148 ][ 249 ],
   alphaCSR[ 148 ][ 250 ],
   alphaCSR[ 148 ][ 251 ],
   alphaCSR[ 148 ][ 252 ],
   alphaCSR[ 148 ][ 253 ],
   alphaCSR[ 148 ][ 254 ],
   alphaCSR[ 148 ][ 255 ],
   alphaCSR[ 148 ][ 256 ],
   alphaCSR[ 148 ][ 257 ],
   alphaCSR[ 148 ][ 258 ],
   alphaCSR[ 148 ][ 259 ],
   alphaCSR[ 148 ][ 260 ],
   alphaCSR[ 148 ][ 261 ],
   alphaCSR[ 148 ][ 262 ],
   alphaCSR[ 148 ][ 263 ],
   alphaCSR[ 148 ][ 264 ],
   alphaCSR[ 148 ][ 265 ],
   alphaCSR[ 148 ][ 266 ],
   alphaCSR[ 148 ][ 267 ],
   alphaCSR[ 148 ][ 268 ],
   alphaCSR[ 148 ][ 269 ],
   alphaCSR[ 148 ][ 270 ],
   alphaCSR[ 148 ][ 271 ],
   alphaCSR[ 148 ][ 272 ],
   alphaCSR[ 148 ][ 273 ],
   alphaCSR[ 148 ][ 274 ],
   alphaCSR[ 148 ][ 275 ],
   alphaCSR[ 148 ][ 276 ],
   alphaCSR[ 148 ][ 277 ],
   alphaCSR[ 148 ][ 278 ],
   alphaCSR[ 148 ][ 279 ],
   alphaCSR[ 148 ][ 280 ],
   alphaCSR[ 148 ][ 281 ],
   alphaCSR[ 148 ][ 282 ],
   alphaCSR[ 148 ][ 283 ],
   alphaCSR[ 148 ][ 284 ],
   alphaCSR[ 148 ][ 285 ],
   alphaCSR[ 148 ][ 286 ],
   alphaCSR[ 148 ][ 287 ],
   alphaCSR[ 148 ][ 288 ],
   alphaCSR[ 148 ][ 289 ],
   alphaCSR[ 148 ][ 290 ],
   alphaCSR[ 148 ][ 291 ],
   alphaCSR[ 148 ][ 292 ],
   alphaCSR[ 148 ][ 293 ],
   alphaCSR[ 148 ][ 294 ],
   alphaCSR[ 148 ][ 295 ],
   alphaCSR[ 148 ][ 296 ],
   alphaCSR[ 148 ][ 297 ],
   alphaCSR[ 148 ][ 298 ],
   alphaCSR[ 148 ][ 299 ],
   alphaCSR[ 148 ][ 300 ],
   alphaCSR[ 148 ][ 301 ],
   alphaCSR[ 148 ][ 302 ],
   alphaCSR[ 148 ][ 303 ],
   alphaCSR[ 148 ][ 304 ],
   alphaCSR[ 148 ][ 305 ],
   alphaCSR[ 148 ][ 306 ],
   alphaCSR[ 148 ][ 307 ],
   alphaCSR[ 148 ][ 308 ],
   alphaCSR[ 148 ][ 309 ],
   alphaCSR[ 148 ][ 310 ],
   alphaCSR[ 148 ][ 311 ],
   alphaCSR[ 148 ][ 312 ],
   alphaCSR[ 148 ][ 313 ],
   alphaCSR[ 148 ][ 314 ],
   alphaCSR[ 148 ][ 315 ],
   alphaCSR[ 148 ][ 316 ],
   alphaCSR[ 148 ][ 317 ],
   alphaCSR[ 148 ][ 318 ],
   alphaCSR[ 148 ][ 319 ],
   alphaCSR[ 148 ][ 320 ],
   alphaCSR[ 148 ][ 321 ],
   alphaCSR[ 148 ][ 322 ],
   alphaCSR[ 148 ][ 323 ],
   alphaCSR[ 148 ][ 324 ],
   alphaCSR[ 148 ][ 325 ],
   alphaCSR[ 148 ][ 326 ],
   alphaCSR[ 148 ][ 327 ],
   alphaCSR[ 148 ][ 328 ],
   alphaCSR[ 148 ][ 329 ],
   alphaCSR[ 148 ][ 330 ],
   alphaCSR[ 148 ][ 331 ],
   alphaCSR[ 148 ][ 332 ],
   alphaCSR[ 148 ][ 333 ],
   alphaCSR[ 148 ][ 334 ],
   alphaCSR[ 148 ][ 335 ],
   alphaCSR[ 148 ][ 336 ],
   alphaCSR[ 148 ][ 337 ],
   alphaCSR[ 148 ][ 338 ],
   alphaCSR[ 148 ][ 339 ],
   alphaCSR[ 148 ][ 340 ],
   alphaCSR[ 148 ][ 341 ],
   alphaCSR[ 148 ][ 342 ],
   alphaCSR[ 148 ][ 343 ],
   alphaCSR[ 148 ][ 344 ],
   alphaCSR[ 148 ][ 345 ],
   alphaCSR[ 148 ][ 346 ],
   alphaCSR[ 148 ][ 347 ],
   alphaCSR[ 148 ][ 348 ],
   alphaCSR[ 148 ][ 349 ],
   alphaCSR[ 148 ][ 350 ],
   alphaCSR[ 148 ][ 351 ],
   alphaCSR[ 148 ][ 352 ],
   alphaCSR[ 148 ][ 353 ],
   alphaCSR[ 148 ][ 354 ],
   alphaCSR[ 148 ][ 355 ],
   alphaCSR[ 148 ][ 356 ],
   alphaCSR[ 148 ][ 357 ],
   alphaCSR[ 148 ][ 358 ],
   alphaCSR[ 148 ][ 359 ],
   alphaCSR[ 148 ][ 360 ],
   alphaCSR[ 148 ][ 361 ],
   alphaCSR[ 148 ][ 362 ],
   alphaCSR[ 148 ][ 363 ],
   alphaCSR[ 148 ][ 364 ],
   alphaCSR[ 148 ][ 365 ],
   alphaCSR[ 148 ][ 366 ],
   alphaCSR[ 148 ][ 367 ],
   alphaCSR[ 148 ][ 368 ],
   alphaCSR[ 148 ][ 369 ],
   alphaCSR[ 148 ][ 370 ],
   alphaCSR[ 148 ][ 371 ],
   alphaCSR[ 148 ][ 372 ],
   alphaCSR[ 148 ][ 373 ],
   alphaCSR[ 148 ][ 374 ],
   alphaCSR[ 148 ][ 375 ],
   alphaCSR[ 148 ][ 376 ],
   alphaCSR[ 148 ][ 377 ],
   alphaCSR[ 148 ][ 378 ],
   alphaCSR[ 148 ][ 379 ],
   alphaCSR[ 148 ][ 380 ],
   alphaCSR[ 148 ][ 381 ],
   alphaCSR[ 148 ][ 382 ],
   alphaCSR[ 148 ][ 383 ],
   alphaCSR[ 149 ][ 0 ],
   alphaCSR[ 149 ][ 1 ],
   alphaCSR[ 149 ][ 2 ],
   alphaCSR[ 149 ][ 3 ],
   alphaCSR[ 149 ][ 4 ],
   alphaCSR[ 149 ][ 5 ],
   alphaCSR[ 149 ][ 6 ],
   alphaCSR[ 149 ][ 7 ],
   alphaCSR[ 149 ][ 8 ],
   alphaCSR[ 149 ][ 9 ],
   alphaCSR[ 149 ][ 10 ],
   alphaCSR[ 149 ][ 11 ],
   alphaCSR[ 149 ][ 12 ],
   alphaCSR[ 149 ][ 13 ],
   alphaCSR[ 149 ][ 14 ],
   alphaCSR[ 149 ][ 15 ],
   alphaCSR[ 149 ][ 16 ],
   alphaCSR[ 149 ][ 17 ],
   alphaCSR[ 149 ][ 18 ],
   alphaCSR[ 149 ][ 19 ],
   alphaCSR[ 149 ][ 20 ],
   alphaCSR[ 149 ][ 21 ],
   alphaCSR[ 149 ][ 22 ],
   alphaCSR[ 149 ][ 23 ],
   alphaCSR[ 149 ][ 24 ],
   alphaCSR[ 149 ][ 25 ],
   alphaCSR[ 149 ][ 26 ],
   alphaCSR[ 149 ][ 27 ],
   alphaCSR[ 149 ][ 28 ],
   alphaCSR[ 149 ][ 29 ],
   alphaCSR[ 149 ][ 30 ],
   alphaCSR[ 149 ][ 31 ],
   alphaCSR[ 149 ][ 32 ],
   alphaCSR[ 149 ][ 33 ],
   alphaCSR[ 149 ][ 34 ],
   alphaCSR[ 149 ][ 35 ],
   alphaCSR[ 149 ][ 36 ],
   alphaCSR[ 149 ][ 37 ],
   alphaCSR[ 149 ][ 38 ],
   alphaCSR[ 149 ][ 39 ],
   alphaCSR[ 149 ][ 40 ],
   alphaCSR[ 149 ][ 41 ],
   alphaCSR[ 149 ][ 42 ],
   alphaCSR[ 149 ][ 43 ],
   alphaCSR[ 149 ][ 44 ],
   alphaCSR[ 149 ][ 45 ],
   alphaCSR[ 149 ][ 46 ],
   alphaCSR[ 149 ][ 47 ],
   alphaCSR[ 149 ][ 48 ],
   alphaCSR[ 149 ][ 49 ],
   alphaCSR[ 149 ][ 50 ],
   alphaCSR[ 149 ][ 51 ],
   alphaCSR[ 149 ][ 52 ],
   alphaCSR[ 149 ][ 53 ],
   alphaCSR[ 149 ][ 54 ],
   alphaCSR[ 149 ][ 55 ],
   alphaCSR[ 149 ][ 56 ],
   alphaCSR[ 149 ][ 57 ],
   alphaCSR[ 149 ][ 58 ],
   alphaCSR[ 149 ][ 59 ],
   alphaCSR[ 149 ][ 60 ],
   alphaCSR[ 149 ][ 61 ],
   alphaCSR[ 149 ][ 62 ],
   alphaCSR[ 149 ][ 63 ],
   alphaCSR[ 149 ][ 64 ],
   alphaCSR[ 149 ][ 65 ],
   alphaCSR[ 149 ][ 66 ],
   alphaCSR[ 149 ][ 67 ],
   alphaCSR[ 149 ][ 68 ],
   alphaCSR[ 149 ][ 69 ],
   alphaCSR[ 149 ][ 70 ],
   alphaCSR[ 149 ][ 71 ],
   alphaCSR[ 149 ][ 72 ],
   alphaCSR[ 149 ][ 73 ],
   alphaCSR[ 149 ][ 74 ],
   alphaCSR[ 149 ][ 75 ],
   alphaCSR[ 149 ][ 76 ],
   alphaCSR[ 149 ][ 77 ],
   alphaCSR[ 149 ][ 78 ],
   alphaCSR[ 149 ][ 79 ],
   alphaCSR[ 149 ][ 80 ],
   alphaCSR[ 149 ][ 81 ],
   alphaCSR[ 149 ][ 82 ],
   alphaCSR[ 149 ][ 83 ],
   alphaCSR[ 149 ][ 84 ],
   alphaCSR[ 149 ][ 85 ],
   alphaCSR[ 149 ][ 86 ],
   alphaCSR[ 149 ][ 87 ],
   alphaCSR[ 149 ][ 88 ],
   alphaCSR[ 149 ][ 89 ],
   alphaCSR[ 149 ][ 90 ],
   alphaCSR[ 149 ][ 91 ],
   alphaCSR[ 149 ][ 92 ],
   alphaCSR[ 149 ][ 93 ],
   alphaCSR[ 149 ][ 94 ],
   alphaCSR[ 149 ][ 95 ],
   alphaCSR[ 149 ][ 96 ],
   alphaCSR[ 149 ][ 97 ],
   alphaCSR[ 149 ][ 98 ],
   alphaCSR[ 149 ][ 99 ],
   alphaCSR[ 149 ][ 100 ],
   alphaCSR[ 149 ][ 101 ],
   alphaCSR[ 149 ][ 102 ],
   alphaCSR[ 149 ][ 103 ],
   alphaCSR[ 149 ][ 104 ],
   alphaCSR[ 149 ][ 105 ],
   alphaCSR[ 149 ][ 106 ],
   alphaCSR[ 149 ][ 107 ],
   alphaCSR[ 149 ][ 108 ],
   alphaCSR[ 149 ][ 109 ],
   alphaCSR[ 149 ][ 110 ],
   alphaCSR[ 149 ][ 111 ],
   alphaCSR[ 149 ][ 112 ],
   alphaCSR[ 149 ][ 113 ],
   alphaCSR[ 149 ][ 114 ],
   alphaCSR[ 149 ][ 115 ],
   alphaCSR[ 149 ][ 116 ],
   alphaCSR[ 149 ][ 117 ],
   alphaCSR[ 149 ][ 118 ],
   alphaCSR[ 149 ][ 119 ],
   alphaCSR[ 149 ][ 120 ],
   alphaCSR[ 149 ][ 121 ],
   alphaCSR[ 149 ][ 122 ],
   alphaCSR[ 149 ][ 123 ],
   alphaCSR[ 149 ][ 124 ],
   alphaCSR[ 149 ][ 125 ],
   alphaCSR[ 149 ][ 126 ],
   alphaCSR[ 149 ][ 127 ],
   alphaCSR[ 149 ][ 128 ],
   alphaCSR[ 149 ][ 129 ],
   alphaCSR[ 149 ][ 130 ],
   alphaCSR[ 149 ][ 131 ],
   alphaCSR[ 149 ][ 132 ],
   alphaCSR[ 149 ][ 133 ],
   alphaCSR[ 149 ][ 134 ],
   alphaCSR[ 149 ][ 135 ],
   alphaCSR[ 149 ][ 136 ],
   alphaCSR[ 149 ][ 137 ],
   alphaCSR[ 149 ][ 138 ],
   alphaCSR[ 149 ][ 139 ],
   alphaCSR[ 149 ][ 140 ],
   alphaCSR[ 149 ][ 141 ],
   alphaCSR[ 149 ][ 142 ],
   alphaCSR[ 149 ][ 143 ],
   alphaCSR[ 149 ][ 144 ],
   alphaCSR[ 149 ][ 145 ],
   alphaCSR[ 149 ][ 146 ],
   alphaCSR[ 149 ][ 147 ],
   alphaCSR[ 149 ][ 148 ],
   alphaCSR[ 149 ][ 149 ],
   alphaCSR[ 149 ][ 150 ],
   alphaCSR[ 149 ][ 151 ],
   alphaCSR[ 149 ][ 152 ],
   alphaCSR[ 149 ][ 153 ],
   alphaCSR[ 149 ][ 154 ],
   alphaCSR[ 149 ][ 155 ],
   alphaCSR[ 149 ][ 156 ],
   alphaCSR[ 149 ][ 157 ],
   alphaCSR[ 149 ][ 158 ],
   alphaCSR[ 149 ][ 159 ],
   alphaCSR[ 149 ][ 160 ],
   alphaCSR[ 149 ][ 161 ],
   alphaCSR[ 149 ][ 162 ],
   alphaCSR[ 149 ][ 163 ],
   alphaCSR[ 149 ][ 164 ],
   alphaCSR[ 149 ][ 165 ],
   alphaCSR[ 149 ][ 166 ],
   alphaCSR[ 149 ][ 167 ],
   alphaCSR[ 149 ][ 168 ],
   alphaCSR[ 149 ][ 169 ],
   alphaCSR[ 149 ][ 170 ],
   alphaCSR[ 149 ][ 171 ],
   alphaCSR[ 149 ][ 172 ],
   alphaCSR[ 149 ][ 173 ],
   alphaCSR[ 149 ][ 174 ],
   alphaCSR[ 149 ][ 175 ],
   alphaCSR[ 149 ][ 176 ],
   alphaCSR[ 149 ][ 177 ],
   alphaCSR[ 149 ][ 178 ],
   alphaCSR[ 149 ][ 179 ],
   alphaCSR[ 149 ][ 180 ],
   alphaCSR[ 149 ][ 181 ],
   alphaCSR[ 149 ][ 182 ],
   alphaCSR[ 149 ][ 183 ],
   alphaCSR[ 149 ][ 184 ],
   alphaCSR[ 149 ][ 185 ],
   alphaCSR[ 149 ][ 186 ],
   alphaCSR[ 149 ][ 187 ],
   alphaCSR[ 149 ][ 188 ],
   alphaCSR[ 149 ][ 189 ],
   alphaCSR[ 149 ][ 190 ],
   alphaCSR[ 149 ][ 191 ],
   alphaCSR[ 149 ][ 192 ],
   alphaCSR[ 149 ][ 193 ],
   alphaCSR[ 149 ][ 194 ],
   alphaCSR[ 149 ][ 195 ],
   alphaCSR[ 149 ][ 196 ],
   alphaCSR[ 149 ][ 197 ],
   alphaCSR[ 149 ][ 198 ],
   alphaCSR[ 149 ][ 199 ],
   alphaCSR[ 149 ][ 200 ],
   alphaCSR[ 149 ][ 201 ],
   alphaCSR[ 149 ][ 202 ],
   alphaCSR[ 149 ][ 203 ],
   alphaCSR[ 149 ][ 204 ],
   alphaCSR[ 149 ][ 205 ],
   alphaCSR[ 149 ][ 206 ],
   alphaCSR[ 149 ][ 207 ],
   alphaCSR[ 149 ][ 208 ],
   alphaCSR[ 149 ][ 209 ],
   alphaCSR[ 149 ][ 210 ],
   alphaCSR[ 149 ][ 211 ],
   alphaCSR[ 149 ][ 212 ],
   alphaCSR[ 149 ][ 213 ],
   alphaCSR[ 149 ][ 214 ],
   alphaCSR[ 149 ][ 215 ],
   alphaCSR[ 149 ][ 216 ],
   alphaCSR[ 149 ][ 217 ],
   alphaCSR[ 149 ][ 218 ],
   alphaCSR[ 149 ][ 219 ],
   alphaCSR[ 149 ][ 220 ],
   alphaCSR[ 149 ][ 221 ],
   alphaCSR[ 149 ][ 222 ],
   alphaCSR[ 149 ][ 223 ],
   alphaCSR[ 149 ][ 224 ],
   alphaCSR[ 149 ][ 225 ],
   alphaCSR[ 149 ][ 226 ],
   alphaCSR[ 149 ][ 227 ],
   alphaCSR[ 149 ][ 228 ],
   alphaCSR[ 149 ][ 229 ],
   alphaCSR[ 149 ][ 230 ],
   alphaCSR[ 149 ][ 231 ],
   alphaCSR[ 149 ][ 232 ],
   alphaCSR[ 149 ][ 233 ],
   alphaCSR[ 149 ][ 234 ],
   alphaCSR[ 149 ][ 235 ],
   alphaCSR[ 149 ][ 236 ],
   alphaCSR[ 149 ][ 237 ],
   alphaCSR[ 149 ][ 238 ],
   alphaCSR[ 149 ][ 239 ],
   alphaCSR[ 149 ][ 240 ],
   alphaCSR[ 149 ][ 241 ],
   alphaCSR[ 149 ][ 242 ],
   alphaCSR[ 149 ][ 243 ],
   alphaCSR[ 149 ][ 244 ],
   alphaCSR[ 149 ][ 245 ],
   alphaCSR[ 149 ][ 246 ],
   alphaCSR[ 149 ][ 247 ],
   alphaCSR[ 149 ][ 248 ],
   alphaCSR[ 149 ][ 249 ],
   alphaCSR[ 149 ][ 250 ],
   alphaCSR[ 149 ][ 251 ],
   alphaCSR[ 149 ][ 252 ],
   alphaCSR[ 149 ][ 253 ],
   alphaCSR[ 149 ][ 254 ],
   alphaCSR[ 149 ][ 255 ],
   alphaCSR[ 149 ][ 256 ],
   alphaCSR[ 149 ][ 257 ],
   alphaCSR[ 149 ][ 258 ],
   alphaCSR[ 149 ][ 259 ],
   alphaCSR[ 149 ][ 260 ],
   alphaCSR[ 149 ][ 261 ],
   alphaCSR[ 149 ][ 262 ],
   alphaCSR[ 149 ][ 263 ],
   alphaCSR[ 149 ][ 264 ],
   alphaCSR[ 149 ][ 265 ],
   alphaCSR[ 149 ][ 266 ],
   alphaCSR[ 149 ][ 267 ],
   alphaCSR[ 149 ][ 268 ],
   alphaCSR[ 149 ][ 269 ],
   alphaCSR[ 149 ][ 270 ],
   alphaCSR[ 149 ][ 271 ],
   alphaCSR[ 149 ][ 272 ],
   alphaCSR[ 149 ][ 273 ],
   alphaCSR[ 149 ][ 274 ],
   alphaCSR[ 149 ][ 275 ],
   alphaCSR[ 149 ][ 276 ],
   alphaCSR[ 149 ][ 277 ],
   alphaCSR[ 149 ][ 278 ],
   alphaCSR[ 149 ][ 279 ],
   alphaCSR[ 149 ][ 280 ],
   alphaCSR[ 149 ][ 281 ],
   alphaCSR[ 149 ][ 282 ],
   alphaCSR[ 149 ][ 283 ],
   alphaCSR[ 149 ][ 284 ],
   alphaCSR[ 149 ][ 285 ],
   alphaCSR[ 149 ][ 286 ],
   alphaCSR[ 149 ][ 287 ],
   alphaCSR[ 149 ][ 288 ],
   alphaCSR[ 149 ][ 289 ],
   alphaCSR[ 149 ][ 290 ],
   alphaCSR[ 149 ][ 291 ],
   alphaCSR[ 149 ][ 292 ],
   alphaCSR[ 149 ][ 293 ],
   alphaCSR[ 149 ][ 294 ],
   alphaCSR[ 149 ][ 295 ],
   alphaCSR[ 149 ][ 296 ],
   alphaCSR[ 149 ][ 297 ],
   alphaCSR[ 149 ][ 298 ],
   alphaCSR[ 149 ][ 299 ],
   alphaCSR[ 149 ][ 300 ],
   alphaCSR[ 149 ][ 301 ],
   alphaCSR[ 149 ][ 302 ],
   alphaCSR[ 149 ][ 303 ],
   alphaCSR[ 149 ][ 304 ],
   alphaCSR[ 149 ][ 305 ],
   alphaCSR[ 149 ][ 306 ],
   alphaCSR[ 149 ][ 307 ],
   alphaCSR[ 149 ][ 308 ],
   alphaCSR[ 149 ][ 309 ],
   alphaCSR[ 149 ][ 310 ],
   alphaCSR[ 149 ][ 311 ],
   alphaCSR[ 149 ][ 312 ],
   alphaCSR[ 149 ][ 313 ],
   alphaCSR[ 149 ][ 314 ],
   alphaCSR[ 149 ][ 315 ],
   alphaCSR[ 149 ][ 316 ],
   alphaCSR[ 149 ][ 317 ],
   alphaCSR[ 149 ][ 318 ],
   alphaCSR[ 149 ][ 319 ],
   alphaCSR[ 149 ][ 320 ],
   alphaCSR[ 149 ][ 321 ],
   alphaCSR[ 149 ][ 322 ],
   alphaCSR[ 149 ][ 323 ],
   alphaCSR[ 149 ][ 324 ],
   alphaCSR[ 149 ][ 325 ],
   alphaCSR[ 149 ][ 326 ],
   alphaCSR[ 149 ][ 327 ],
   alphaCSR[ 149 ][ 328 ],
   alphaCSR[ 149 ][ 329 ],
   alphaCSR[ 149 ][ 330 ],
   alphaCSR[ 149 ][ 331 ],
   alphaCSR[ 149 ][ 332 ],
   alphaCSR[ 149 ][ 333 ],
   alphaCSR[ 149 ][ 334 ],
   alphaCSR[ 149 ][ 335 ],
   alphaCSR[ 149 ][ 336 ],
   alphaCSR[ 149 ][ 337 ],
   alphaCSR[ 149 ][ 338 ],
   alphaCSR[ 149 ][ 339 ],
   alphaCSR[ 149 ][ 340 ],
   alphaCSR[ 149 ][ 341 ],
   alphaCSR[ 149 ][ 342 ],
   alphaCSR[ 149 ][ 343 ],
   alphaCSR[ 149 ][ 344 ],
   alphaCSR[ 149 ][ 345 ],
   alphaCSR[ 149 ][ 346 ],
   alphaCSR[ 149 ][ 347 ],
   alphaCSR[ 149 ][ 348 ],
   alphaCSR[ 149 ][ 349 ],
   alphaCSR[ 149 ][ 350 ],
   alphaCSR[ 149 ][ 351 ],
   alphaCSR[ 149 ][ 352 ],
   alphaCSR[ 149 ][ 353 ],
   alphaCSR[ 149 ][ 354 ],
   alphaCSR[ 149 ][ 355 ],
   alphaCSR[ 149 ][ 356 ],
   alphaCSR[ 149 ][ 357 ],
   alphaCSR[ 149 ][ 358 ],
   alphaCSR[ 149 ][ 359 ],
   alphaCSR[ 149 ][ 360 ],
   alphaCSR[ 149 ][ 361 ],
   alphaCSR[ 149 ][ 362 ],
   alphaCSR[ 149 ][ 363 ],
   alphaCSR[ 149 ][ 364 ],
   alphaCSR[ 149 ][ 365 ],
   alphaCSR[ 149 ][ 366 ],
   alphaCSR[ 149 ][ 367 ],
   alphaCSR[ 149 ][ 368 ],
   alphaCSR[ 149 ][ 369 ],
   alphaCSR[ 149 ][ 370 ],
   alphaCSR[ 149 ][ 371 ],
   alphaCSR[ 149 ][ 372 ],
   alphaCSR[ 149 ][ 373 ],
   alphaCSR[ 149 ][ 374 ],
   alphaCSR[ 149 ][ 375 ],
   alphaCSR[ 149 ][ 376 ],
   alphaCSR[ 149 ][ 377 ],
   alphaCSR[ 149 ][ 378 ],
   alphaCSR[ 149 ][ 379 ],
   alphaCSR[ 149 ][ 380 ],
   alphaCSR[ 149 ][ 381 ],
   alphaCSR[ 149 ][ 382 ],
   alphaCSR[ 149 ][ 383 ],
   alphaCSR[ 150 ][ 0 ],
   alphaCSR[ 150 ][ 1 ],
   alphaCSR[ 150 ][ 2 ],
   alphaCSR[ 150 ][ 3 ],
   alphaCSR[ 150 ][ 4 ],
   alphaCSR[ 150 ][ 5 ],
   alphaCSR[ 150 ][ 6 ],
   alphaCSR[ 150 ][ 7 ],
   alphaCSR[ 150 ][ 8 ],
   alphaCSR[ 150 ][ 9 ],
   alphaCSR[ 150 ][ 10 ],
   alphaCSR[ 150 ][ 11 ],
   alphaCSR[ 150 ][ 12 ],
   alphaCSR[ 150 ][ 13 ],
   alphaCSR[ 150 ][ 14 ],
   alphaCSR[ 150 ][ 15 ],
   alphaCSR[ 150 ][ 16 ],
   alphaCSR[ 150 ][ 17 ],
   alphaCSR[ 150 ][ 18 ],
   alphaCSR[ 150 ][ 19 ],
   alphaCSR[ 150 ][ 20 ],
   alphaCSR[ 150 ][ 21 ],
   alphaCSR[ 150 ][ 22 ],
   alphaCSR[ 150 ][ 23 ],
   alphaCSR[ 150 ][ 24 ],
   alphaCSR[ 150 ][ 25 ],
   alphaCSR[ 150 ][ 26 ],
   alphaCSR[ 150 ][ 27 ],
   alphaCSR[ 150 ][ 28 ],
   alphaCSR[ 150 ][ 29 ],
   alphaCSR[ 150 ][ 30 ],
   alphaCSR[ 150 ][ 31 ],
   alphaCSR[ 150 ][ 32 ],
   alphaCSR[ 150 ][ 33 ],
   alphaCSR[ 150 ][ 34 ],
   alphaCSR[ 150 ][ 35 ],
   alphaCSR[ 150 ][ 36 ],
   alphaCSR[ 150 ][ 37 ],
   alphaCSR[ 150 ][ 38 ],
   alphaCSR[ 150 ][ 39 ],
   alphaCSR[ 150 ][ 40 ],
   alphaCSR[ 150 ][ 41 ],
   alphaCSR[ 150 ][ 42 ],
   alphaCSR[ 150 ][ 43 ],
   alphaCSR[ 150 ][ 44 ],
   alphaCSR[ 150 ][ 45 ],
   alphaCSR[ 150 ][ 46 ],
   alphaCSR[ 150 ][ 47 ],
   alphaCSR[ 150 ][ 48 ],
   alphaCSR[ 150 ][ 49 ],
   alphaCSR[ 150 ][ 50 ],
   alphaCSR[ 150 ][ 51 ],
   alphaCSR[ 150 ][ 52 ],
   alphaCSR[ 150 ][ 53 ],
   alphaCSR[ 150 ][ 54 ],
   alphaCSR[ 150 ][ 55 ],
   alphaCSR[ 150 ][ 56 ],
   alphaCSR[ 150 ][ 57 ],
   alphaCSR[ 150 ][ 58 ],
   alphaCSR[ 150 ][ 59 ],
   alphaCSR[ 150 ][ 60 ],
   alphaCSR[ 150 ][ 61 ],
   alphaCSR[ 150 ][ 62 ],
   alphaCSR[ 150 ][ 63 ],
   alphaCSR[ 150 ][ 64 ],
   alphaCSR[ 150 ][ 65 ],
   alphaCSR[ 150 ][ 66 ],
   alphaCSR[ 150 ][ 67 ],
   alphaCSR[ 150 ][ 68 ],
   alphaCSR[ 150 ][ 69 ],
   alphaCSR[ 150 ][ 70 ],
   alphaCSR[ 150 ][ 71 ],
   alphaCSR[ 150 ][ 72 ],
   alphaCSR[ 150 ][ 73 ],
   alphaCSR[ 150 ][ 74 ],
   alphaCSR[ 150 ][ 75 ],
   alphaCSR[ 150 ][ 76 ],
   alphaCSR[ 150 ][ 77 ],
   alphaCSR[ 150 ][ 78 ],
   alphaCSR[ 150 ][ 79 ],
   alphaCSR[ 150 ][ 80 ],
   alphaCSR[ 150 ][ 81 ],
   alphaCSR[ 150 ][ 82 ],
   alphaCSR[ 150 ][ 83 ],
   alphaCSR[ 150 ][ 84 ],
   alphaCSR[ 150 ][ 85 ],
   alphaCSR[ 150 ][ 86 ],
   alphaCSR[ 150 ][ 87 ],
   alphaCSR[ 150 ][ 88 ],
   alphaCSR[ 150 ][ 89 ],
   alphaCSR[ 150 ][ 90 ],
   alphaCSR[ 150 ][ 91 ],
   alphaCSR[ 150 ][ 92 ],
   alphaCSR[ 150 ][ 93 ],
   alphaCSR[ 150 ][ 94 ],
   alphaCSR[ 150 ][ 95 ],
   alphaCSR[ 150 ][ 96 ],
   alphaCSR[ 150 ][ 97 ],
   alphaCSR[ 150 ][ 98 ],
   alphaCSR[ 150 ][ 99 ],
   alphaCSR[ 150 ][ 100 ],
   alphaCSR[ 150 ][ 101 ],
   alphaCSR[ 150 ][ 102 ],
   alphaCSR[ 150 ][ 103 ],
   alphaCSR[ 150 ][ 104 ],
   alphaCSR[ 150 ][ 105 ],
   alphaCSR[ 150 ][ 106 ],
   alphaCSR[ 150 ][ 107 ],
   alphaCSR[ 150 ][ 108 ],
   alphaCSR[ 150 ][ 109 ],
   alphaCSR[ 150 ][ 110 ],
   alphaCSR[ 150 ][ 111 ],
   alphaCSR[ 150 ][ 112 ],
   alphaCSR[ 150 ][ 113 ],
   alphaCSR[ 150 ][ 114 ],
   alphaCSR[ 150 ][ 115 ],
   alphaCSR[ 150 ][ 116 ],
   alphaCSR[ 150 ][ 117 ],
   alphaCSR[ 150 ][ 118 ],
   alphaCSR[ 150 ][ 119 ],
   alphaCSR[ 150 ][ 120 ],
   alphaCSR[ 150 ][ 121 ],
   alphaCSR[ 150 ][ 122 ],
   alphaCSR[ 150 ][ 123 ],
   alphaCSR[ 150 ][ 124 ],
   alphaCSR[ 150 ][ 125 ],
   alphaCSR[ 150 ][ 126 ],
   alphaCSR[ 150 ][ 127 ],
   alphaCSR[ 150 ][ 128 ],
   alphaCSR[ 150 ][ 129 ],
   alphaCSR[ 150 ][ 130 ],
   alphaCSR[ 150 ][ 131 ],
   alphaCSR[ 150 ][ 132 ],
   alphaCSR[ 150 ][ 133 ],
   alphaCSR[ 150 ][ 134 ],
   alphaCSR[ 150 ][ 135 ],
   alphaCSR[ 150 ][ 136 ],
   alphaCSR[ 150 ][ 137 ],
   alphaCSR[ 150 ][ 138 ],
   alphaCSR[ 150 ][ 139 ],
   alphaCSR[ 150 ][ 140 ],
   alphaCSR[ 150 ][ 141 ],
   alphaCSR[ 150 ][ 142 ],
   alphaCSR[ 150 ][ 143 ],
   alphaCSR[ 150 ][ 144 ],
   alphaCSR[ 150 ][ 145 ],
   alphaCSR[ 150 ][ 146 ],
   alphaCSR[ 150 ][ 147 ],
   alphaCSR[ 150 ][ 148 ],
   alphaCSR[ 150 ][ 149 ],
   alphaCSR[ 150 ][ 150 ],
   alphaCSR[ 150 ][ 151 ],
   alphaCSR[ 150 ][ 152 ],
   alphaCSR[ 150 ][ 153 ],
   alphaCSR[ 150 ][ 154 ],
   alphaCSR[ 150 ][ 155 ],
   alphaCSR[ 150 ][ 156 ],
   alphaCSR[ 150 ][ 157 ],
   alphaCSR[ 150 ][ 158 ],
   alphaCSR[ 150 ][ 159 ],
   alphaCSR[ 150 ][ 160 ],
   alphaCSR[ 150 ][ 161 ],
   alphaCSR[ 150 ][ 162 ],
   alphaCSR[ 150 ][ 163 ],
   alphaCSR[ 150 ][ 164 ],
   alphaCSR[ 150 ][ 165 ],
   alphaCSR[ 150 ][ 166 ],
   alphaCSR[ 150 ][ 167 ],
   alphaCSR[ 150 ][ 168 ],
   alphaCSR[ 150 ][ 169 ],
   alphaCSR[ 150 ][ 170 ],
   alphaCSR[ 150 ][ 171 ],
   alphaCSR[ 150 ][ 172 ],
   alphaCSR[ 150 ][ 173 ],
   alphaCSR[ 150 ][ 174 ],
   alphaCSR[ 150 ][ 175 ],
   alphaCSR[ 150 ][ 176 ],
   alphaCSR[ 150 ][ 177 ],
   alphaCSR[ 150 ][ 178 ],
   alphaCSR[ 150 ][ 179 ],
   alphaCSR[ 150 ][ 180 ],
   alphaCSR[ 150 ][ 181 ],
   alphaCSR[ 150 ][ 182 ],
   alphaCSR[ 150 ][ 183 ],
   alphaCSR[ 150 ][ 184 ],
   alphaCSR[ 150 ][ 185 ],
   alphaCSR[ 150 ][ 186 ],
   alphaCSR[ 150 ][ 187 ],
   alphaCSR[ 150 ][ 188 ],
   alphaCSR[ 150 ][ 189 ],
   alphaCSR[ 150 ][ 190 ],
   alphaCSR[ 150 ][ 191 ],
   alphaCSR[ 150 ][ 192 ],
   alphaCSR[ 150 ][ 193 ],
   alphaCSR[ 150 ][ 194 ],
   alphaCSR[ 150 ][ 195 ],
   alphaCSR[ 150 ][ 196 ],
   alphaCSR[ 150 ][ 197 ],
   alphaCSR[ 150 ][ 198 ],
   alphaCSR[ 150 ][ 199 ],
   alphaCSR[ 150 ][ 200 ],
   alphaCSR[ 150 ][ 201 ],
   alphaCSR[ 150 ][ 202 ],
   alphaCSR[ 150 ][ 203 ],
   alphaCSR[ 150 ][ 204 ],
   alphaCSR[ 150 ][ 205 ],
   alphaCSR[ 150 ][ 206 ],
   alphaCSR[ 150 ][ 207 ],
   alphaCSR[ 150 ][ 208 ],
   alphaCSR[ 150 ][ 209 ],
   alphaCSR[ 150 ][ 210 ],
   alphaCSR[ 150 ][ 211 ],
   alphaCSR[ 150 ][ 212 ],
   alphaCSR[ 150 ][ 213 ],
   alphaCSR[ 150 ][ 214 ],
   alphaCSR[ 150 ][ 215 ],
   alphaCSR[ 150 ][ 216 ],
   alphaCSR[ 150 ][ 217 ],
   alphaCSR[ 150 ][ 218 ],
   alphaCSR[ 150 ][ 219 ],
   alphaCSR[ 150 ][ 220 ],
   alphaCSR[ 150 ][ 221 ],
   alphaCSR[ 150 ][ 222 ],
   alphaCSR[ 150 ][ 223 ],
   alphaCSR[ 150 ][ 224 ],
   alphaCSR[ 150 ][ 225 ],
   alphaCSR[ 150 ][ 226 ],
   alphaCSR[ 150 ][ 227 ],
   alphaCSR[ 150 ][ 228 ],
   alphaCSR[ 150 ][ 229 ],
   alphaCSR[ 150 ][ 230 ],
   alphaCSR[ 150 ][ 231 ],
   alphaCSR[ 150 ][ 232 ],
   alphaCSR[ 150 ][ 233 ],
   alphaCSR[ 150 ][ 234 ],
   alphaCSR[ 150 ][ 235 ],
   alphaCSR[ 150 ][ 236 ],
   alphaCSR[ 150 ][ 237 ],
   alphaCSR[ 150 ][ 238 ],
   alphaCSR[ 150 ][ 239 ],
   alphaCSR[ 150 ][ 240 ],
   alphaCSR[ 150 ][ 241 ],
   alphaCSR[ 150 ][ 242 ],
   alphaCSR[ 150 ][ 243 ],
   alphaCSR[ 150 ][ 244 ],
   alphaCSR[ 150 ][ 245 ],
   alphaCSR[ 150 ][ 246 ],
   alphaCSR[ 150 ][ 247 ],
   alphaCSR[ 150 ][ 248 ],
   alphaCSR[ 150 ][ 249 ],
   alphaCSR[ 150 ][ 250 ],
   alphaCSR[ 150 ][ 251 ],
   alphaCSR[ 150 ][ 252 ],
   alphaCSR[ 150 ][ 253 ],
   alphaCSR[ 150 ][ 254 ],
   alphaCSR[ 150 ][ 255 ],
   alphaCSR[ 150 ][ 256 ],
   alphaCSR[ 150 ][ 257 ],
   alphaCSR[ 150 ][ 258 ],
   alphaCSR[ 150 ][ 259 ],
   alphaCSR[ 150 ][ 260 ],
   alphaCSR[ 150 ][ 261 ],
   alphaCSR[ 150 ][ 262 ],
   alphaCSR[ 150 ][ 263 ],
   alphaCSR[ 150 ][ 264 ],
   alphaCSR[ 150 ][ 265 ],
   alphaCSR[ 150 ][ 266 ],
   alphaCSR[ 150 ][ 267 ],
   alphaCSR[ 150 ][ 268 ],
   alphaCSR[ 150 ][ 269 ],
   alphaCSR[ 150 ][ 270 ],
   alphaCSR[ 150 ][ 271 ],
   alphaCSR[ 150 ][ 272 ],
   alphaCSR[ 150 ][ 273 ],
   alphaCSR[ 150 ][ 274 ],
   alphaCSR[ 150 ][ 275 ],
   alphaCSR[ 150 ][ 276 ],
   alphaCSR[ 150 ][ 277 ],
   alphaCSR[ 150 ][ 278 ],
   alphaCSR[ 150 ][ 279 ],
   alphaCSR[ 150 ][ 280 ],
   alphaCSR[ 150 ][ 281 ],
   alphaCSR[ 150 ][ 282 ],
   alphaCSR[ 150 ][ 283 ],
   alphaCSR[ 150 ][ 284 ],
   alphaCSR[ 150 ][ 285 ],
   alphaCSR[ 150 ][ 286 ],
   alphaCSR[ 150 ][ 287 ],
   alphaCSR[ 150 ][ 288 ],
   alphaCSR[ 150 ][ 289 ],
   alphaCSR[ 150 ][ 290 ],
   alphaCSR[ 150 ][ 291 ],
   alphaCSR[ 150 ][ 292 ],
   alphaCSR[ 150 ][ 293 ],
   alphaCSR[ 150 ][ 294 ],
   alphaCSR[ 150 ][ 295 ],
   alphaCSR[ 150 ][ 296 ],
   alphaCSR[ 150 ][ 297 ],
   alphaCSR[ 150 ][ 298 ],
   alphaCSR[ 150 ][ 299 ],
   alphaCSR[ 150 ][ 300 ],
   alphaCSR[ 150 ][ 301 ],
   alphaCSR[ 150 ][ 302 ],
   alphaCSR[ 150 ][ 303 ],
   alphaCSR[ 150 ][ 304 ],
   alphaCSR[ 150 ][ 305 ],
   alphaCSR[ 150 ][ 306 ],
   alphaCSR[ 150 ][ 307 ],
   alphaCSR[ 150 ][ 308 ],
   alphaCSR[ 150 ][ 309 ],
   alphaCSR[ 150 ][ 310 ],
   alphaCSR[ 150 ][ 311 ],
   alphaCSR[ 150 ][ 312 ],
   alphaCSR[ 150 ][ 313 ],
   alphaCSR[ 150 ][ 314 ],
   alphaCSR[ 150 ][ 315 ],
   alphaCSR[ 150 ][ 316 ],
   alphaCSR[ 150 ][ 317 ],
   alphaCSR[ 150 ][ 318 ],
   alphaCSR[ 150 ][ 319 ],
   alphaCSR[ 150 ][ 320 ],
   alphaCSR[ 150 ][ 321 ],
   alphaCSR[ 150 ][ 322 ],
   alphaCSR[ 150 ][ 323 ],
   alphaCSR[ 150 ][ 324 ],
   alphaCSR[ 150 ][ 325 ],
   alphaCSR[ 150 ][ 326 ],
   alphaCSR[ 150 ][ 327 ],
   alphaCSR[ 150 ][ 328 ],
   alphaCSR[ 150 ][ 329 ],
   alphaCSR[ 150 ][ 330 ],
   alphaCSR[ 150 ][ 331 ],
   alphaCSR[ 150 ][ 332 ],
   alphaCSR[ 150 ][ 333 ],
   alphaCSR[ 150 ][ 334 ],
   alphaCSR[ 150 ][ 335 ],
   alphaCSR[ 150 ][ 336 ],
   alphaCSR[ 150 ][ 337 ],
   alphaCSR[ 150 ][ 338 ],
   alphaCSR[ 150 ][ 339 ],
   alphaCSR[ 150 ][ 340 ],
   alphaCSR[ 150 ][ 341 ],
   alphaCSR[ 150 ][ 342 ],
   alphaCSR[ 150 ][ 343 ],
   alphaCSR[ 150 ][ 344 ],
   alphaCSR[ 150 ][ 345 ],
   alphaCSR[ 150 ][ 346 ],
   alphaCSR[ 150 ][ 347 ],
   alphaCSR[ 150 ][ 348 ],
   alphaCSR[ 150 ][ 349 ],
   alphaCSR[ 150 ][ 350 ],
   alphaCSR[ 150 ][ 351 ],
   alphaCSR[ 150 ][ 352 ],
   alphaCSR[ 150 ][ 353 ],
   alphaCSR[ 150 ][ 354 ],
   alphaCSR[ 150 ][ 355 ],
   alphaCSR[ 150 ][ 356 ],
   alphaCSR[ 150 ][ 357 ],
   alphaCSR[ 150 ][ 358 ],
   alphaCSR[ 150 ][ 359 ],
   alphaCSR[ 150 ][ 360 ],
   alphaCSR[ 150 ][ 361 ],
   alphaCSR[ 150 ][ 362 ],
   alphaCSR[ 150 ][ 363 ],
   alphaCSR[ 150 ][ 364 ],
   alphaCSR[ 150 ][ 365 ],
   alphaCSR[ 150 ][ 366 ],
   alphaCSR[ 150 ][ 367 ],
   alphaCSR[ 150 ][ 368 ],
   alphaCSR[ 150 ][ 369 ],
   alphaCSR[ 150 ][ 370 ],
   alphaCSR[ 150 ][ 371 ],
   alphaCSR[ 150 ][ 372 ],
   alphaCSR[ 150 ][ 373 ],
   alphaCSR[ 150 ][ 374 ],
   alphaCSR[ 150 ][ 375 ],
   alphaCSR[ 150 ][ 376 ],
   alphaCSR[ 150 ][ 377 ],
   alphaCSR[ 150 ][ 378 ],
   alphaCSR[ 150 ][ 379 ],
   alphaCSR[ 150 ][ 380 ],
   alphaCSR[ 150 ][ 381 ],
   alphaCSR[ 150 ][ 382 ],
   alphaCSR[ 150 ][ 383 ],
   alphaCSR[ 151 ][ 0 ],
   alphaCSR[ 151 ][ 1 ],
   alphaCSR[ 151 ][ 2 ],
   alphaCSR[ 151 ][ 3 ],
   alphaCSR[ 151 ][ 4 ],
   alphaCSR[ 151 ][ 5 ],
   alphaCSR[ 151 ][ 6 ],
   alphaCSR[ 151 ][ 7 ],
   alphaCSR[ 151 ][ 8 ],
   alphaCSR[ 151 ][ 9 ],
   alphaCSR[ 151 ][ 10 ],
   alphaCSR[ 151 ][ 11 ],
   alphaCSR[ 151 ][ 12 ],
   alphaCSR[ 151 ][ 13 ],
   alphaCSR[ 151 ][ 14 ],
   alphaCSR[ 151 ][ 15 ],
   alphaCSR[ 151 ][ 16 ],
   alphaCSR[ 151 ][ 17 ],
   alphaCSR[ 151 ][ 18 ],
   alphaCSR[ 151 ][ 19 ],
   alphaCSR[ 151 ][ 20 ],
   alphaCSR[ 151 ][ 21 ],
   alphaCSR[ 151 ][ 22 ],
   alphaCSR[ 151 ][ 23 ],
   alphaCSR[ 151 ][ 24 ],
   alphaCSR[ 151 ][ 25 ],
   alphaCSR[ 151 ][ 26 ],
   alphaCSR[ 151 ][ 27 ],
   alphaCSR[ 151 ][ 28 ],
   alphaCSR[ 151 ][ 29 ],
   alphaCSR[ 151 ][ 30 ],
   alphaCSR[ 151 ][ 31 ],
   alphaCSR[ 151 ][ 32 ],
   alphaCSR[ 151 ][ 33 ],
   alphaCSR[ 151 ][ 34 ],
   alphaCSR[ 151 ][ 35 ],
   alphaCSR[ 151 ][ 36 ],
   alphaCSR[ 151 ][ 37 ],
   alphaCSR[ 151 ][ 38 ],
   alphaCSR[ 151 ][ 39 ],
   alphaCSR[ 151 ][ 40 ],
   alphaCSR[ 151 ][ 41 ],
   alphaCSR[ 151 ][ 42 ],
   alphaCSR[ 151 ][ 43 ],
   alphaCSR[ 151 ][ 44 ],
   alphaCSR[ 151 ][ 45 ],
   alphaCSR[ 151 ][ 46 ],
   alphaCSR[ 151 ][ 47 ],
   alphaCSR[ 151 ][ 48 ],
   alphaCSR[ 151 ][ 49 ],
   alphaCSR[ 151 ][ 50 ],
   alphaCSR[ 151 ][ 51 ],
   alphaCSR[ 151 ][ 52 ],
   alphaCSR[ 151 ][ 53 ],
   alphaCSR[ 151 ][ 54 ],
   alphaCSR[ 151 ][ 55 ],
   alphaCSR[ 151 ][ 56 ],
   alphaCSR[ 151 ][ 57 ],
   alphaCSR[ 151 ][ 58 ],
   alphaCSR[ 151 ][ 59 ],
   alphaCSR[ 151 ][ 60 ],
   alphaCSR[ 151 ][ 61 ],
   alphaCSR[ 151 ][ 62 ],
   alphaCSR[ 151 ][ 63 ],
   alphaCSR[ 151 ][ 64 ],
   alphaCSR[ 151 ][ 65 ],
   alphaCSR[ 151 ][ 66 ],
   alphaCSR[ 151 ][ 67 ],
   alphaCSR[ 151 ][ 68 ],
   alphaCSR[ 151 ][ 69 ],
   alphaCSR[ 151 ][ 70 ],
   alphaCSR[ 151 ][ 71 ],
   alphaCSR[ 151 ][ 72 ],
   alphaCSR[ 151 ][ 73 ],
   alphaCSR[ 151 ][ 74 ],
   alphaCSR[ 151 ][ 75 ],
   alphaCSR[ 151 ][ 76 ],
   alphaCSR[ 151 ][ 77 ],
   alphaCSR[ 151 ][ 78 ],
   alphaCSR[ 151 ][ 79 ],
   alphaCSR[ 151 ][ 80 ],
   alphaCSR[ 151 ][ 81 ],
   alphaCSR[ 151 ][ 82 ],
   alphaCSR[ 151 ][ 83 ],
   alphaCSR[ 151 ][ 84 ],
   alphaCSR[ 151 ][ 85 ],
   alphaCSR[ 151 ][ 86 ],
   alphaCSR[ 151 ][ 87 ],
   alphaCSR[ 151 ][ 88 ],
   alphaCSR[ 151 ][ 89 ],
   alphaCSR[ 151 ][ 90 ],
   alphaCSR[ 151 ][ 91 ],
   alphaCSR[ 151 ][ 92 ],
   alphaCSR[ 151 ][ 93 ],
   alphaCSR[ 151 ][ 94 ],
   alphaCSR[ 151 ][ 95 ],
   alphaCSR[ 151 ][ 96 ],
   alphaCSR[ 151 ][ 97 ],
   alphaCSR[ 151 ][ 98 ],
   alphaCSR[ 151 ][ 99 ],
   alphaCSR[ 151 ][ 100 ],
   alphaCSR[ 151 ][ 101 ],
   alphaCSR[ 151 ][ 102 ],
   alphaCSR[ 151 ][ 103 ],
   alphaCSR[ 151 ][ 104 ],
   alphaCSR[ 151 ][ 105 ],
   alphaCSR[ 151 ][ 106 ],
   alphaCSR[ 151 ][ 107 ],
   alphaCSR[ 151 ][ 108 ],
   alphaCSR[ 151 ][ 109 ],
   alphaCSR[ 151 ][ 110 ],
   alphaCSR[ 151 ][ 111 ],
   alphaCSR[ 151 ][ 112 ],
   alphaCSR[ 151 ][ 113 ],
   alphaCSR[ 151 ][ 114 ],
   alphaCSR[ 151 ][ 115 ],
   alphaCSR[ 151 ][ 116 ],
   alphaCSR[ 151 ][ 117 ],
   alphaCSR[ 151 ][ 118 ],
   alphaCSR[ 151 ][ 119 ],
   alphaCSR[ 151 ][ 120 ],
   alphaCSR[ 151 ][ 121 ],
   alphaCSR[ 151 ][ 122 ],
   alphaCSR[ 151 ][ 123 ],
   alphaCSR[ 151 ][ 124 ],
   alphaCSR[ 151 ][ 125 ],
   alphaCSR[ 151 ][ 126 ],
   alphaCSR[ 151 ][ 127 ],
   alphaCSR[ 151 ][ 128 ],
   alphaCSR[ 151 ][ 129 ],
   alphaCSR[ 151 ][ 130 ],
   alphaCSR[ 151 ][ 131 ],
   alphaCSR[ 151 ][ 132 ],
   alphaCSR[ 151 ][ 133 ],
   alphaCSR[ 151 ][ 134 ],
   alphaCSR[ 151 ][ 135 ],
   alphaCSR[ 151 ][ 136 ],
   alphaCSR[ 151 ][ 137 ],
   alphaCSR[ 151 ][ 138 ],
   alphaCSR[ 151 ][ 139 ],
   alphaCSR[ 151 ][ 140 ],
   alphaCSR[ 151 ][ 141 ],
   alphaCSR[ 151 ][ 142 ],
   alphaCSR[ 151 ][ 143 ],
   alphaCSR[ 151 ][ 144 ],
   alphaCSR[ 151 ][ 145 ],
   alphaCSR[ 151 ][ 146 ],
   alphaCSR[ 151 ][ 147 ],
   alphaCSR[ 151 ][ 148 ],
   alphaCSR[ 151 ][ 149 ],
   alphaCSR[ 151 ][ 150 ],
   alphaCSR[ 151 ][ 151 ],
   alphaCSR[ 151 ][ 152 ],
   alphaCSR[ 151 ][ 153 ],
   alphaCSR[ 151 ][ 154 ],
   alphaCSR[ 151 ][ 155 ],
   alphaCSR[ 151 ][ 156 ],
   alphaCSR[ 151 ][ 157 ],
   alphaCSR[ 151 ][ 158 ],
   alphaCSR[ 151 ][ 159 ],
   alphaCSR[ 151 ][ 160 ],
   alphaCSR[ 151 ][ 161 ],
   alphaCSR[ 151 ][ 162 ],
   alphaCSR[ 151 ][ 163 ],
   alphaCSR[ 151 ][ 164 ],
   alphaCSR[ 151 ][ 165 ],
   alphaCSR[ 151 ][ 166 ],
   alphaCSR[ 151 ][ 167 ],
   alphaCSR[ 151 ][ 168 ],
   alphaCSR[ 151 ][ 169 ],
   alphaCSR[ 151 ][ 170 ],
   alphaCSR[ 151 ][ 171 ],
   alphaCSR[ 151 ][ 172 ],
   alphaCSR[ 151 ][ 173 ],
   alphaCSR[ 151 ][ 174 ],
   alphaCSR[ 151 ][ 175 ],
   alphaCSR[ 151 ][ 176 ],
   alphaCSR[ 151 ][ 177 ],
   alphaCSR[ 151 ][ 178 ],
   alphaCSR[ 151 ][ 179 ],
   alphaCSR[ 151 ][ 180 ],
   alphaCSR[ 151 ][ 181 ],
   alphaCSR[ 151 ][ 182 ],
   alphaCSR[ 151 ][ 183 ],
   alphaCSR[ 151 ][ 184 ],
   alphaCSR[ 151 ][ 185 ],
   alphaCSR[ 151 ][ 186 ],
   alphaCSR[ 151 ][ 187 ],
   alphaCSR[ 151 ][ 188 ],
   alphaCSR[ 151 ][ 189 ],
   alphaCSR[ 151 ][ 190 ],
   alphaCSR[ 151 ][ 191 ],
   alphaCSR[ 151 ][ 192 ],
   alphaCSR[ 151 ][ 193 ],
   alphaCSR[ 151 ][ 194 ],
   alphaCSR[ 151 ][ 195 ],
   alphaCSR[ 151 ][ 196 ],
   alphaCSR[ 151 ][ 197 ],
   alphaCSR[ 151 ][ 198 ],
   alphaCSR[ 151 ][ 199 ],
   alphaCSR[ 151 ][ 200 ],
   alphaCSR[ 151 ][ 201 ],
   alphaCSR[ 151 ][ 202 ],
   alphaCSR[ 151 ][ 203 ],
   alphaCSR[ 151 ][ 204 ],
   alphaCSR[ 151 ][ 205 ],
   alphaCSR[ 151 ][ 206 ],
   alphaCSR[ 151 ][ 207 ],
   alphaCSR[ 151 ][ 208 ],
   alphaCSR[ 151 ][ 209 ],
   alphaCSR[ 151 ][ 210 ],
   alphaCSR[ 151 ][ 211 ],
   alphaCSR[ 151 ][ 212 ],
   alphaCSR[ 151 ][ 213 ],
   alphaCSR[ 151 ][ 214 ],
   alphaCSR[ 151 ][ 215 ],
   alphaCSR[ 151 ][ 216 ],
   alphaCSR[ 151 ][ 217 ],
   alphaCSR[ 151 ][ 218 ],
   alphaCSR[ 151 ][ 219 ],
   alphaCSR[ 151 ][ 220 ],
   alphaCSR[ 151 ][ 221 ],
   alphaCSR[ 151 ][ 222 ],
   alphaCSR[ 151 ][ 223 ],
   alphaCSR[ 151 ][ 224 ],
   alphaCSR[ 151 ][ 225 ],
   alphaCSR[ 151 ][ 226 ],
   alphaCSR[ 151 ][ 227 ],
   alphaCSR[ 151 ][ 228 ],
   alphaCSR[ 151 ][ 229 ],
   alphaCSR[ 151 ][ 230 ],
   alphaCSR[ 151 ][ 231 ],
   alphaCSR[ 151 ][ 232 ],
   alphaCSR[ 151 ][ 233 ],
   alphaCSR[ 151 ][ 234 ],
   alphaCSR[ 151 ][ 235 ],
   alphaCSR[ 151 ][ 236 ],
   alphaCSR[ 151 ][ 237 ],
   alphaCSR[ 151 ][ 238 ],
   alphaCSR[ 151 ][ 239 ],
   alphaCSR[ 151 ][ 240 ],
   alphaCSR[ 151 ][ 241 ],
   alphaCSR[ 151 ][ 242 ],
   alphaCSR[ 151 ][ 243 ],
   alphaCSR[ 151 ][ 244 ],
   alphaCSR[ 151 ][ 245 ],
   alphaCSR[ 151 ][ 246 ],
   alphaCSR[ 151 ][ 247 ],
   alphaCSR[ 151 ][ 248 ],
   alphaCSR[ 151 ][ 249 ],
   alphaCSR[ 151 ][ 250 ],
   alphaCSR[ 151 ][ 251 ],
   alphaCSR[ 151 ][ 252 ],
   alphaCSR[ 151 ][ 253 ],
   alphaCSR[ 151 ][ 254 ],
   alphaCSR[ 151 ][ 255 ],
   alphaCSR[ 151 ][ 256 ],
   alphaCSR[ 151 ][ 257 ],
   alphaCSR[ 151 ][ 258 ],
   alphaCSR[ 151 ][ 259 ],
   alphaCSR[ 151 ][ 260 ],
   alphaCSR[ 151 ][ 261 ],
   alphaCSR[ 151 ][ 262 ],
   alphaCSR[ 151 ][ 263 ],
   alphaCSR[ 151 ][ 264 ],
   alphaCSR[ 151 ][ 265 ],
   alphaCSR[ 151 ][ 266 ],
   alphaCSR[ 151 ][ 267 ],
   alphaCSR[ 151 ][ 268 ],
   alphaCSR[ 151 ][ 269 ],
   alphaCSR[ 151 ][ 270 ],
   alphaCSR[ 151 ][ 271 ],
   alphaCSR[ 151 ][ 272 ],
   alphaCSR[ 151 ][ 273 ],
   alphaCSR[ 151 ][ 274 ],
   alphaCSR[ 151 ][ 275 ],
   alphaCSR[ 151 ][ 276 ],
   alphaCSR[ 151 ][ 277 ],
   alphaCSR[ 151 ][ 278 ],
   alphaCSR[ 151 ][ 279 ],
   alphaCSR[ 151 ][ 280 ],
   alphaCSR[ 151 ][ 281 ],
   alphaCSR[ 151 ][ 282 ],
   alphaCSR[ 151 ][ 283 ],
   alphaCSR[ 151 ][ 284 ],
   alphaCSR[ 151 ][ 285 ],
   alphaCSR[ 151 ][ 286 ],
   alphaCSR[ 151 ][ 287 ],
   alphaCSR[ 151 ][ 288 ],
   alphaCSR[ 151 ][ 289 ],
   alphaCSR[ 151 ][ 290 ],
   alphaCSR[ 151 ][ 291 ],
   alphaCSR[ 151 ][ 292 ],
   alphaCSR[ 151 ][ 293 ],
   alphaCSR[ 151 ][ 294 ],
   alphaCSR[ 151 ][ 295 ],
   alphaCSR[ 151 ][ 296 ],
   alphaCSR[ 151 ][ 297 ],
   alphaCSR[ 151 ][ 298 ],
   alphaCSR[ 151 ][ 299 ],
   alphaCSR[ 151 ][ 300 ],
   alphaCSR[ 151 ][ 301 ],
   alphaCSR[ 151 ][ 302 ],
   alphaCSR[ 151 ][ 303 ],
   alphaCSR[ 151 ][ 304 ],
   alphaCSR[ 151 ][ 305 ],
   alphaCSR[ 151 ][ 306 ],
   alphaCSR[ 151 ][ 307 ],
   alphaCSR[ 151 ][ 308 ],
   alphaCSR[ 151 ][ 309 ],
   alphaCSR[ 151 ][ 310 ],
   alphaCSR[ 151 ][ 311 ],
   alphaCSR[ 151 ][ 312 ],
   alphaCSR[ 151 ][ 313 ],
   alphaCSR[ 151 ][ 314 ],
   alphaCSR[ 151 ][ 315 ],
   alphaCSR[ 151 ][ 316 ],
   alphaCSR[ 151 ][ 317 ],
   alphaCSR[ 151 ][ 318 ],
   alphaCSR[ 151 ][ 319 ],
   alphaCSR[ 151 ][ 320 ],
   alphaCSR[ 151 ][ 321 ],
   alphaCSR[ 151 ][ 322 ],
   alphaCSR[ 151 ][ 323 ],
   alphaCSR[ 151 ][ 324 ],
   alphaCSR[ 151 ][ 325 ],
   alphaCSR[ 151 ][ 326 ],
   alphaCSR[ 151 ][ 327 ],
   alphaCSR[ 151 ][ 328 ],
   alphaCSR[ 151 ][ 329 ],
   alphaCSR[ 151 ][ 330 ],
   alphaCSR[ 151 ][ 331 ],
   alphaCSR[ 151 ][ 332 ],
   alphaCSR[ 151 ][ 333 ],
   alphaCSR[ 151 ][ 334 ],
   alphaCSR[ 151 ][ 335 ],
   alphaCSR[ 151 ][ 336 ],
   alphaCSR[ 151 ][ 337 ],
   alphaCSR[ 151 ][ 338 ],
   alphaCSR[ 151 ][ 339 ],
   alphaCSR[ 151 ][ 340 ],
   alphaCSR[ 151 ][ 341 ],
   alphaCSR[ 151 ][ 342 ],
   alphaCSR[ 151 ][ 343 ],
   alphaCSR[ 151 ][ 344 ],
   alphaCSR[ 151 ][ 345 ],
   alphaCSR[ 151 ][ 346 ],
   alphaCSR[ 151 ][ 347 ],
   alphaCSR[ 151 ][ 348 ],
   alphaCSR[ 151 ][ 349 ],
   alphaCSR[ 151 ][ 350 ],
   alphaCSR[ 151 ][ 351 ],
   alphaCSR[ 151 ][ 352 ],
   alphaCSR[ 151 ][ 353 ],
   alphaCSR[ 151 ][ 354 ],
   alphaCSR[ 151 ][ 355 ],
   alphaCSR[ 151 ][ 356 ],
   alphaCSR[ 151 ][ 357 ],
   alphaCSR[ 151 ][ 358 ],
   alphaCSR[ 151 ][ 359 ],
   alphaCSR[ 151 ][ 360 ],
   alphaCSR[ 151 ][ 361 ],
   alphaCSR[ 151 ][ 362 ],
   alphaCSR[ 151 ][ 363 ],
   alphaCSR[ 151 ][ 364 ],
   alphaCSR[ 151 ][ 365 ],
   alphaCSR[ 151 ][ 366 ],
   alphaCSR[ 151 ][ 367 ],
   alphaCSR[ 151 ][ 368 ],
   alphaCSR[ 151 ][ 369 ],
   alphaCSR[ 151 ][ 370 ],
   alphaCSR[ 151 ][ 371 ],
   alphaCSR[ 151 ][ 372 ],
   alphaCSR[ 151 ][ 373 ],
   alphaCSR[ 151 ][ 374 ],
   alphaCSR[ 151 ][ 375 ],
   alphaCSR[ 151 ][ 376 ],
   alphaCSR[ 151 ][ 377 ],
   alphaCSR[ 151 ][ 378 ],
   alphaCSR[ 151 ][ 379 ],
   alphaCSR[ 151 ][ 380 ],
   alphaCSR[ 151 ][ 381 ],
   alphaCSR[ 151 ][ 382 ],
   alphaCSR[ 151 ][ 383 ],
   alphaCSR[ 152 ][ 0 ],
   alphaCSR[ 152 ][ 1 ],
   alphaCSR[ 152 ][ 2 ],
   alphaCSR[ 152 ][ 3 ],
   alphaCSR[ 152 ][ 4 ],
   alphaCSR[ 152 ][ 5 ],
   alphaCSR[ 152 ][ 6 ],
   alphaCSR[ 152 ][ 7 ],
   alphaCSR[ 152 ][ 8 ],
   alphaCSR[ 152 ][ 9 ],
   alphaCSR[ 152 ][ 10 ],
   alphaCSR[ 152 ][ 11 ],
   alphaCSR[ 152 ][ 12 ],
   alphaCSR[ 152 ][ 13 ],
   alphaCSR[ 152 ][ 14 ],
   alphaCSR[ 152 ][ 15 ],
   alphaCSR[ 152 ][ 16 ],
   alphaCSR[ 152 ][ 17 ],
   alphaCSR[ 152 ][ 18 ],
   alphaCSR[ 152 ][ 19 ],
   alphaCSR[ 152 ][ 20 ],
   alphaCSR[ 152 ][ 21 ],
   alphaCSR[ 152 ][ 22 ],
   alphaCSR[ 152 ][ 23 ],
   alphaCSR[ 152 ][ 24 ],
   alphaCSR[ 152 ][ 25 ],
   alphaCSR[ 152 ][ 26 ],
   alphaCSR[ 152 ][ 27 ],
   alphaCSR[ 152 ][ 28 ],
   alphaCSR[ 152 ][ 29 ],
   alphaCSR[ 152 ][ 30 ],
   alphaCSR[ 152 ][ 31 ],
   alphaCSR[ 152 ][ 32 ],
   alphaCSR[ 152 ][ 33 ],
   alphaCSR[ 152 ][ 34 ],
   alphaCSR[ 152 ][ 35 ],
   alphaCSR[ 152 ][ 36 ],
   alphaCSR[ 152 ][ 37 ],
   alphaCSR[ 152 ][ 38 ],
   alphaCSR[ 152 ][ 39 ],
   alphaCSR[ 152 ][ 40 ],
   alphaCSR[ 152 ][ 41 ],
   alphaCSR[ 152 ][ 42 ],
   alphaCSR[ 152 ][ 43 ],
   alphaCSR[ 152 ][ 44 ],
   alphaCSR[ 152 ][ 45 ],
   alphaCSR[ 152 ][ 46 ],
   alphaCSR[ 152 ][ 47 ],
   alphaCSR[ 152 ][ 48 ],
   alphaCSR[ 152 ][ 49 ],
   alphaCSR[ 152 ][ 50 ],
   alphaCSR[ 152 ][ 51 ],
   alphaCSR[ 152 ][ 52 ],
   alphaCSR[ 152 ][ 53 ],
   alphaCSR[ 152 ][ 54 ],
   alphaCSR[ 152 ][ 55 ],
   alphaCSR[ 152 ][ 56 ],
   alphaCSR[ 152 ][ 57 ],
   alphaCSR[ 152 ][ 58 ],
   alphaCSR[ 152 ][ 59 ],
   alphaCSR[ 152 ][ 60 ],
   alphaCSR[ 152 ][ 61 ],
   alphaCSR[ 152 ][ 62 ],
   alphaCSR[ 152 ][ 63 ],
   alphaCSR[ 152 ][ 64 ],
   alphaCSR[ 152 ][ 65 ],
   alphaCSR[ 152 ][ 66 ],
   alphaCSR[ 152 ][ 67 ],
   alphaCSR[ 152 ][ 68 ],
   alphaCSR[ 152 ][ 69 ],
   alphaCSR[ 152 ][ 70 ],
   alphaCSR[ 152 ][ 71 ],
   alphaCSR[ 152 ][ 72 ],
   alphaCSR[ 152 ][ 73 ],
   alphaCSR[ 152 ][ 74 ],
   alphaCSR[ 152 ][ 75 ],
   alphaCSR[ 152 ][ 76 ],
   alphaCSR[ 152 ][ 77 ],
   alphaCSR[ 152 ][ 78 ],
   alphaCSR[ 152 ][ 79 ],
   alphaCSR[ 152 ][ 80 ],
   alphaCSR[ 152 ][ 81 ],
   alphaCSR[ 152 ][ 82 ],
   alphaCSR[ 152 ][ 83 ],
   alphaCSR[ 152 ][ 84 ],
   alphaCSR[ 152 ][ 85 ],
   alphaCSR[ 152 ][ 86 ],
   alphaCSR[ 152 ][ 87 ],
   alphaCSR[ 152 ][ 88 ],
   alphaCSR[ 152 ][ 89 ],
   alphaCSR[ 152 ][ 90 ],
   alphaCSR[ 152 ][ 91 ],
   alphaCSR[ 152 ][ 92 ],
   alphaCSR[ 152 ][ 93 ],
   alphaCSR[ 152 ][ 94 ],
   alphaCSR[ 152 ][ 95 ],
   alphaCSR[ 152 ][ 96 ],
   alphaCSR[ 152 ][ 97 ],
   alphaCSR[ 152 ][ 98 ],
   alphaCSR[ 152 ][ 99 ],
   alphaCSR[ 152 ][ 100 ],
   alphaCSR[ 152 ][ 101 ],
   alphaCSR[ 152 ][ 102 ],
   alphaCSR[ 152 ][ 103 ],
   alphaCSR[ 152 ][ 104 ],
   alphaCSR[ 152 ][ 105 ],
   alphaCSR[ 152 ][ 106 ],
   alphaCSR[ 152 ][ 107 ],
   alphaCSR[ 152 ][ 108 ],
   alphaCSR[ 152 ][ 109 ],
   alphaCSR[ 152 ][ 110 ],
   alphaCSR[ 152 ][ 111 ],
   alphaCSR[ 152 ][ 112 ],
   alphaCSR[ 152 ][ 113 ],
   alphaCSR[ 152 ][ 114 ],
   alphaCSR[ 152 ][ 115 ],
   alphaCSR[ 152 ][ 116 ],
   alphaCSR[ 152 ][ 117 ],
   alphaCSR[ 152 ][ 118 ],
   alphaCSR[ 152 ][ 119 ],
   alphaCSR[ 152 ][ 120 ],
   alphaCSR[ 152 ][ 121 ],
   alphaCSR[ 152 ][ 122 ],
   alphaCSR[ 152 ][ 123 ],
   alphaCSR[ 152 ][ 124 ],
   alphaCSR[ 152 ][ 125 ],
   alphaCSR[ 152 ][ 126 ],
   alphaCSR[ 152 ][ 127 ],
   alphaCSR[ 152 ][ 128 ],
   alphaCSR[ 152 ][ 129 ],
   alphaCSR[ 152 ][ 130 ],
   alphaCSR[ 152 ][ 131 ],
   alphaCSR[ 152 ][ 132 ],
   alphaCSR[ 152 ][ 133 ],
   alphaCSR[ 152 ][ 134 ],
   alphaCSR[ 152 ][ 135 ],
   alphaCSR[ 152 ][ 136 ],
   alphaCSR[ 152 ][ 137 ],
   alphaCSR[ 152 ][ 138 ],
   alphaCSR[ 152 ][ 139 ],
   alphaCSR[ 152 ][ 140 ],
   alphaCSR[ 152 ][ 141 ],
   alphaCSR[ 152 ][ 142 ],
   alphaCSR[ 152 ][ 143 ],
   alphaCSR[ 152 ][ 144 ],
   alphaCSR[ 152 ][ 145 ],
   alphaCSR[ 152 ][ 146 ],
   alphaCSR[ 152 ][ 147 ],
   alphaCSR[ 152 ][ 148 ],
   alphaCSR[ 152 ][ 149 ],
   alphaCSR[ 152 ][ 150 ],
   alphaCSR[ 152 ][ 151 ],
   alphaCSR[ 152 ][ 152 ],
   alphaCSR[ 152 ][ 153 ],
   alphaCSR[ 152 ][ 154 ],
   alphaCSR[ 152 ][ 155 ],
   alphaCSR[ 152 ][ 156 ],
   alphaCSR[ 152 ][ 157 ],
   alphaCSR[ 152 ][ 158 ],
   alphaCSR[ 152 ][ 159 ],
   alphaCSR[ 152 ][ 160 ],
   alphaCSR[ 152 ][ 161 ],
   alphaCSR[ 152 ][ 162 ],
   alphaCSR[ 152 ][ 163 ],
   alphaCSR[ 152 ][ 164 ],
   alphaCSR[ 152 ][ 165 ],
   alphaCSR[ 152 ][ 166 ],
   alphaCSR[ 152 ][ 167 ],
   alphaCSR[ 152 ][ 168 ],
   alphaCSR[ 152 ][ 169 ],
   alphaCSR[ 152 ][ 170 ],
   alphaCSR[ 152 ][ 171 ],
   alphaCSR[ 152 ][ 172 ],
   alphaCSR[ 152 ][ 173 ],
   alphaCSR[ 152 ][ 174 ],
   alphaCSR[ 152 ][ 175 ],
   alphaCSR[ 152 ][ 176 ],
   alphaCSR[ 152 ][ 177 ],
   alphaCSR[ 152 ][ 178 ],
   alphaCSR[ 152 ][ 179 ],
   alphaCSR[ 152 ][ 180 ],
   alphaCSR[ 152 ][ 181 ],
   alphaCSR[ 152 ][ 182 ],
   alphaCSR[ 152 ][ 183 ],
   alphaCSR[ 152 ][ 184 ],
   alphaCSR[ 152 ][ 185 ],
   alphaCSR[ 152 ][ 186 ],
   alphaCSR[ 152 ][ 187 ],
   alphaCSR[ 152 ][ 188 ],
   alphaCSR[ 152 ][ 189 ],
   alphaCSR[ 152 ][ 190 ],
   alphaCSR[ 152 ][ 191 ],
   alphaCSR[ 152 ][ 192 ],
   alphaCSR[ 152 ][ 193 ],
   alphaCSR[ 152 ][ 194 ],
   alphaCSR[ 152 ][ 195 ],
   alphaCSR[ 152 ][ 196 ],
   alphaCSR[ 152 ][ 197 ],
   alphaCSR[ 152 ][ 198 ],
   alphaCSR[ 152 ][ 199 ],
   alphaCSR[ 152 ][ 200 ],
   alphaCSR[ 152 ][ 201 ],
   alphaCSR[ 152 ][ 202 ],
   alphaCSR[ 152 ][ 203 ],
   alphaCSR[ 152 ][ 204 ],
   alphaCSR[ 152 ][ 205 ],
   alphaCSR[ 152 ][ 206 ],
   alphaCSR[ 152 ][ 207 ],
   alphaCSR[ 152 ][ 208 ],
   alphaCSR[ 152 ][ 209 ],
   alphaCSR[ 152 ][ 210 ],
   alphaCSR[ 152 ][ 211 ],
   alphaCSR[ 152 ][ 212 ],
   alphaCSR[ 152 ][ 213 ],
   alphaCSR[ 152 ][ 214 ],
   alphaCSR[ 152 ][ 215 ],
   alphaCSR[ 152 ][ 216 ],
   alphaCSR[ 152 ][ 217 ],
   alphaCSR[ 152 ][ 218 ],
   alphaCSR[ 152 ][ 219 ],
   alphaCSR[ 152 ][ 220 ],
   alphaCSR[ 152 ][ 221 ],
   alphaCSR[ 152 ][ 222 ],
   alphaCSR[ 152 ][ 223 ],
   alphaCSR[ 152 ][ 224 ],
   alphaCSR[ 152 ][ 225 ],
   alphaCSR[ 152 ][ 226 ],
   alphaCSR[ 152 ][ 227 ],
   alphaCSR[ 152 ][ 228 ],
   alphaCSR[ 152 ][ 229 ],
   alphaCSR[ 152 ][ 230 ],
   alphaCSR[ 152 ][ 231 ],
   alphaCSR[ 152 ][ 232 ],
   alphaCSR[ 152 ][ 233 ],
   alphaCSR[ 152 ][ 234 ],
   alphaCSR[ 152 ][ 235 ],
   alphaCSR[ 152 ][ 236 ],
   alphaCSR[ 152 ][ 237 ],
   alphaCSR[ 152 ][ 238 ],
   alphaCSR[ 152 ][ 239 ],
   alphaCSR[ 152 ][ 240 ],
   alphaCSR[ 152 ][ 241 ],
   alphaCSR[ 152 ][ 242 ],
   alphaCSR[ 152 ][ 243 ],
   alphaCSR[ 152 ][ 244 ],
   alphaCSR[ 152 ][ 245 ],
   alphaCSR[ 152 ][ 246 ],
   alphaCSR[ 152 ][ 247 ],
   alphaCSR[ 152 ][ 248 ],
   alphaCSR[ 152 ][ 249 ],
   alphaCSR[ 152 ][ 250 ],
   alphaCSR[ 152 ][ 251 ],
   alphaCSR[ 152 ][ 252 ],
   alphaCSR[ 152 ][ 253 ],
   alphaCSR[ 152 ][ 254 ],
   alphaCSR[ 152 ][ 255 ],
   alphaCSR[ 152 ][ 256 ],
   alphaCSR[ 152 ][ 257 ],
   alphaCSR[ 152 ][ 258 ],
   alphaCSR[ 152 ][ 259 ],
   alphaCSR[ 152 ][ 260 ],
   alphaCSR[ 152 ][ 261 ],
   alphaCSR[ 152 ][ 262 ],
   alphaCSR[ 152 ][ 263 ],
   alphaCSR[ 152 ][ 264 ],
   alphaCSR[ 152 ][ 265 ],
   alphaCSR[ 152 ][ 266 ],
   alphaCSR[ 152 ][ 267 ],
   alphaCSR[ 152 ][ 268 ],
   alphaCSR[ 152 ][ 269 ],
   alphaCSR[ 152 ][ 270 ],
   alphaCSR[ 152 ][ 271 ],
   alphaCSR[ 152 ][ 272 ],
   alphaCSR[ 152 ][ 273 ],
   alphaCSR[ 152 ][ 274 ],
   alphaCSR[ 152 ][ 275 ],
   alphaCSR[ 152 ][ 276 ],
   alphaCSR[ 152 ][ 277 ],
   alphaCSR[ 152 ][ 278 ],
   alphaCSR[ 152 ][ 279 ],
   alphaCSR[ 152 ][ 280 ],
   alphaCSR[ 152 ][ 281 ],
   alphaCSR[ 152 ][ 282 ],
   alphaCSR[ 152 ][ 283 ],
   alphaCSR[ 152 ][ 284 ],
   alphaCSR[ 152 ][ 285 ],
   alphaCSR[ 152 ][ 286 ],
   alphaCSR[ 152 ][ 287 ],
   alphaCSR[ 152 ][ 288 ],
   alphaCSR[ 152 ][ 289 ],
   alphaCSR[ 152 ][ 290 ],
   alphaCSR[ 152 ][ 291 ],
   alphaCSR[ 152 ][ 292 ],
   alphaCSR[ 152 ][ 293 ],
   alphaCSR[ 152 ][ 294 ],
   alphaCSR[ 152 ][ 295 ],
   alphaCSR[ 152 ][ 296 ],
   alphaCSR[ 152 ][ 297 ],
   alphaCSR[ 152 ][ 298 ],
   alphaCSR[ 152 ][ 299 ],
   alphaCSR[ 152 ][ 300 ],
   alphaCSR[ 152 ][ 301 ],
   alphaCSR[ 152 ][ 302 ],
   alphaCSR[ 152 ][ 303 ],
   alphaCSR[ 152 ][ 304 ],
   alphaCSR[ 152 ][ 305 ],
   alphaCSR[ 152 ][ 306 ],
   alphaCSR[ 152 ][ 307 ],
   alphaCSR[ 152 ][ 308 ],
   alphaCSR[ 152 ][ 309 ],
   alphaCSR[ 152 ][ 310 ],
   alphaCSR[ 152 ][ 311 ],
   alphaCSR[ 152 ][ 312 ],
   alphaCSR[ 152 ][ 313 ],
   alphaCSR[ 152 ][ 314 ],
   alphaCSR[ 152 ][ 315 ],
   alphaCSR[ 152 ][ 316 ],
   alphaCSR[ 152 ][ 317 ],
   alphaCSR[ 152 ][ 318 ],
   alphaCSR[ 152 ][ 319 ],
   alphaCSR[ 152 ][ 320 ],
   alphaCSR[ 152 ][ 321 ],
   alphaCSR[ 152 ][ 322 ],
   alphaCSR[ 152 ][ 323 ],
   alphaCSR[ 152 ][ 324 ],
   alphaCSR[ 152 ][ 325 ],
   alphaCSR[ 152 ][ 326 ],
   alphaCSR[ 152 ][ 327 ],
   alphaCSR[ 152 ][ 328 ],
   alphaCSR[ 152 ][ 329 ],
   alphaCSR[ 152 ][ 330 ],
   alphaCSR[ 152 ][ 331 ],
   alphaCSR[ 152 ][ 332 ],
   alphaCSR[ 152 ][ 333 ],
   alphaCSR[ 152 ][ 334 ],
   alphaCSR[ 152 ][ 335 ],
   alphaCSR[ 152 ][ 336 ],
   alphaCSR[ 152 ][ 337 ],
   alphaCSR[ 152 ][ 338 ],
   alphaCSR[ 152 ][ 339 ],
   alphaCSR[ 152 ][ 340 ],
   alphaCSR[ 152 ][ 341 ],
   alphaCSR[ 152 ][ 342 ],
   alphaCSR[ 152 ][ 343 ],
   alphaCSR[ 152 ][ 344 ],
   alphaCSR[ 152 ][ 345 ],
   alphaCSR[ 152 ][ 346 ],
   alphaCSR[ 152 ][ 347 ],
   alphaCSR[ 152 ][ 348 ],
   alphaCSR[ 152 ][ 349 ],
   alphaCSR[ 152 ][ 350 ],
   alphaCSR[ 152 ][ 351 ],
   alphaCSR[ 152 ][ 352 ],
   alphaCSR[ 152 ][ 353 ],
   alphaCSR[ 152 ][ 354 ],
   alphaCSR[ 152 ][ 355 ],
   alphaCSR[ 152 ][ 356 ],
   alphaCSR[ 152 ][ 357 ],
   alphaCSR[ 152 ][ 358 ],
   alphaCSR[ 152 ][ 359 ],
   alphaCSR[ 152 ][ 360 ],
   alphaCSR[ 152 ][ 361 ],
   alphaCSR[ 152 ][ 362 ],
   alphaCSR[ 152 ][ 363 ],
   alphaCSR[ 152 ][ 364 ],
   alphaCSR[ 152 ][ 365 ],
   alphaCSR[ 152 ][ 366 ],
   alphaCSR[ 152 ][ 367 ],
   alphaCSR[ 152 ][ 368 ],
   alphaCSR[ 152 ][ 369 ],
   alphaCSR[ 152 ][ 370 ],
   alphaCSR[ 152 ][ 371 ],
   alphaCSR[ 152 ][ 372 ],
   alphaCSR[ 152 ][ 373 ],
   alphaCSR[ 152 ][ 374 ],
   alphaCSR[ 152 ][ 375 ],
   alphaCSR[ 152 ][ 376 ],
   alphaCSR[ 152 ][ 377 ],
   alphaCSR[ 152 ][ 378 ],
   alphaCSR[ 152 ][ 379 ],
   alphaCSR[ 152 ][ 380 ],
   alphaCSR[ 152 ][ 381 ],
   alphaCSR[ 152 ][ 382 ],
   alphaCSR[ 152 ][ 383 ],
   alphaCSR[ 153 ][ 0 ],
   alphaCSR[ 153 ][ 1 ],
   alphaCSR[ 153 ][ 2 ],
   alphaCSR[ 153 ][ 3 ],
   alphaCSR[ 153 ][ 4 ],
   alphaCSR[ 153 ][ 5 ],
   alphaCSR[ 153 ][ 6 ],
   alphaCSR[ 153 ][ 7 ],
   alphaCSR[ 153 ][ 8 ],
   alphaCSR[ 153 ][ 9 ],
   alphaCSR[ 153 ][ 10 ],
   alphaCSR[ 153 ][ 11 ],
   alphaCSR[ 153 ][ 12 ],
   alphaCSR[ 153 ][ 13 ],
   alphaCSR[ 153 ][ 14 ],
   alphaCSR[ 153 ][ 15 ],
   alphaCSR[ 153 ][ 16 ],
   alphaCSR[ 153 ][ 17 ],
   alphaCSR[ 153 ][ 18 ],
   alphaCSR[ 153 ][ 19 ],
   alphaCSR[ 153 ][ 20 ],
   alphaCSR[ 153 ][ 21 ],
   alphaCSR[ 153 ][ 22 ],
   alphaCSR[ 153 ][ 23 ],
   alphaCSR[ 153 ][ 24 ],
   alphaCSR[ 153 ][ 25 ],
   alphaCSR[ 153 ][ 26 ],
   alphaCSR[ 153 ][ 27 ],
   alphaCSR[ 153 ][ 28 ],
   alphaCSR[ 153 ][ 29 ],
   alphaCSR[ 153 ][ 30 ],
   alphaCSR[ 153 ][ 31 ],
   alphaCSR[ 153 ][ 32 ],
   alphaCSR[ 153 ][ 33 ],
   alphaCSR[ 153 ][ 34 ],
   alphaCSR[ 153 ][ 35 ],
   alphaCSR[ 153 ][ 36 ],
   alphaCSR[ 153 ][ 37 ],
   alphaCSR[ 153 ][ 38 ],
   alphaCSR[ 153 ][ 39 ],
   alphaCSR[ 153 ][ 40 ],
   alphaCSR[ 153 ][ 41 ],
   alphaCSR[ 153 ][ 42 ],
   alphaCSR[ 153 ][ 43 ],
   alphaCSR[ 153 ][ 44 ],
   alphaCSR[ 153 ][ 45 ],
   alphaCSR[ 153 ][ 46 ],
   alphaCSR[ 153 ][ 47 ],
   alphaCSR[ 153 ][ 48 ],
   alphaCSR[ 153 ][ 49 ],
   alphaCSR[ 153 ][ 50 ],
   alphaCSR[ 153 ][ 51 ],
   alphaCSR[ 153 ][ 52 ],
   alphaCSR[ 153 ][ 53 ],
   alphaCSR[ 153 ][ 54 ],
   alphaCSR[ 153 ][ 55 ],
   alphaCSR[ 153 ][ 56 ],
   alphaCSR[ 153 ][ 57 ],
   alphaCSR[ 153 ][ 58 ],
   alphaCSR[ 153 ][ 59 ],
   alphaCSR[ 153 ][ 60 ],
   alphaCSR[ 153 ][ 61 ],
   alphaCSR[ 153 ][ 62 ],
   alphaCSR[ 153 ][ 63 ],
   alphaCSR[ 153 ][ 64 ],
   alphaCSR[ 153 ][ 65 ],
   alphaCSR[ 153 ][ 66 ],
   alphaCSR[ 153 ][ 67 ],
   alphaCSR[ 153 ][ 68 ],
   alphaCSR[ 153 ][ 69 ],
   alphaCSR[ 153 ][ 70 ],
   alphaCSR[ 153 ][ 71 ],
   alphaCSR[ 153 ][ 72 ],
   alphaCSR[ 153 ][ 73 ],
   alphaCSR[ 153 ][ 74 ],
   alphaCSR[ 153 ][ 75 ],
   alphaCSR[ 153 ][ 76 ],
   alphaCSR[ 153 ][ 77 ],
   alphaCSR[ 153 ][ 78 ],
   alphaCSR[ 153 ][ 79 ],
   alphaCSR[ 153 ][ 80 ],
   alphaCSR[ 153 ][ 81 ],
   alphaCSR[ 153 ][ 82 ],
   alphaCSR[ 153 ][ 83 ],
   alphaCSR[ 153 ][ 84 ],
   alphaCSR[ 153 ][ 85 ],
   alphaCSR[ 153 ][ 86 ],
   alphaCSR[ 153 ][ 87 ],
   alphaCSR[ 153 ][ 88 ],
   alphaCSR[ 153 ][ 89 ],
   alphaCSR[ 153 ][ 90 ],
   alphaCSR[ 153 ][ 91 ],
   alphaCSR[ 153 ][ 92 ],
   alphaCSR[ 153 ][ 93 ],
   alphaCSR[ 153 ][ 94 ],
   alphaCSR[ 153 ][ 95 ],
   alphaCSR[ 153 ][ 96 ],
   alphaCSR[ 153 ][ 97 ],
   alphaCSR[ 153 ][ 98 ],
   alphaCSR[ 153 ][ 99 ],
   alphaCSR[ 153 ][ 100 ],
   alphaCSR[ 153 ][ 101 ],
   alphaCSR[ 153 ][ 102 ],
   alphaCSR[ 153 ][ 103 ],
   alphaCSR[ 153 ][ 104 ],
   alphaCSR[ 153 ][ 105 ],
   alphaCSR[ 153 ][ 106 ],
   alphaCSR[ 153 ][ 107 ],
   alphaCSR[ 153 ][ 108 ],
   alphaCSR[ 153 ][ 109 ],
   alphaCSR[ 153 ][ 110 ],
   alphaCSR[ 153 ][ 111 ],
   alphaCSR[ 153 ][ 112 ],
   alphaCSR[ 153 ][ 113 ],
   alphaCSR[ 153 ][ 114 ],
   alphaCSR[ 153 ][ 115 ],
   alphaCSR[ 153 ][ 116 ],
   alphaCSR[ 153 ][ 117 ],
   alphaCSR[ 153 ][ 118 ],
   alphaCSR[ 153 ][ 119 ],
   alphaCSR[ 153 ][ 120 ],
   alphaCSR[ 153 ][ 121 ],
   alphaCSR[ 153 ][ 122 ],
   alphaCSR[ 153 ][ 123 ],
   alphaCSR[ 153 ][ 124 ],
   alphaCSR[ 153 ][ 125 ],
   alphaCSR[ 153 ][ 126 ],
   alphaCSR[ 153 ][ 127 ],
   alphaCSR[ 153 ][ 128 ],
   alphaCSR[ 153 ][ 129 ],
   alphaCSR[ 153 ][ 130 ],
   alphaCSR[ 153 ][ 131 ],
   alphaCSR[ 153 ][ 132 ],
   alphaCSR[ 153 ][ 133 ],
   alphaCSR[ 153 ][ 134 ],
   alphaCSR[ 153 ][ 135 ],
   alphaCSR[ 153 ][ 136 ],
   alphaCSR[ 153 ][ 137 ],
   alphaCSR[ 153 ][ 138 ],
   alphaCSR[ 153 ][ 139 ],
   alphaCSR[ 153 ][ 140 ],
   alphaCSR[ 153 ][ 141 ],
   alphaCSR[ 153 ][ 142 ],
   alphaCSR[ 153 ][ 143 ],
   alphaCSR[ 153 ][ 144 ],
   alphaCSR[ 153 ][ 145 ],
   alphaCSR[ 153 ][ 146 ],
   alphaCSR[ 153 ][ 147 ],
   alphaCSR[ 153 ][ 148 ],
   alphaCSR[ 153 ][ 149 ],
   alphaCSR[ 153 ][ 150 ],
   alphaCSR[ 153 ][ 151 ],
   alphaCSR[ 153 ][ 152 ],
   alphaCSR[ 153 ][ 153 ],
   alphaCSR[ 153 ][ 154 ],
   alphaCSR[ 153 ][ 155 ],
   alphaCSR[ 153 ][ 156 ],
   alphaCSR[ 153 ][ 157 ],
   alphaCSR[ 153 ][ 158 ],
   alphaCSR[ 153 ][ 159 ],
   alphaCSR[ 153 ][ 160 ],
   alphaCSR[ 153 ][ 161 ],
   alphaCSR[ 153 ][ 162 ],
   alphaCSR[ 153 ][ 163 ],
   alphaCSR[ 153 ][ 164 ],
   alphaCSR[ 153 ][ 165 ],
   alphaCSR[ 153 ][ 166 ],
   alphaCSR[ 153 ][ 167 ],
   alphaCSR[ 153 ][ 168 ],
   alphaCSR[ 153 ][ 169 ],
   alphaCSR[ 153 ][ 170 ],
   alphaCSR[ 153 ][ 171 ],
   alphaCSR[ 153 ][ 172 ],
   alphaCSR[ 153 ][ 173 ],
   alphaCSR[ 153 ][ 174 ],
   alphaCSR[ 153 ][ 175 ],
   alphaCSR[ 153 ][ 176 ],
   alphaCSR[ 153 ][ 177 ],
   alphaCSR[ 153 ][ 178 ],
   alphaCSR[ 153 ][ 179 ],
   alphaCSR[ 153 ][ 180 ],
   alphaCSR[ 153 ][ 181 ],
   alphaCSR[ 153 ][ 182 ],
   alphaCSR[ 153 ][ 183 ],
   alphaCSR[ 153 ][ 184 ],
   alphaCSR[ 153 ][ 185 ],
   alphaCSR[ 153 ][ 186 ],
   alphaCSR[ 153 ][ 187 ],
   alphaCSR[ 153 ][ 188 ],
   alphaCSR[ 153 ][ 189 ],
   alphaCSR[ 153 ][ 190 ],
   alphaCSR[ 153 ][ 191 ],
   alphaCSR[ 153 ][ 192 ],
   alphaCSR[ 153 ][ 193 ],
   alphaCSR[ 153 ][ 194 ],
   alphaCSR[ 153 ][ 195 ],
   alphaCSR[ 153 ][ 196 ],
   alphaCSR[ 153 ][ 197 ],
   alphaCSR[ 153 ][ 198 ],
   alphaCSR[ 153 ][ 199 ],
   alphaCSR[ 153 ][ 200 ],
   alphaCSR[ 153 ][ 201 ],
   alphaCSR[ 153 ][ 202 ],
   alphaCSR[ 153 ][ 203 ],
   alphaCSR[ 153 ][ 204 ],
   alphaCSR[ 153 ][ 205 ],
   alphaCSR[ 153 ][ 206 ],
   alphaCSR[ 153 ][ 207 ],
   alphaCSR[ 153 ][ 208 ],
   alphaCSR[ 153 ][ 209 ],
   alphaCSR[ 153 ][ 210 ],
   alphaCSR[ 153 ][ 211 ],
   alphaCSR[ 153 ][ 212 ],
   alphaCSR[ 153 ][ 213 ],
   alphaCSR[ 153 ][ 214 ],
   alphaCSR[ 153 ][ 215 ],
   alphaCSR[ 153 ][ 216 ],
   alphaCSR[ 153 ][ 217 ],
   alphaCSR[ 153 ][ 218 ],
   alphaCSR[ 153 ][ 219 ],
   alphaCSR[ 153 ][ 220 ],
   alphaCSR[ 153 ][ 221 ],
   alphaCSR[ 153 ][ 222 ],
   alphaCSR[ 153 ][ 223 ],
   alphaCSR[ 153 ][ 224 ],
   alphaCSR[ 153 ][ 225 ],
   alphaCSR[ 153 ][ 226 ],
   alphaCSR[ 153 ][ 227 ],
   alphaCSR[ 153 ][ 228 ],
   alphaCSR[ 153 ][ 229 ],
   alphaCSR[ 153 ][ 230 ],
   alphaCSR[ 153 ][ 231 ],
   alphaCSR[ 153 ][ 232 ],
   alphaCSR[ 153 ][ 233 ],
   alphaCSR[ 153 ][ 234 ],
   alphaCSR[ 153 ][ 235 ],
   alphaCSR[ 153 ][ 236 ],
   alphaCSR[ 153 ][ 237 ],
   alphaCSR[ 153 ][ 238 ],
   alphaCSR[ 153 ][ 239 ],
   alphaCSR[ 153 ][ 240 ],
   alphaCSR[ 153 ][ 241 ],
   alphaCSR[ 153 ][ 242 ],
   alphaCSR[ 153 ][ 243 ],
   alphaCSR[ 153 ][ 244 ],
   alphaCSR[ 153 ][ 245 ],
   alphaCSR[ 153 ][ 246 ],
   alphaCSR[ 153 ][ 247 ],
   alphaCSR[ 153 ][ 248 ],
   alphaCSR[ 153 ][ 249 ],
   alphaCSR[ 153 ][ 250 ],
   alphaCSR[ 153 ][ 251 ],
   alphaCSR[ 153 ][ 252 ],
   alphaCSR[ 153 ][ 253 ],
   alphaCSR[ 153 ][ 254 ],
   alphaCSR[ 153 ][ 255 ],
   alphaCSR[ 153 ][ 256 ],
   alphaCSR[ 153 ][ 257 ],
   alphaCSR[ 153 ][ 258 ],
   alphaCSR[ 153 ][ 259 ],
   alphaCSR[ 153 ][ 260 ],
   alphaCSR[ 153 ][ 261 ],
   alphaCSR[ 153 ][ 262 ],
   alphaCSR[ 153 ][ 263 ],
   alphaCSR[ 153 ][ 264 ],
   alphaCSR[ 153 ][ 265 ],
   alphaCSR[ 153 ][ 266 ],
   alphaCSR[ 153 ][ 267 ],
   alphaCSR[ 153 ][ 268 ],
   alphaCSR[ 153 ][ 269 ],
   alphaCSR[ 153 ][ 270 ],
   alphaCSR[ 153 ][ 271 ],
   alphaCSR[ 153 ][ 272 ],
   alphaCSR[ 153 ][ 273 ],
   alphaCSR[ 153 ][ 274 ],
   alphaCSR[ 153 ][ 275 ],
   alphaCSR[ 153 ][ 276 ],
   alphaCSR[ 153 ][ 277 ],
   alphaCSR[ 153 ][ 278 ],
   alphaCSR[ 153 ][ 279 ],
   alphaCSR[ 153 ][ 280 ],
   alphaCSR[ 153 ][ 281 ],
   alphaCSR[ 153 ][ 282 ],
   alphaCSR[ 153 ][ 283 ],
   alphaCSR[ 153 ][ 284 ],
   alphaCSR[ 153 ][ 285 ],
   alphaCSR[ 153 ][ 286 ],
   alphaCSR[ 153 ][ 287 ],
   alphaCSR[ 153 ][ 288 ],
   alphaCSR[ 153 ][ 289 ],
   alphaCSR[ 153 ][ 290 ],
   alphaCSR[ 153 ][ 291 ],
   alphaCSR[ 153 ][ 292 ],
   alphaCSR[ 153 ][ 293 ],
   alphaCSR[ 153 ][ 294 ],
   alphaCSR[ 153 ][ 295 ],
   alphaCSR[ 153 ][ 296 ],
   alphaCSR[ 153 ][ 297 ],
   alphaCSR[ 153 ][ 298 ],
   alphaCSR[ 153 ][ 299 ],
   alphaCSR[ 153 ][ 300 ],
   alphaCSR[ 153 ][ 301 ],
   alphaCSR[ 153 ][ 302 ],
   alphaCSR[ 153 ][ 303 ],
   alphaCSR[ 153 ][ 304 ],
   alphaCSR[ 153 ][ 305 ],
   alphaCSR[ 153 ][ 306 ],
   alphaCSR[ 153 ][ 307 ],
   alphaCSR[ 153 ][ 308 ],
   alphaCSR[ 153 ][ 309 ],
   alphaCSR[ 153 ][ 310 ],
   alphaCSR[ 153 ][ 311 ],
   alphaCSR[ 153 ][ 312 ],
   alphaCSR[ 153 ][ 313 ],
   alphaCSR[ 153 ][ 314 ],
   alphaCSR[ 153 ][ 315 ],
   alphaCSR[ 153 ][ 316 ],
   alphaCSR[ 153 ][ 317 ],
   alphaCSR[ 153 ][ 318 ],
   alphaCSR[ 153 ][ 319 ],
   alphaCSR[ 153 ][ 320 ],
   alphaCSR[ 153 ][ 321 ],
   alphaCSR[ 153 ][ 322 ],
   alphaCSR[ 153 ][ 323 ],
   alphaCSR[ 153 ][ 324 ],
   alphaCSR[ 153 ][ 325 ],
   alphaCSR[ 153 ][ 326 ],
   alphaCSR[ 153 ][ 327 ],
   alphaCSR[ 153 ][ 328 ],
   alphaCSR[ 153 ][ 329 ],
   alphaCSR[ 153 ][ 330 ],
   alphaCSR[ 153 ][ 331 ],
   alphaCSR[ 153 ][ 332 ],
   alphaCSR[ 153 ][ 333 ],
   alphaCSR[ 153 ][ 334 ],
   alphaCSR[ 153 ][ 335 ],
   alphaCSR[ 153 ][ 336 ],
   alphaCSR[ 153 ][ 337 ],
   alphaCSR[ 153 ][ 338 ],
   alphaCSR[ 153 ][ 339 ],
   alphaCSR[ 153 ][ 340 ],
   alphaCSR[ 153 ][ 341 ],
   alphaCSR[ 153 ][ 342 ],
   alphaCSR[ 153 ][ 343 ],
   alphaCSR[ 153 ][ 344 ],
   alphaCSR[ 153 ][ 345 ],
   alphaCSR[ 153 ][ 346 ],
   alphaCSR[ 153 ][ 347 ],
   alphaCSR[ 153 ][ 348 ],
   alphaCSR[ 153 ][ 349 ],
   alphaCSR[ 153 ][ 350 ],
   alphaCSR[ 153 ][ 351 ],
   alphaCSR[ 153 ][ 352 ],
   alphaCSR[ 153 ][ 353 ],
   alphaCSR[ 153 ][ 354 ],
   alphaCSR[ 153 ][ 355 ],
   alphaCSR[ 153 ][ 356 ],
   alphaCSR[ 153 ][ 357 ],
   alphaCSR[ 153 ][ 358 ],
   alphaCSR[ 153 ][ 359 ],
   alphaCSR[ 153 ][ 360 ],
   alphaCSR[ 153 ][ 361 ],
   alphaCSR[ 153 ][ 362 ],
   alphaCSR[ 153 ][ 363 ],
   alphaCSR[ 153 ][ 364 ],
   alphaCSR[ 153 ][ 365 ],
   alphaCSR[ 153 ][ 366 ],
   alphaCSR[ 153 ][ 367 ],
   alphaCSR[ 153 ][ 368 ],
   alphaCSR[ 153 ][ 369 ],
   alphaCSR[ 153 ][ 370 ],
   alphaCSR[ 153 ][ 371 ],
   alphaCSR[ 153 ][ 372 ],
   alphaCSR[ 153 ][ 373 ],
   alphaCSR[ 153 ][ 374 ],
   alphaCSR[ 153 ][ 375 ],
   alphaCSR[ 153 ][ 376 ],
   alphaCSR[ 153 ][ 377 ],
   alphaCSR[ 153 ][ 378 ],
   alphaCSR[ 153 ][ 379 ],
   alphaCSR[ 153 ][ 380 ],
   alphaCSR[ 153 ][ 381 ],
   alphaCSR[ 153 ][ 382 ],
   alphaCSR[ 153 ][ 383 ],
   alphaCSR[ 154 ][ 0 ],
   alphaCSR[ 154 ][ 1 ],
   alphaCSR[ 154 ][ 2 ],
   alphaCSR[ 154 ][ 3 ],
   alphaCSR[ 154 ][ 4 ],
   alphaCSR[ 154 ][ 5 ],
   alphaCSR[ 154 ][ 6 ],
   alphaCSR[ 154 ][ 7 ],
   alphaCSR[ 154 ][ 8 ],
   alphaCSR[ 154 ][ 9 ],
   alphaCSR[ 154 ][ 10 ],
   alphaCSR[ 154 ][ 11 ],
   alphaCSR[ 154 ][ 12 ],
   alphaCSR[ 154 ][ 13 ],
   alphaCSR[ 154 ][ 14 ],
   alphaCSR[ 154 ][ 15 ],
   alphaCSR[ 154 ][ 16 ],
   alphaCSR[ 154 ][ 17 ],
   alphaCSR[ 154 ][ 18 ],
   alphaCSR[ 154 ][ 19 ],
   alphaCSR[ 154 ][ 20 ],
   alphaCSR[ 154 ][ 21 ],
   alphaCSR[ 154 ][ 22 ],
   alphaCSR[ 154 ][ 23 ],
   alphaCSR[ 154 ][ 24 ],
   alphaCSR[ 154 ][ 25 ],
   alphaCSR[ 154 ][ 26 ],
   alphaCSR[ 154 ][ 27 ],
   alphaCSR[ 154 ][ 28 ],
   alphaCSR[ 154 ][ 29 ],
   alphaCSR[ 154 ][ 30 ],
   alphaCSR[ 154 ][ 31 ],
   alphaCSR[ 154 ][ 32 ],
   alphaCSR[ 154 ][ 33 ],
   alphaCSR[ 154 ][ 34 ],
   alphaCSR[ 154 ][ 35 ],
   alphaCSR[ 154 ][ 36 ],
   alphaCSR[ 154 ][ 37 ],
   alphaCSR[ 154 ][ 38 ],
   alphaCSR[ 154 ][ 39 ],
   alphaCSR[ 154 ][ 40 ],
   alphaCSR[ 154 ][ 41 ],
   alphaCSR[ 154 ][ 42 ],
   alphaCSR[ 154 ][ 43 ],
   alphaCSR[ 154 ][ 44 ],
   alphaCSR[ 154 ][ 45 ],
   alphaCSR[ 154 ][ 46 ],
   alphaCSR[ 154 ][ 47 ],
   alphaCSR[ 154 ][ 48 ],
   alphaCSR[ 154 ][ 49 ],
   alphaCSR[ 154 ][ 50 ],
   alphaCSR[ 154 ][ 51 ],
   alphaCSR[ 154 ][ 52 ],
   alphaCSR[ 154 ][ 53 ],
   alphaCSR[ 154 ][ 54 ],
   alphaCSR[ 154 ][ 55 ],
   alphaCSR[ 154 ][ 56 ],
   alphaCSR[ 154 ][ 57 ],
   alphaCSR[ 154 ][ 58 ],
   alphaCSR[ 154 ][ 59 ],
   alphaCSR[ 154 ][ 60 ],
   alphaCSR[ 154 ][ 61 ],
   alphaCSR[ 154 ][ 62 ],
   alphaCSR[ 154 ][ 63 ],
   alphaCSR[ 154 ][ 64 ],
   alphaCSR[ 154 ][ 65 ],
   alphaCSR[ 154 ][ 66 ],
   alphaCSR[ 154 ][ 67 ],
   alphaCSR[ 154 ][ 68 ],
   alphaCSR[ 154 ][ 69 ],
   alphaCSR[ 154 ][ 70 ],
   alphaCSR[ 154 ][ 71 ],
   alphaCSR[ 154 ][ 72 ],
   alphaCSR[ 154 ][ 73 ],
   alphaCSR[ 154 ][ 74 ],
   alphaCSR[ 154 ][ 75 ],
   alphaCSR[ 154 ][ 76 ],
   alphaCSR[ 154 ][ 77 ],
   alphaCSR[ 154 ][ 78 ],
   alphaCSR[ 154 ][ 79 ],
   alphaCSR[ 154 ][ 80 ],
   alphaCSR[ 154 ][ 81 ],
   alphaCSR[ 154 ][ 82 ],
   alphaCSR[ 154 ][ 83 ],
   alphaCSR[ 154 ][ 84 ],
   alphaCSR[ 154 ][ 85 ],
   alphaCSR[ 154 ][ 86 ],
   alphaCSR[ 154 ][ 87 ],
   alphaCSR[ 154 ][ 88 ],
   alphaCSR[ 154 ][ 89 ],
   alphaCSR[ 154 ][ 90 ],
   alphaCSR[ 154 ][ 91 ],
   alphaCSR[ 154 ][ 92 ],
   alphaCSR[ 154 ][ 93 ],
   alphaCSR[ 154 ][ 94 ],
   alphaCSR[ 154 ][ 95 ],
   alphaCSR[ 154 ][ 96 ],
   alphaCSR[ 154 ][ 97 ],
   alphaCSR[ 154 ][ 98 ],
   alphaCSR[ 154 ][ 99 ],
   alphaCSR[ 154 ][ 100 ],
   alphaCSR[ 154 ][ 101 ],
   alphaCSR[ 154 ][ 102 ],
   alphaCSR[ 154 ][ 103 ],
   alphaCSR[ 154 ][ 104 ],
   alphaCSR[ 154 ][ 105 ],
   alphaCSR[ 154 ][ 106 ],
   alphaCSR[ 154 ][ 107 ],
   alphaCSR[ 154 ][ 108 ],
   alphaCSR[ 154 ][ 109 ],
   alphaCSR[ 154 ][ 110 ],
   alphaCSR[ 154 ][ 111 ],
   alphaCSR[ 154 ][ 112 ],
   alphaCSR[ 154 ][ 113 ],
   alphaCSR[ 154 ][ 114 ],
   alphaCSR[ 154 ][ 115 ],
   alphaCSR[ 154 ][ 116 ],
   alphaCSR[ 154 ][ 117 ],
   alphaCSR[ 154 ][ 118 ],
   alphaCSR[ 154 ][ 119 ],
   alphaCSR[ 154 ][ 120 ],
   alphaCSR[ 154 ][ 121 ],
   alphaCSR[ 154 ][ 122 ],
   alphaCSR[ 154 ][ 123 ],
   alphaCSR[ 154 ][ 124 ],
   alphaCSR[ 154 ][ 125 ],
   alphaCSR[ 154 ][ 126 ],
   alphaCSR[ 154 ][ 127 ],
   alphaCSR[ 154 ][ 128 ],
   alphaCSR[ 154 ][ 129 ],
   alphaCSR[ 154 ][ 130 ],
   alphaCSR[ 154 ][ 131 ],
   alphaCSR[ 154 ][ 132 ],
   alphaCSR[ 154 ][ 133 ],
   alphaCSR[ 154 ][ 134 ],
   alphaCSR[ 154 ][ 135 ],
   alphaCSR[ 154 ][ 136 ],
   alphaCSR[ 154 ][ 137 ],
   alphaCSR[ 154 ][ 138 ],
   alphaCSR[ 154 ][ 139 ],
   alphaCSR[ 154 ][ 140 ],
   alphaCSR[ 154 ][ 141 ],
   alphaCSR[ 154 ][ 142 ],
   alphaCSR[ 154 ][ 143 ],
   alphaCSR[ 154 ][ 144 ],
   alphaCSR[ 154 ][ 145 ],
   alphaCSR[ 154 ][ 146 ],
   alphaCSR[ 154 ][ 147 ],
   alphaCSR[ 154 ][ 148 ],
   alphaCSR[ 154 ][ 149 ],
   alphaCSR[ 154 ][ 150 ],
   alphaCSR[ 154 ][ 151 ],
   alphaCSR[ 154 ][ 152 ],
   alphaCSR[ 154 ][ 153 ],
   alphaCSR[ 154 ][ 154 ],
   alphaCSR[ 154 ][ 155 ],
   alphaCSR[ 154 ][ 156 ],
   alphaCSR[ 154 ][ 157 ],
   alphaCSR[ 154 ][ 158 ],
   alphaCSR[ 154 ][ 159 ],
   alphaCSR[ 154 ][ 160 ],
   alphaCSR[ 154 ][ 161 ],
   alphaCSR[ 154 ][ 162 ],
   alphaCSR[ 154 ][ 163 ],
   alphaCSR[ 154 ][ 164 ],
   alphaCSR[ 154 ][ 165 ],
   alphaCSR[ 154 ][ 166 ],
   alphaCSR[ 154 ][ 167 ],
   alphaCSR[ 154 ][ 168 ],
   alphaCSR[ 154 ][ 169 ],
   alphaCSR[ 154 ][ 170 ],
   alphaCSR[ 154 ][ 171 ],
   alphaCSR[ 154 ][ 172 ],
   alphaCSR[ 154 ][ 173 ],
   alphaCSR[ 154 ][ 174 ],
   alphaCSR[ 154 ][ 175 ],
   alphaCSR[ 154 ][ 176 ],
   alphaCSR[ 154 ][ 177 ],
   alphaCSR[ 154 ][ 178 ],
   alphaCSR[ 154 ][ 179 ],
   alphaCSR[ 154 ][ 180 ],
   alphaCSR[ 154 ][ 181 ],
   alphaCSR[ 154 ][ 182 ],
   alphaCSR[ 154 ][ 183 ],
   alphaCSR[ 154 ][ 184 ],
   alphaCSR[ 154 ][ 185 ],
   alphaCSR[ 154 ][ 186 ],
   alphaCSR[ 154 ][ 187 ],
   alphaCSR[ 154 ][ 188 ],
   alphaCSR[ 154 ][ 189 ],
   alphaCSR[ 154 ][ 190 ],
   alphaCSR[ 154 ][ 191 ],
   alphaCSR[ 154 ][ 192 ],
   alphaCSR[ 154 ][ 193 ],
   alphaCSR[ 154 ][ 194 ],
   alphaCSR[ 154 ][ 195 ],
   alphaCSR[ 154 ][ 196 ],
   alphaCSR[ 154 ][ 197 ],
   alphaCSR[ 154 ][ 198 ],
   alphaCSR[ 154 ][ 199 ],
   alphaCSR[ 154 ][ 200 ],
   alphaCSR[ 154 ][ 201 ],
   alphaCSR[ 154 ][ 202 ],
   alphaCSR[ 154 ][ 203 ],
   alphaCSR[ 154 ][ 204 ],
   alphaCSR[ 154 ][ 205 ],
   alphaCSR[ 154 ][ 206 ],
   alphaCSR[ 154 ][ 207 ],
   alphaCSR[ 154 ][ 208 ],
   alphaCSR[ 154 ][ 209 ],
   alphaCSR[ 154 ][ 210 ],
   alphaCSR[ 154 ][ 211 ],
   alphaCSR[ 154 ][ 212 ],
   alphaCSR[ 154 ][ 213 ],
   alphaCSR[ 154 ][ 214 ],
   alphaCSR[ 154 ][ 215 ],
   alphaCSR[ 154 ][ 216 ],
   alphaCSR[ 154 ][ 217 ],
   alphaCSR[ 154 ][ 218 ],
   alphaCSR[ 154 ][ 219 ],
   alphaCSR[ 154 ][ 220 ],
   alphaCSR[ 154 ][ 221 ],
   alphaCSR[ 154 ][ 222 ],
   alphaCSR[ 154 ][ 223 ],
   alphaCSR[ 154 ][ 224 ],
   alphaCSR[ 154 ][ 225 ],
   alphaCSR[ 154 ][ 226 ],
   alphaCSR[ 154 ][ 227 ],
   alphaCSR[ 154 ][ 228 ],
   alphaCSR[ 154 ][ 229 ],
   alphaCSR[ 154 ][ 230 ],
   alphaCSR[ 154 ][ 231 ],
   alphaCSR[ 154 ][ 232 ],
   alphaCSR[ 154 ][ 233 ],
   alphaCSR[ 154 ][ 234 ],
   alphaCSR[ 154 ][ 235 ],
   alphaCSR[ 154 ][ 236 ],
   alphaCSR[ 154 ][ 237 ],
   alphaCSR[ 154 ][ 238 ],
   alphaCSR[ 154 ][ 239 ],
   alphaCSR[ 154 ][ 240 ],
   alphaCSR[ 154 ][ 241 ],
   alphaCSR[ 154 ][ 242 ],
   alphaCSR[ 154 ][ 243 ],
   alphaCSR[ 154 ][ 244 ],
   alphaCSR[ 154 ][ 245 ],
   alphaCSR[ 154 ][ 246 ],
   alphaCSR[ 154 ][ 247 ],
   alphaCSR[ 154 ][ 248 ],
   alphaCSR[ 154 ][ 249 ],
   alphaCSR[ 154 ][ 250 ],
   alphaCSR[ 154 ][ 251 ],
   alphaCSR[ 154 ][ 252 ],
   alphaCSR[ 154 ][ 253 ],
   alphaCSR[ 154 ][ 254 ],
   alphaCSR[ 154 ][ 255 ],
   alphaCSR[ 154 ][ 256 ],
   alphaCSR[ 154 ][ 257 ],
   alphaCSR[ 154 ][ 258 ],
   alphaCSR[ 154 ][ 259 ],
   alphaCSR[ 154 ][ 260 ],
   alphaCSR[ 154 ][ 261 ],
   alphaCSR[ 154 ][ 262 ],
   alphaCSR[ 154 ][ 263 ],
   alphaCSR[ 154 ][ 264 ],
   alphaCSR[ 154 ][ 265 ],
   alphaCSR[ 154 ][ 266 ],
   alphaCSR[ 154 ][ 267 ],
   alphaCSR[ 154 ][ 268 ],
   alphaCSR[ 154 ][ 269 ],
   alphaCSR[ 154 ][ 270 ],
   alphaCSR[ 154 ][ 271 ],
   alphaCSR[ 154 ][ 272 ],
   alphaCSR[ 154 ][ 273 ],
   alphaCSR[ 154 ][ 274 ],
   alphaCSR[ 154 ][ 275 ],
   alphaCSR[ 154 ][ 276 ],
   alphaCSR[ 154 ][ 277 ],
   alphaCSR[ 154 ][ 278 ],
   alphaCSR[ 154 ][ 279 ],
   alphaCSR[ 154 ][ 280 ],
   alphaCSR[ 154 ][ 281 ],
   alphaCSR[ 154 ][ 282 ],
   alphaCSR[ 154 ][ 283 ],
   alphaCSR[ 154 ][ 284 ],
   alphaCSR[ 154 ][ 285 ],
   alphaCSR[ 154 ][ 286 ],
   alphaCSR[ 154 ][ 287 ],
   alphaCSR[ 154 ][ 288 ],
   alphaCSR[ 154 ][ 289 ],
   alphaCSR[ 154 ][ 290 ],
   alphaCSR[ 154 ][ 291 ],
   alphaCSR[ 154 ][ 292 ],
   alphaCSR[ 154 ][ 293 ],
   alphaCSR[ 154 ][ 294 ],
   alphaCSR[ 154 ][ 295 ],
   alphaCSR[ 154 ][ 296 ],
   alphaCSR[ 154 ][ 297 ],
   alphaCSR[ 154 ][ 298 ],
   alphaCSR[ 154 ][ 299 ],
   alphaCSR[ 154 ][ 300 ],
   alphaCSR[ 154 ][ 301 ],
   alphaCSR[ 154 ][ 302 ],
   alphaCSR[ 154 ][ 303 ],
   alphaCSR[ 154 ][ 304 ],
   alphaCSR[ 154 ][ 305 ],
   alphaCSR[ 154 ][ 306 ],
   alphaCSR[ 154 ][ 307 ],
   alphaCSR[ 154 ][ 308 ],
   alphaCSR[ 154 ][ 309 ],
   alphaCSR[ 154 ][ 310 ],
   alphaCSR[ 154 ][ 311 ],
   alphaCSR[ 154 ][ 312 ],
   alphaCSR[ 154 ][ 313 ],
   alphaCSR[ 154 ][ 314 ],
   alphaCSR[ 154 ][ 315 ],
   alphaCSR[ 154 ][ 316 ],
   alphaCSR[ 154 ][ 317 ],
   alphaCSR[ 154 ][ 318 ],
   alphaCSR[ 154 ][ 319 ],
   alphaCSR[ 154 ][ 320 ],
   alphaCSR[ 154 ][ 321 ],
   alphaCSR[ 154 ][ 322 ],
   alphaCSR[ 154 ][ 323 ],
   alphaCSR[ 154 ][ 324 ],
   alphaCSR[ 154 ][ 325 ],
   alphaCSR[ 154 ][ 326 ],
   alphaCSR[ 154 ][ 327 ],
   alphaCSR[ 154 ][ 328 ],
   alphaCSR[ 154 ][ 329 ],
   alphaCSR[ 154 ][ 330 ],
   alphaCSR[ 154 ][ 331 ],
   alphaCSR[ 154 ][ 332 ],
   alphaCSR[ 154 ][ 333 ],
   alphaCSR[ 154 ][ 334 ],
   alphaCSR[ 154 ][ 335 ],
   alphaCSR[ 154 ][ 336 ],
   alphaCSR[ 154 ][ 337 ],
   alphaCSR[ 154 ][ 338 ],
   alphaCSR[ 154 ][ 339 ],
   alphaCSR[ 154 ][ 340 ],
   alphaCSR[ 154 ][ 341 ],
   alphaCSR[ 154 ][ 342 ],
   alphaCSR[ 154 ][ 343 ],
   alphaCSR[ 154 ][ 344 ],
   alphaCSR[ 154 ][ 345 ],
   alphaCSR[ 154 ][ 346 ],
   alphaCSR[ 154 ][ 347 ],
   alphaCSR[ 154 ][ 348 ],
   alphaCSR[ 154 ][ 349 ],
   alphaCSR[ 154 ][ 350 ],
   alphaCSR[ 154 ][ 351 ],
   alphaCSR[ 154 ][ 352 ],
   alphaCSR[ 154 ][ 353 ],
   alphaCSR[ 154 ][ 354 ],
   alphaCSR[ 154 ][ 355 ],
   alphaCSR[ 154 ][ 356 ],
   alphaCSR[ 154 ][ 357 ],
   alphaCSR[ 154 ][ 358 ],
   alphaCSR[ 154 ][ 359 ],
   alphaCSR[ 154 ][ 360 ],
   alphaCSR[ 154 ][ 361 ],
   alphaCSR[ 154 ][ 362 ],
   alphaCSR[ 154 ][ 363 ],
   alphaCSR[ 154 ][ 364 ],
   alphaCSR[ 154 ][ 365 ],
   alphaCSR[ 154 ][ 366 ],
   alphaCSR[ 154 ][ 367 ],
   alphaCSR[ 154 ][ 368 ],
   alphaCSR[ 154 ][ 369 ],
   alphaCSR[ 154 ][ 370 ],
   alphaCSR[ 154 ][ 371 ],
   alphaCSR[ 154 ][ 372 ],
   alphaCSR[ 154 ][ 373 ],
   alphaCSR[ 154 ][ 374 ],
   alphaCSR[ 154 ][ 375 ],
   alphaCSR[ 154 ][ 376 ],
   alphaCSR[ 154 ][ 377 ],
   alphaCSR[ 154 ][ 378 ],
   alphaCSR[ 154 ][ 379 ],
   alphaCSR[ 154 ][ 380 ],
   alphaCSR[ 154 ][ 381 ],
   alphaCSR[ 154 ][ 382 ],
   alphaCSR[ 154 ][ 383 ],
   alphaCSR[ 155 ][ 0 ],
   alphaCSR[ 155 ][ 1 ],
   alphaCSR[ 155 ][ 2 ],
   alphaCSR[ 155 ][ 3 ],
   alphaCSR[ 155 ][ 4 ],
   alphaCSR[ 155 ][ 5 ],
   alphaCSR[ 155 ][ 6 ],
   alphaCSR[ 155 ][ 7 ],
   alphaCSR[ 155 ][ 8 ],
   alphaCSR[ 155 ][ 9 ],
   alphaCSR[ 155 ][ 10 ],
   alphaCSR[ 155 ][ 11 ],
   alphaCSR[ 155 ][ 12 ],
   alphaCSR[ 155 ][ 13 ],
   alphaCSR[ 155 ][ 14 ],
   alphaCSR[ 155 ][ 15 ],
   alphaCSR[ 155 ][ 16 ],
   alphaCSR[ 155 ][ 17 ],
   alphaCSR[ 155 ][ 18 ],
   alphaCSR[ 155 ][ 19 ],
   alphaCSR[ 155 ][ 20 ],
   alphaCSR[ 155 ][ 21 ],
   alphaCSR[ 155 ][ 22 ],
   alphaCSR[ 155 ][ 23 ],
   alphaCSR[ 155 ][ 24 ],
   alphaCSR[ 155 ][ 25 ],
   alphaCSR[ 155 ][ 26 ],
   alphaCSR[ 155 ][ 27 ],
   alphaCSR[ 155 ][ 28 ],
   alphaCSR[ 155 ][ 29 ],
   alphaCSR[ 155 ][ 30 ],
   alphaCSR[ 155 ][ 31 ],
   alphaCSR[ 155 ][ 32 ],
   alphaCSR[ 155 ][ 33 ],
   alphaCSR[ 155 ][ 34 ],
   alphaCSR[ 155 ][ 35 ],
   alphaCSR[ 155 ][ 36 ],
   alphaCSR[ 155 ][ 37 ],
   alphaCSR[ 155 ][ 38 ],
   alphaCSR[ 155 ][ 39 ],
   alphaCSR[ 155 ][ 40 ],
   alphaCSR[ 155 ][ 41 ],
   alphaCSR[ 155 ][ 42 ],
   alphaCSR[ 155 ][ 43 ],
   alphaCSR[ 155 ][ 44 ],
   alphaCSR[ 155 ][ 45 ],
   alphaCSR[ 155 ][ 46 ],
   alphaCSR[ 155 ][ 47 ],
   alphaCSR[ 155 ][ 48 ],
   alphaCSR[ 155 ][ 49 ],
   alphaCSR[ 155 ][ 50 ],
   alphaCSR[ 155 ][ 51 ],
   alphaCSR[ 155 ][ 52 ],
   alphaCSR[ 155 ][ 53 ],
   alphaCSR[ 155 ][ 54 ],
   alphaCSR[ 155 ][ 55 ],
   alphaCSR[ 155 ][ 56 ],
   alphaCSR[ 155 ][ 57 ],
   alphaCSR[ 155 ][ 58 ],
   alphaCSR[ 155 ][ 59 ],
   alphaCSR[ 155 ][ 60 ],
   alphaCSR[ 155 ][ 61 ],
   alphaCSR[ 155 ][ 62 ],
   alphaCSR[ 155 ][ 63 ],
   alphaCSR[ 155 ][ 64 ],
   alphaCSR[ 155 ][ 65 ],
   alphaCSR[ 155 ][ 66 ],
   alphaCSR[ 155 ][ 67 ],
   alphaCSR[ 155 ][ 68 ],
   alphaCSR[ 155 ][ 69 ],
   alphaCSR[ 155 ][ 70 ],
   alphaCSR[ 155 ][ 71 ],
   alphaCSR[ 155 ][ 72 ],
   alphaCSR[ 155 ][ 73 ],
   alphaCSR[ 155 ][ 74 ],
   alphaCSR[ 155 ][ 75 ],
   alphaCSR[ 155 ][ 76 ],
   alphaCSR[ 155 ][ 77 ],
   alphaCSR[ 155 ][ 78 ],
   alphaCSR[ 155 ][ 79 ],
   alphaCSR[ 155 ][ 80 ],
   alphaCSR[ 155 ][ 81 ],
   alphaCSR[ 155 ][ 82 ],
   alphaCSR[ 155 ][ 83 ],
   alphaCSR[ 155 ][ 84 ],
   alphaCSR[ 155 ][ 85 ],
   alphaCSR[ 155 ][ 86 ],
   alphaCSR[ 155 ][ 87 ],
   alphaCSR[ 155 ][ 88 ],
   alphaCSR[ 155 ][ 89 ],
   alphaCSR[ 155 ][ 90 ],
   alphaCSR[ 155 ][ 91 ],
   alphaCSR[ 155 ][ 92 ],
   alphaCSR[ 155 ][ 93 ],
   alphaCSR[ 155 ][ 94 ],
   alphaCSR[ 155 ][ 95 ],
   alphaCSR[ 155 ][ 96 ],
   alphaCSR[ 155 ][ 97 ],
   alphaCSR[ 155 ][ 98 ],
   alphaCSR[ 155 ][ 99 ],
   alphaCSR[ 155 ][ 100 ],
   alphaCSR[ 155 ][ 101 ],
   alphaCSR[ 155 ][ 102 ],
   alphaCSR[ 155 ][ 103 ],
   alphaCSR[ 155 ][ 104 ],
   alphaCSR[ 155 ][ 105 ],
   alphaCSR[ 155 ][ 106 ],
   alphaCSR[ 155 ][ 107 ],
   alphaCSR[ 155 ][ 108 ],
   alphaCSR[ 155 ][ 109 ],
   alphaCSR[ 155 ][ 110 ],
   alphaCSR[ 155 ][ 111 ],
   alphaCSR[ 155 ][ 112 ],
   alphaCSR[ 155 ][ 113 ],
   alphaCSR[ 155 ][ 114 ],
   alphaCSR[ 155 ][ 115 ],
   alphaCSR[ 155 ][ 116 ],
   alphaCSR[ 155 ][ 117 ],
   alphaCSR[ 155 ][ 118 ],
   alphaCSR[ 155 ][ 119 ],
   alphaCSR[ 155 ][ 120 ],
   alphaCSR[ 155 ][ 121 ],
   alphaCSR[ 155 ][ 122 ],
   alphaCSR[ 155 ][ 123 ],
   alphaCSR[ 155 ][ 124 ],
   alphaCSR[ 155 ][ 125 ],
   alphaCSR[ 155 ][ 126 ],
   alphaCSR[ 155 ][ 127 ],
   alphaCSR[ 155 ][ 128 ],
   alphaCSR[ 155 ][ 129 ],
   alphaCSR[ 155 ][ 130 ],
   alphaCSR[ 155 ][ 131 ],
   alphaCSR[ 155 ][ 132 ],
   alphaCSR[ 155 ][ 133 ],
   alphaCSR[ 155 ][ 134 ],
   alphaCSR[ 155 ][ 135 ],
   alphaCSR[ 155 ][ 136 ],
   alphaCSR[ 155 ][ 137 ],
   alphaCSR[ 155 ][ 138 ],
   alphaCSR[ 155 ][ 139 ],
   alphaCSR[ 155 ][ 140 ],
   alphaCSR[ 155 ][ 141 ],
   alphaCSR[ 155 ][ 142 ],
   alphaCSR[ 155 ][ 143 ],
   alphaCSR[ 155 ][ 144 ],
   alphaCSR[ 155 ][ 145 ],
   alphaCSR[ 155 ][ 146 ],
   alphaCSR[ 155 ][ 147 ],
   alphaCSR[ 155 ][ 148 ],
   alphaCSR[ 155 ][ 149 ],
   alphaCSR[ 155 ][ 150 ],
   alphaCSR[ 155 ][ 151 ],
   alphaCSR[ 155 ][ 152 ],
   alphaCSR[ 155 ][ 153 ],
   alphaCSR[ 155 ][ 154 ],
   alphaCSR[ 155 ][ 155 ],
   alphaCSR[ 155 ][ 156 ],
   alphaCSR[ 155 ][ 157 ],
   alphaCSR[ 155 ][ 158 ],
   alphaCSR[ 155 ][ 159 ],
   alphaCSR[ 155 ][ 160 ],
   alphaCSR[ 155 ][ 161 ],
   alphaCSR[ 155 ][ 162 ],
   alphaCSR[ 155 ][ 163 ],
   alphaCSR[ 155 ][ 164 ],
   alphaCSR[ 155 ][ 165 ],
   alphaCSR[ 155 ][ 166 ],
   alphaCSR[ 155 ][ 167 ],
   alphaCSR[ 155 ][ 168 ],
   alphaCSR[ 155 ][ 169 ],
   alphaCSR[ 155 ][ 170 ],
   alphaCSR[ 155 ][ 171 ],
   alphaCSR[ 155 ][ 172 ],
   alphaCSR[ 155 ][ 173 ],
   alphaCSR[ 155 ][ 174 ],
   alphaCSR[ 155 ][ 175 ],
   alphaCSR[ 155 ][ 176 ],
   alphaCSR[ 155 ][ 177 ],
   alphaCSR[ 155 ][ 178 ],
   alphaCSR[ 155 ][ 179 ],
   alphaCSR[ 155 ][ 180 ],
   alphaCSR[ 155 ][ 181 ],
   alphaCSR[ 155 ][ 182 ],
   alphaCSR[ 155 ][ 183 ],
   alphaCSR[ 155 ][ 184 ],
   alphaCSR[ 155 ][ 185 ],
   alphaCSR[ 155 ][ 186 ],
   alphaCSR[ 155 ][ 187 ],
   alphaCSR[ 155 ][ 188 ],
   alphaCSR[ 155 ][ 189 ],
   alphaCSR[ 155 ][ 190 ],
   alphaCSR[ 155 ][ 191 ],
   alphaCSR[ 155 ][ 192 ],
   alphaCSR[ 155 ][ 193 ],
   alphaCSR[ 155 ][ 194 ],
   alphaCSR[ 155 ][ 195 ],
   alphaCSR[ 155 ][ 196 ],
   alphaCSR[ 155 ][ 197 ],
   alphaCSR[ 155 ][ 198 ],
   alphaCSR[ 155 ][ 199 ],
   alphaCSR[ 155 ][ 200 ],
   alphaCSR[ 155 ][ 201 ],
   alphaCSR[ 155 ][ 202 ],
   alphaCSR[ 155 ][ 203 ],
   alphaCSR[ 155 ][ 204 ],
   alphaCSR[ 155 ][ 205 ],
   alphaCSR[ 155 ][ 206 ],
   alphaCSR[ 155 ][ 207 ],
   alphaCSR[ 155 ][ 208 ],
   alphaCSR[ 155 ][ 209 ],
   alphaCSR[ 155 ][ 210 ],
   alphaCSR[ 155 ][ 211 ],
   alphaCSR[ 155 ][ 212 ],
   alphaCSR[ 155 ][ 213 ],
   alphaCSR[ 155 ][ 214 ],
   alphaCSR[ 155 ][ 215 ],
   alphaCSR[ 155 ][ 216 ],
   alphaCSR[ 155 ][ 217 ],
   alphaCSR[ 155 ][ 218 ],
   alphaCSR[ 155 ][ 219 ],
   alphaCSR[ 155 ][ 220 ],
   alphaCSR[ 155 ][ 221 ],
   alphaCSR[ 155 ][ 222 ],
   alphaCSR[ 155 ][ 223 ],
   alphaCSR[ 155 ][ 224 ],
   alphaCSR[ 155 ][ 225 ],
   alphaCSR[ 155 ][ 226 ],
   alphaCSR[ 155 ][ 227 ],
   alphaCSR[ 155 ][ 228 ],
   alphaCSR[ 155 ][ 229 ],
   alphaCSR[ 155 ][ 230 ],
   alphaCSR[ 155 ][ 231 ],
   alphaCSR[ 155 ][ 232 ],
   alphaCSR[ 155 ][ 233 ],
   alphaCSR[ 155 ][ 234 ],
   alphaCSR[ 155 ][ 235 ],
   alphaCSR[ 155 ][ 236 ],
   alphaCSR[ 155 ][ 237 ],
   alphaCSR[ 155 ][ 238 ],
   alphaCSR[ 155 ][ 239 ],
   alphaCSR[ 155 ][ 240 ],
   alphaCSR[ 155 ][ 241 ],
   alphaCSR[ 155 ][ 242 ],
   alphaCSR[ 155 ][ 243 ],
   alphaCSR[ 155 ][ 244 ],
   alphaCSR[ 155 ][ 245 ],
   alphaCSR[ 155 ][ 246 ],
   alphaCSR[ 155 ][ 247 ],
   alphaCSR[ 155 ][ 248 ],
   alphaCSR[ 155 ][ 249 ],
   alphaCSR[ 155 ][ 250 ],
   alphaCSR[ 155 ][ 251 ],
   alphaCSR[ 155 ][ 252 ],
   alphaCSR[ 155 ][ 253 ],
   alphaCSR[ 155 ][ 254 ],
   alphaCSR[ 155 ][ 255 ],
   alphaCSR[ 155 ][ 256 ],
   alphaCSR[ 155 ][ 257 ],
   alphaCSR[ 155 ][ 258 ],
   alphaCSR[ 155 ][ 259 ],
   alphaCSR[ 155 ][ 260 ],
   alphaCSR[ 155 ][ 261 ],
   alphaCSR[ 155 ][ 262 ],
   alphaCSR[ 155 ][ 263 ],
   alphaCSR[ 155 ][ 264 ],
   alphaCSR[ 155 ][ 265 ],
   alphaCSR[ 155 ][ 266 ],
   alphaCSR[ 155 ][ 267 ],
   alphaCSR[ 155 ][ 268 ],
   alphaCSR[ 155 ][ 269 ],
   alphaCSR[ 155 ][ 270 ],
   alphaCSR[ 155 ][ 271 ],
   alphaCSR[ 155 ][ 272 ],
   alphaCSR[ 155 ][ 273 ],
   alphaCSR[ 155 ][ 274 ],
   alphaCSR[ 155 ][ 275 ],
   alphaCSR[ 155 ][ 276 ],
   alphaCSR[ 155 ][ 277 ],
   alphaCSR[ 155 ][ 278 ],
   alphaCSR[ 155 ][ 279 ],
   alphaCSR[ 155 ][ 280 ],
   alphaCSR[ 155 ][ 281 ],
   alphaCSR[ 155 ][ 282 ],
   alphaCSR[ 155 ][ 283 ],
   alphaCSR[ 155 ][ 284 ],
   alphaCSR[ 155 ][ 285 ],
   alphaCSR[ 155 ][ 286 ],
   alphaCSR[ 155 ][ 287 ],
   alphaCSR[ 155 ][ 288 ],
   alphaCSR[ 155 ][ 289 ],
   alphaCSR[ 155 ][ 290 ],
   alphaCSR[ 155 ][ 291 ],
   alphaCSR[ 155 ][ 292 ],
   alphaCSR[ 155 ][ 293 ],
   alphaCSR[ 155 ][ 294 ],
   alphaCSR[ 155 ][ 295 ],
   alphaCSR[ 155 ][ 296 ],
   alphaCSR[ 155 ][ 297 ],
   alphaCSR[ 155 ][ 298 ],
   alphaCSR[ 155 ][ 299 ],
   alphaCSR[ 155 ][ 300 ],
   alphaCSR[ 155 ][ 301 ],
   alphaCSR[ 155 ][ 302 ],
   alphaCSR[ 155 ][ 303 ],
   alphaCSR[ 155 ][ 304 ],
   alphaCSR[ 155 ][ 305 ],
   alphaCSR[ 155 ][ 306 ],
   alphaCSR[ 155 ][ 307 ],
   alphaCSR[ 155 ][ 308 ],
   alphaCSR[ 155 ][ 309 ],
   alphaCSR[ 155 ][ 310 ],
   alphaCSR[ 155 ][ 311 ],
   alphaCSR[ 155 ][ 312 ],
   alphaCSR[ 155 ][ 313 ],
   alphaCSR[ 155 ][ 314 ],
   alphaCSR[ 155 ][ 315 ],
   alphaCSR[ 155 ][ 316 ],
   alphaCSR[ 155 ][ 317 ],
   alphaCSR[ 155 ][ 318 ],
   alphaCSR[ 155 ][ 319 ],
   alphaCSR[ 155 ][ 320 ],
   alphaCSR[ 155 ][ 321 ],
   alphaCSR[ 155 ][ 322 ],
   alphaCSR[ 155 ][ 323 ],
   alphaCSR[ 155 ][ 324 ],
   alphaCSR[ 155 ][ 325 ],
   alphaCSR[ 155 ][ 326 ],
   alphaCSR[ 155 ][ 327 ],
   alphaCSR[ 155 ][ 328 ],
   alphaCSR[ 155 ][ 329 ],
   alphaCSR[ 155 ][ 330 ],
   alphaCSR[ 155 ][ 331 ],
   alphaCSR[ 155 ][ 332 ],
   alphaCSR[ 155 ][ 333 ],
   alphaCSR[ 155 ][ 334 ],
   alphaCSR[ 155 ][ 335 ],
   alphaCSR[ 155 ][ 336 ],
   alphaCSR[ 155 ][ 337 ],
   alphaCSR[ 155 ][ 338 ],
   alphaCSR[ 155 ][ 339 ],
   alphaCSR[ 155 ][ 340 ],
   alphaCSR[ 155 ][ 341 ],
   alphaCSR[ 155 ][ 342 ],
   alphaCSR[ 155 ][ 343 ],
   alphaCSR[ 155 ][ 344 ],
   alphaCSR[ 155 ][ 345 ],
   alphaCSR[ 155 ][ 346 ],
   alphaCSR[ 155 ][ 347 ],
   alphaCSR[ 155 ][ 348 ],
   alphaCSR[ 155 ][ 349 ],
   alphaCSR[ 155 ][ 350 ],
   alphaCSR[ 155 ][ 351 ],
   alphaCSR[ 155 ][ 352 ],
   alphaCSR[ 155 ][ 353 ],
   alphaCSR[ 155 ][ 354 ],
   alphaCSR[ 155 ][ 355 ],
   alphaCSR[ 155 ][ 356 ],
   alphaCSR[ 155 ][ 357 ],
   alphaCSR[ 155 ][ 358 ],
   alphaCSR[ 155 ][ 359 ],
   alphaCSR[ 155 ][ 360 ],
   alphaCSR[ 155 ][ 361 ],
   alphaCSR[ 155 ][ 362 ],
   alphaCSR[ 155 ][ 363 ],
   alphaCSR[ 155 ][ 364 ],
   alphaCSR[ 155 ][ 365 ],
   alphaCSR[ 155 ][ 366 ],
   alphaCSR[ 155 ][ 367 ],
   alphaCSR[ 155 ][ 368 ],
   alphaCSR[ 155 ][ 369 ],
   alphaCSR[ 155 ][ 370 ],
   alphaCSR[ 155 ][ 371 ],
   alphaCSR[ 155 ][ 372 ],
   alphaCSR[ 155 ][ 373 ],
   alphaCSR[ 155 ][ 374 ],
   alphaCSR[ 155 ][ 375 ],
   alphaCSR[ 155 ][ 376 ],
   alphaCSR[ 155 ][ 377 ],
   alphaCSR[ 155 ][ 378 ],
   alphaCSR[ 155 ][ 379 ],
   alphaCSR[ 155 ][ 380 ],
   alphaCSR[ 155 ][ 381 ],
   alphaCSR[ 155 ][ 382 ],
   alphaCSR[ 155 ][ 383 ],
   alphaCSR[ 156 ][ 0 ],
   alphaCSR[ 156 ][ 1 ],
   alphaCSR[ 156 ][ 2 ],
   alphaCSR[ 156 ][ 3 ],
   alphaCSR[ 156 ][ 4 ],
   alphaCSR[ 156 ][ 5 ],
   alphaCSR[ 156 ][ 6 ],
   alphaCSR[ 156 ][ 7 ],
   alphaCSR[ 156 ][ 8 ],
   alphaCSR[ 156 ][ 9 ],
   alphaCSR[ 156 ][ 10 ],
   alphaCSR[ 156 ][ 11 ],
   alphaCSR[ 156 ][ 12 ],
   alphaCSR[ 156 ][ 13 ],
   alphaCSR[ 156 ][ 14 ],
   alphaCSR[ 156 ][ 15 ],
   alphaCSR[ 156 ][ 16 ],
   alphaCSR[ 156 ][ 17 ],
   alphaCSR[ 156 ][ 18 ],
   alphaCSR[ 156 ][ 19 ],
   alphaCSR[ 156 ][ 20 ],
   alphaCSR[ 156 ][ 21 ],
   alphaCSR[ 156 ][ 22 ],
   alphaCSR[ 156 ][ 23 ],
   alphaCSR[ 156 ][ 24 ],
   alphaCSR[ 156 ][ 25 ],
   alphaCSR[ 156 ][ 26 ],
   alphaCSR[ 156 ][ 27 ],
   alphaCSR[ 156 ][ 28 ],
   alphaCSR[ 156 ][ 29 ],
   alphaCSR[ 156 ][ 30 ],
   alphaCSR[ 156 ][ 31 ],
   alphaCSR[ 156 ][ 32 ],
   alphaCSR[ 156 ][ 33 ],
   alphaCSR[ 156 ][ 34 ],
   alphaCSR[ 156 ][ 35 ],
   alphaCSR[ 156 ][ 36 ],
   alphaCSR[ 156 ][ 37 ],
   alphaCSR[ 156 ][ 38 ],
   alphaCSR[ 156 ][ 39 ],
   alphaCSR[ 156 ][ 40 ],
   alphaCSR[ 156 ][ 41 ],
   alphaCSR[ 156 ][ 42 ],
   alphaCSR[ 156 ][ 43 ],
   alphaCSR[ 156 ][ 44 ],
   alphaCSR[ 156 ][ 45 ],
   alphaCSR[ 156 ][ 46 ],
   alphaCSR[ 156 ][ 47 ],
   alphaCSR[ 156 ][ 48 ],
   alphaCSR[ 156 ][ 49 ],
   alphaCSR[ 156 ][ 50 ],
   alphaCSR[ 156 ][ 51 ],
   alphaCSR[ 156 ][ 52 ],
   alphaCSR[ 156 ][ 53 ],
   alphaCSR[ 156 ][ 54 ],
   alphaCSR[ 156 ][ 55 ],
   alphaCSR[ 156 ][ 56 ],
   alphaCSR[ 156 ][ 57 ],
   alphaCSR[ 156 ][ 58 ],
   alphaCSR[ 156 ][ 59 ],
   alphaCSR[ 156 ][ 60 ],
   alphaCSR[ 156 ][ 61 ],
   alphaCSR[ 156 ][ 62 ],
   alphaCSR[ 156 ][ 63 ],
   alphaCSR[ 156 ][ 64 ],
   alphaCSR[ 156 ][ 65 ],
   alphaCSR[ 156 ][ 66 ],
   alphaCSR[ 156 ][ 67 ],
   alphaCSR[ 156 ][ 68 ],
   alphaCSR[ 156 ][ 69 ],
   alphaCSR[ 156 ][ 70 ],
   alphaCSR[ 156 ][ 71 ],
   alphaCSR[ 156 ][ 72 ],
   alphaCSR[ 156 ][ 73 ],
   alphaCSR[ 156 ][ 74 ],
   alphaCSR[ 156 ][ 75 ],
   alphaCSR[ 156 ][ 76 ],
   alphaCSR[ 156 ][ 77 ],
   alphaCSR[ 156 ][ 78 ],
   alphaCSR[ 156 ][ 79 ],
   alphaCSR[ 156 ][ 80 ],
   alphaCSR[ 156 ][ 81 ],
   alphaCSR[ 156 ][ 82 ],
   alphaCSR[ 156 ][ 83 ],
   alphaCSR[ 156 ][ 84 ],
   alphaCSR[ 156 ][ 85 ],
   alphaCSR[ 156 ][ 86 ],
   alphaCSR[ 156 ][ 87 ],
   alphaCSR[ 156 ][ 88 ],
   alphaCSR[ 156 ][ 89 ],
   alphaCSR[ 156 ][ 90 ],
   alphaCSR[ 156 ][ 91 ],
   alphaCSR[ 156 ][ 92 ],
   alphaCSR[ 156 ][ 93 ],
   alphaCSR[ 156 ][ 94 ],
   alphaCSR[ 156 ][ 95 ],
   alphaCSR[ 156 ][ 96 ],
   alphaCSR[ 156 ][ 97 ],
   alphaCSR[ 156 ][ 98 ],
   alphaCSR[ 156 ][ 99 ],
   alphaCSR[ 156 ][ 100 ],
   alphaCSR[ 156 ][ 101 ],
   alphaCSR[ 156 ][ 102 ],
   alphaCSR[ 156 ][ 103 ],
   alphaCSR[ 156 ][ 104 ],
   alphaCSR[ 156 ][ 105 ],
   alphaCSR[ 156 ][ 106 ],
   alphaCSR[ 156 ][ 107 ],
   alphaCSR[ 156 ][ 108 ],
   alphaCSR[ 156 ][ 109 ],
   alphaCSR[ 156 ][ 110 ],
   alphaCSR[ 156 ][ 111 ],
   alphaCSR[ 156 ][ 112 ],
   alphaCSR[ 156 ][ 113 ],
   alphaCSR[ 156 ][ 114 ],
   alphaCSR[ 156 ][ 115 ],
   alphaCSR[ 156 ][ 116 ],
   alphaCSR[ 156 ][ 117 ],
   alphaCSR[ 156 ][ 118 ],
   alphaCSR[ 156 ][ 119 ],
   alphaCSR[ 156 ][ 120 ],
   alphaCSR[ 156 ][ 121 ],
   alphaCSR[ 156 ][ 122 ],
   alphaCSR[ 156 ][ 123 ],
   alphaCSR[ 156 ][ 124 ],
   alphaCSR[ 156 ][ 125 ],
   alphaCSR[ 156 ][ 126 ],
   alphaCSR[ 156 ][ 127 ],
   alphaCSR[ 156 ][ 128 ],
   alphaCSR[ 156 ][ 129 ],
   alphaCSR[ 156 ][ 130 ],
   alphaCSR[ 156 ][ 131 ],
   alphaCSR[ 156 ][ 132 ],
   alphaCSR[ 156 ][ 133 ],
   alphaCSR[ 156 ][ 134 ],
   alphaCSR[ 156 ][ 135 ],
   alphaCSR[ 156 ][ 136 ],
   alphaCSR[ 156 ][ 137 ],
   alphaCSR[ 156 ][ 138 ],
   alphaCSR[ 156 ][ 139 ],
   alphaCSR[ 156 ][ 140 ],
   alphaCSR[ 156 ][ 141 ],
   alphaCSR[ 156 ][ 142 ],
   alphaCSR[ 156 ][ 143 ],
   alphaCSR[ 156 ][ 144 ],
   alphaCSR[ 156 ][ 145 ],
   alphaCSR[ 156 ][ 146 ],
   alphaCSR[ 156 ][ 147 ],
   alphaCSR[ 156 ][ 148 ],
   alphaCSR[ 156 ][ 149 ],
   alphaCSR[ 156 ][ 150 ],
   alphaCSR[ 156 ][ 151 ],
   alphaCSR[ 156 ][ 152 ],
   alphaCSR[ 156 ][ 153 ],
   alphaCSR[ 156 ][ 154 ],
   alphaCSR[ 156 ][ 155 ],
   alphaCSR[ 156 ][ 156 ],
   alphaCSR[ 156 ][ 157 ],
   alphaCSR[ 156 ][ 158 ],
   alphaCSR[ 156 ][ 159 ],
   alphaCSR[ 156 ][ 160 ],
   alphaCSR[ 156 ][ 161 ],
   alphaCSR[ 156 ][ 162 ],
   alphaCSR[ 156 ][ 163 ],
   alphaCSR[ 156 ][ 164 ],
   alphaCSR[ 156 ][ 165 ],
   alphaCSR[ 156 ][ 166 ],
   alphaCSR[ 156 ][ 167 ],
   alphaCSR[ 156 ][ 168 ],
   alphaCSR[ 156 ][ 169 ],
   alphaCSR[ 156 ][ 170 ],
   alphaCSR[ 156 ][ 171 ],
   alphaCSR[ 156 ][ 172 ],
   alphaCSR[ 156 ][ 173 ],
   alphaCSR[ 156 ][ 174 ],
   alphaCSR[ 156 ][ 175 ],
   alphaCSR[ 156 ][ 176 ],
   alphaCSR[ 156 ][ 177 ],
   alphaCSR[ 156 ][ 178 ],
   alphaCSR[ 156 ][ 179 ],
   alphaCSR[ 156 ][ 180 ],
   alphaCSR[ 156 ][ 181 ],
   alphaCSR[ 156 ][ 182 ],
   alphaCSR[ 156 ][ 183 ],
   alphaCSR[ 156 ][ 184 ],
   alphaCSR[ 156 ][ 185 ],
   alphaCSR[ 156 ][ 186 ],
   alphaCSR[ 156 ][ 187 ],
   alphaCSR[ 156 ][ 188 ],
   alphaCSR[ 156 ][ 189 ],
   alphaCSR[ 156 ][ 190 ],
   alphaCSR[ 156 ][ 191 ],
   alphaCSR[ 156 ][ 192 ],
   alphaCSR[ 156 ][ 193 ],
   alphaCSR[ 156 ][ 194 ],
   alphaCSR[ 156 ][ 195 ],
   alphaCSR[ 156 ][ 196 ],
   alphaCSR[ 156 ][ 197 ],
   alphaCSR[ 156 ][ 198 ],
   alphaCSR[ 156 ][ 199 ],
   alphaCSR[ 156 ][ 200 ],
   alphaCSR[ 156 ][ 201 ],
   alphaCSR[ 156 ][ 202 ],
   alphaCSR[ 156 ][ 203 ],
   alphaCSR[ 156 ][ 204 ],
   alphaCSR[ 156 ][ 205 ],
   alphaCSR[ 156 ][ 206 ],
   alphaCSR[ 156 ][ 207 ],
   alphaCSR[ 156 ][ 208 ],
   alphaCSR[ 156 ][ 209 ],
   alphaCSR[ 156 ][ 210 ],
   alphaCSR[ 156 ][ 211 ],
   alphaCSR[ 156 ][ 212 ],
   alphaCSR[ 156 ][ 213 ],
   alphaCSR[ 156 ][ 214 ],
   alphaCSR[ 156 ][ 215 ],
   alphaCSR[ 156 ][ 216 ],
   alphaCSR[ 156 ][ 217 ],
   alphaCSR[ 156 ][ 218 ],
   alphaCSR[ 156 ][ 219 ],
   alphaCSR[ 156 ][ 220 ],
   alphaCSR[ 156 ][ 221 ],
   alphaCSR[ 156 ][ 222 ],
   alphaCSR[ 156 ][ 223 ],
   alphaCSR[ 156 ][ 224 ],
   alphaCSR[ 156 ][ 225 ],
   alphaCSR[ 156 ][ 226 ],
   alphaCSR[ 156 ][ 227 ],
   alphaCSR[ 156 ][ 228 ],
   alphaCSR[ 156 ][ 229 ],
   alphaCSR[ 156 ][ 230 ],
   alphaCSR[ 156 ][ 231 ],
   alphaCSR[ 156 ][ 232 ],
   alphaCSR[ 156 ][ 233 ],
   alphaCSR[ 156 ][ 234 ],
   alphaCSR[ 156 ][ 235 ],
   alphaCSR[ 156 ][ 236 ],
   alphaCSR[ 156 ][ 237 ],
   alphaCSR[ 156 ][ 238 ],
   alphaCSR[ 156 ][ 239 ],
   alphaCSR[ 156 ][ 240 ],
   alphaCSR[ 156 ][ 241 ],
   alphaCSR[ 156 ][ 242 ],
   alphaCSR[ 156 ][ 243 ],
   alphaCSR[ 156 ][ 244 ],
   alphaCSR[ 156 ][ 245 ],
   alphaCSR[ 156 ][ 246 ],
   alphaCSR[ 156 ][ 247 ],
   alphaCSR[ 156 ][ 248 ],
   alphaCSR[ 156 ][ 249 ],
   alphaCSR[ 156 ][ 250 ],
   alphaCSR[ 156 ][ 251 ],
   alphaCSR[ 156 ][ 252 ],
   alphaCSR[ 156 ][ 253 ],
   alphaCSR[ 156 ][ 254 ],
   alphaCSR[ 156 ][ 255 ],
   alphaCSR[ 156 ][ 256 ],
   alphaCSR[ 156 ][ 257 ],
   alphaCSR[ 156 ][ 258 ],
   alphaCSR[ 156 ][ 259 ],
   alphaCSR[ 156 ][ 260 ],
   alphaCSR[ 156 ][ 261 ],
   alphaCSR[ 156 ][ 262 ],
   alphaCSR[ 156 ][ 263 ],
   alphaCSR[ 156 ][ 264 ],
   alphaCSR[ 156 ][ 265 ],
   alphaCSR[ 156 ][ 266 ],
   alphaCSR[ 156 ][ 267 ],
   alphaCSR[ 156 ][ 268 ],
   alphaCSR[ 156 ][ 269 ],
   alphaCSR[ 156 ][ 270 ],
   alphaCSR[ 156 ][ 271 ],
   alphaCSR[ 156 ][ 272 ],
   alphaCSR[ 156 ][ 273 ],
   alphaCSR[ 156 ][ 274 ],
   alphaCSR[ 156 ][ 275 ],
   alphaCSR[ 156 ][ 276 ],
   alphaCSR[ 156 ][ 277 ],
   alphaCSR[ 156 ][ 278 ],
   alphaCSR[ 156 ][ 279 ],
   alphaCSR[ 156 ][ 280 ],
   alphaCSR[ 156 ][ 281 ],
   alphaCSR[ 156 ][ 282 ],
   alphaCSR[ 156 ][ 283 ],
   alphaCSR[ 156 ][ 284 ],
   alphaCSR[ 156 ][ 285 ],
   alphaCSR[ 156 ][ 286 ],
   alphaCSR[ 156 ][ 287 ],
   alphaCSR[ 156 ][ 288 ],
   alphaCSR[ 156 ][ 289 ],
   alphaCSR[ 156 ][ 290 ],
   alphaCSR[ 156 ][ 291 ],
   alphaCSR[ 156 ][ 292 ],
   alphaCSR[ 156 ][ 293 ],
   alphaCSR[ 156 ][ 294 ],
   alphaCSR[ 156 ][ 295 ],
   alphaCSR[ 156 ][ 296 ],
   alphaCSR[ 156 ][ 297 ],
   alphaCSR[ 156 ][ 298 ],
   alphaCSR[ 156 ][ 299 ],
   alphaCSR[ 156 ][ 300 ],
   alphaCSR[ 156 ][ 301 ],
   alphaCSR[ 156 ][ 302 ],
   alphaCSR[ 156 ][ 303 ],
   alphaCSR[ 156 ][ 304 ],
   alphaCSR[ 156 ][ 305 ],
   alphaCSR[ 156 ][ 306 ],
   alphaCSR[ 156 ][ 307 ],
   alphaCSR[ 156 ][ 308 ],
   alphaCSR[ 156 ][ 309 ],
   alphaCSR[ 156 ][ 310 ],
   alphaCSR[ 156 ][ 311 ],
   alphaCSR[ 156 ][ 312 ],
   alphaCSR[ 156 ][ 313 ],
   alphaCSR[ 156 ][ 314 ],
   alphaCSR[ 156 ][ 315 ],
   alphaCSR[ 156 ][ 316 ],
   alphaCSR[ 156 ][ 317 ],
   alphaCSR[ 156 ][ 318 ],
   alphaCSR[ 156 ][ 319 ],
   alphaCSR[ 156 ][ 320 ],
   alphaCSR[ 156 ][ 321 ],
   alphaCSR[ 156 ][ 322 ],
   alphaCSR[ 156 ][ 323 ],
   alphaCSR[ 156 ][ 324 ],
   alphaCSR[ 156 ][ 325 ],
   alphaCSR[ 156 ][ 326 ],
   alphaCSR[ 156 ][ 327 ],
   alphaCSR[ 156 ][ 328 ],
   alphaCSR[ 156 ][ 329 ],
   alphaCSR[ 156 ][ 330 ],
   alphaCSR[ 156 ][ 331 ],
   alphaCSR[ 156 ][ 332 ],
   alphaCSR[ 156 ][ 333 ],
   alphaCSR[ 156 ][ 334 ],
   alphaCSR[ 156 ][ 335 ],
   alphaCSR[ 156 ][ 336 ],
   alphaCSR[ 156 ][ 337 ],
   alphaCSR[ 156 ][ 338 ],
   alphaCSR[ 156 ][ 339 ],
   alphaCSR[ 156 ][ 340 ],
   alphaCSR[ 156 ][ 341 ],
   alphaCSR[ 156 ][ 342 ],
   alphaCSR[ 156 ][ 343 ],
   alphaCSR[ 156 ][ 344 ],
   alphaCSR[ 156 ][ 345 ],
   alphaCSR[ 156 ][ 346 ],
   alphaCSR[ 156 ][ 347 ],
   alphaCSR[ 156 ][ 348 ],
   alphaCSR[ 156 ][ 349 ],
   alphaCSR[ 156 ][ 350 ],
   alphaCSR[ 156 ][ 351 ],
   alphaCSR[ 156 ][ 352 ],
   alphaCSR[ 156 ][ 353 ],
   alphaCSR[ 156 ][ 354 ],
   alphaCSR[ 156 ][ 355 ],
   alphaCSR[ 156 ][ 356 ],
   alphaCSR[ 156 ][ 357 ],
   alphaCSR[ 156 ][ 358 ],
   alphaCSR[ 156 ][ 359 ],
   alphaCSR[ 156 ][ 360 ],
   alphaCSR[ 156 ][ 361 ],
   alphaCSR[ 156 ][ 362 ],
   alphaCSR[ 156 ][ 363 ],
   alphaCSR[ 156 ][ 364 ],
   alphaCSR[ 156 ][ 365 ],
   alphaCSR[ 156 ][ 366 ],
   alphaCSR[ 156 ][ 367 ],
   alphaCSR[ 156 ][ 368 ],
   alphaCSR[ 156 ][ 369 ],
   alphaCSR[ 156 ][ 370 ],
   alphaCSR[ 156 ][ 371 ],
   alphaCSR[ 156 ][ 372 ],
   alphaCSR[ 156 ][ 373 ],
   alphaCSR[ 156 ][ 374 ],
   alphaCSR[ 156 ][ 375 ],
   alphaCSR[ 156 ][ 376 ],
   alphaCSR[ 156 ][ 377 ],
   alphaCSR[ 156 ][ 378 ],
   alphaCSR[ 156 ][ 379 ],
   alphaCSR[ 156 ][ 380 ],
   alphaCSR[ 156 ][ 381 ],
   alphaCSR[ 156 ][ 382 ],
   alphaCSR[ 156 ][ 383 ],
   alphaCSR[ 157 ][ 0 ],
   alphaCSR[ 157 ][ 1 ],
   alphaCSR[ 157 ][ 2 ],
   alphaCSR[ 157 ][ 3 ],
   alphaCSR[ 157 ][ 4 ],
   alphaCSR[ 157 ][ 5 ],
   alphaCSR[ 157 ][ 6 ],
   alphaCSR[ 157 ][ 7 ],
   alphaCSR[ 157 ][ 8 ],
   alphaCSR[ 157 ][ 9 ],
   alphaCSR[ 157 ][ 10 ],
   alphaCSR[ 157 ][ 11 ],
   alphaCSR[ 157 ][ 12 ],
   alphaCSR[ 157 ][ 13 ],
   alphaCSR[ 157 ][ 14 ],
   alphaCSR[ 157 ][ 15 ],
   alphaCSR[ 157 ][ 16 ],
   alphaCSR[ 157 ][ 17 ],
   alphaCSR[ 157 ][ 18 ],
   alphaCSR[ 157 ][ 19 ],
   alphaCSR[ 157 ][ 20 ],
   alphaCSR[ 157 ][ 21 ],
   alphaCSR[ 157 ][ 22 ],
   alphaCSR[ 157 ][ 23 ],
   alphaCSR[ 157 ][ 24 ],
   alphaCSR[ 157 ][ 25 ],
   alphaCSR[ 157 ][ 26 ],
   alphaCSR[ 157 ][ 27 ],
   alphaCSR[ 157 ][ 28 ],
   alphaCSR[ 157 ][ 29 ],
   alphaCSR[ 157 ][ 30 ],
   alphaCSR[ 157 ][ 31 ],
   alphaCSR[ 157 ][ 32 ],
   alphaCSR[ 157 ][ 33 ],
   alphaCSR[ 157 ][ 34 ],
   alphaCSR[ 157 ][ 35 ],
   alphaCSR[ 157 ][ 36 ],
   alphaCSR[ 157 ][ 37 ],
   alphaCSR[ 157 ][ 38 ],
   alphaCSR[ 157 ][ 39 ],
   alphaCSR[ 157 ][ 40 ],
   alphaCSR[ 157 ][ 41 ],
   alphaCSR[ 157 ][ 42 ],
   alphaCSR[ 157 ][ 43 ],
   alphaCSR[ 157 ][ 44 ],
   alphaCSR[ 157 ][ 45 ],
   alphaCSR[ 157 ][ 46 ],
   alphaCSR[ 157 ][ 47 ],
   alphaCSR[ 157 ][ 48 ],
   alphaCSR[ 157 ][ 49 ],
   alphaCSR[ 157 ][ 50 ],
   alphaCSR[ 157 ][ 51 ],
   alphaCSR[ 157 ][ 52 ],
   alphaCSR[ 157 ][ 53 ],
   alphaCSR[ 157 ][ 54 ],
   alphaCSR[ 157 ][ 55 ],
   alphaCSR[ 157 ][ 56 ],
   alphaCSR[ 157 ][ 57 ],
   alphaCSR[ 157 ][ 58 ],
   alphaCSR[ 157 ][ 59 ],
   alphaCSR[ 157 ][ 60 ],
   alphaCSR[ 157 ][ 61 ],
   alphaCSR[ 157 ][ 62 ],
   alphaCSR[ 157 ][ 63 ],
   alphaCSR[ 157 ][ 64 ],
   alphaCSR[ 157 ][ 65 ],
   alphaCSR[ 157 ][ 66 ],
   alphaCSR[ 157 ][ 67 ],
   alphaCSR[ 157 ][ 68 ],
   alphaCSR[ 157 ][ 69 ],
   alphaCSR[ 157 ][ 70 ],
   alphaCSR[ 157 ][ 71 ],
   alphaCSR[ 157 ][ 72 ],
   alphaCSR[ 157 ][ 73 ],
   alphaCSR[ 157 ][ 74 ],
   alphaCSR[ 157 ][ 75 ],
   alphaCSR[ 157 ][ 76 ],
   alphaCSR[ 157 ][ 77 ],
   alphaCSR[ 157 ][ 78 ],
   alphaCSR[ 157 ][ 79 ],
   alphaCSR[ 157 ][ 80 ],
   alphaCSR[ 157 ][ 81 ],
   alphaCSR[ 157 ][ 82 ],
   alphaCSR[ 157 ][ 83 ],
   alphaCSR[ 157 ][ 84 ],
   alphaCSR[ 157 ][ 85 ],
   alphaCSR[ 157 ][ 86 ],
   alphaCSR[ 157 ][ 87 ],
   alphaCSR[ 157 ][ 88 ],
   alphaCSR[ 157 ][ 89 ],
   alphaCSR[ 157 ][ 90 ],
   alphaCSR[ 157 ][ 91 ],
   alphaCSR[ 157 ][ 92 ],
   alphaCSR[ 157 ][ 93 ],
   alphaCSR[ 157 ][ 94 ],
   alphaCSR[ 157 ][ 95 ],
   alphaCSR[ 157 ][ 96 ],
   alphaCSR[ 157 ][ 97 ],
   alphaCSR[ 157 ][ 98 ],
   alphaCSR[ 157 ][ 99 ],
   alphaCSR[ 157 ][ 100 ],
   alphaCSR[ 157 ][ 101 ],
   alphaCSR[ 157 ][ 102 ],
   alphaCSR[ 157 ][ 103 ],
   alphaCSR[ 157 ][ 104 ],
   alphaCSR[ 157 ][ 105 ],
   alphaCSR[ 157 ][ 106 ],
   alphaCSR[ 157 ][ 107 ],
   alphaCSR[ 157 ][ 108 ],
   alphaCSR[ 157 ][ 109 ],
   alphaCSR[ 157 ][ 110 ],
   alphaCSR[ 157 ][ 111 ],
   alphaCSR[ 157 ][ 112 ],
   alphaCSR[ 157 ][ 113 ],
   alphaCSR[ 157 ][ 114 ],
   alphaCSR[ 157 ][ 115 ],
   alphaCSR[ 157 ][ 116 ],
   alphaCSR[ 157 ][ 117 ],
   alphaCSR[ 157 ][ 118 ],
   alphaCSR[ 157 ][ 119 ],
   alphaCSR[ 157 ][ 120 ],
   alphaCSR[ 157 ][ 121 ],
   alphaCSR[ 157 ][ 122 ],
   alphaCSR[ 157 ][ 123 ],
   alphaCSR[ 157 ][ 124 ],
   alphaCSR[ 157 ][ 125 ],
   alphaCSR[ 157 ][ 126 ],
   alphaCSR[ 157 ][ 127 ],
   alphaCSR[ 157 ][ 128 ],
   alphaCSR[ 157 ][ 129 ],
   alphaCSR[ 157 ][ 130 ],
   alphaCSR[ 157 ][ 131 ],
   alphaCSR[ 157 ][ 132 ],
   alphaCSR[ 157 ][ 133 ],
   alphaCSR[ 157 ][ 134 ],
   alphaCSR[ 157 ][ 135 ],
   alphaCSR[ 157 ][ 136 ],
   alphaCSR[ 157 ][ 137 ],
   alphaCSR[ 157 ][ 138 ],
   alphaCSR[ 157 ][ 139 ],
   alphaCSR[ 157 ][ 140 ],
   alphaCSR[ 157 ][ 141 ],
   alphaCSR[ 157 ][ 142 ],
   alphaCSR[ 157 ][ 143 ],
   alphaCSR[ 157 ][ 144 ],
   alphaCSR[ 157 ][ 145 ],
   alphaCSR[ 157 ][ 146 ],
   alphaCSR[ 157 ][ 147 ],
   alphaCSR[ 157 ][ 148 ],
   alphaCSR[ 157 ][ 149 ],
   alphaCSR[ 157 ][ 150 ],
   alphaCSR[ 157 ][ 151 ],
   alphaCSR[ 157 ][ 152 ],
   alphaCSR[ 157 ][ 153 ],
   alphaCSR[ 157 ][ 154 ],
   alphaCSR[ 157 ][ 155 ],
   alphaCSR[ 157 ][ 156 ],
   alphaCSR[ 157 ][ 157 ],
   alphaCSR[ 157 ][ 158 ],
   alphaCSR[ 157 ][ 159 ],
   alphaCSR[ 157 ][ 160 ],
   alphaCSR[ 157 ][ 161 ],
   alphaCSR[ 157 ][ 162 ],
   alphaCSR[ 157 ][ 163 ],
   alphaCSR[ 157 ][ 164 ],
   alphaCSR[ 157 ][ 165 ],
   alphaCSR[ 157 ][ 166 ],
   alphaCSR[ 157 ][ 167 ],
   alphaCSR[ 157 ][ 168 ],
   alphaCSR[ 157 ][ 169 ],
   alphaCSR[ 157 ][ 170 ],
   alphaCSR[ 157 ][ 171 ],
   alphaCSR[ 157 ][ 172 ],
   alphaCSR[ 157 ][ 173 ],
   alphaCSR[ 157 ][ 174 ],
   alphaCSR[ 157 ][ 175 ],
   alphaCSR[ 157 ][ 176 ],
   alphaCSR[ 157 ][ 177 ],
   alphaCSR[ 157 ][ 178 ],
   alphaCSR[ 157 ][ 179 ],
   alphaCSR[ 157 ][ 180 ],
   alphaCSR[ 157 ][ 181 ],
   alphaCSR[ 157 ][ 182 ],
   alphaCSR[ 157 ][ 183 ],
   alphaCSR[ 157 ][ 184 ],
   alphaCSR[ 157 ][ 185 ],
   alphaCSR[ 157 ][ 186 ],
   alphaCSR[ 157 ][ 187 ],
   alphaCSR[ 157 ][ 188 ],
   alphaCSR[ 157 ][ 189 ],
   alphaCSR[ 157 ][ 190 ],
   alphaCSR[ 157 ][ 191 ],
   alphaCSR[ 157 ][ 192 ],
   alphaCSR[ 157 ][ 193 ],
   alphaCSR[ 157 ][ 194 ],
   alphaCSR[ 157 ][ 195 ],
   alphaCSR[ 157 ][ 196 ],
   alphaCSR[ 157 ][ 197 ],
   alphaCSR[ 157 ][ 198 ],
   alphaCSR[ 157 ][ 199 ],
   alphaCSR[ 157 ][ 200 ],
   alphaCSR[ 157 ][ 201 ],
   alphaCSR[ 157 ][ 202 ],
   alphaCSR[ 157 ][ 203 ],
   alphaCSR[ 157 ][ 204 ],
   alphaCSR[ 157 ][ 205 ],
   alphaCSR[ 157 ][ 206 ],
   alphaCSR[ 157 ][ 207 ],
   alphaCSR[ 157 ][ 208 ],
   alphaCSR[ 157 ][ 209 ],
   alphaCSR[ 157 ][ 210 ],
   alphaCSR[ 157 ][ 211 ],
   alphaCSR[ 157 ][ 212 ],
   alphaCSR[ 157 ][ 213 ],
   alphaCSR[ 157 ][ 214 ],
   alphaCSR[ 157 ][ 215 ],
   alphaCSR[ 157 ][ 216 ],
   alphaCSR[ 157 ][ 217 ],
   alphaCSR[ 157 ][ 218 ],
   alphaCSR[ 157 ][ 219 ],
   alphaCSR[ 157 ][ 220 ],
   alphaCSR[ 157 ][ 221 ],
   alphaCSR[ 157 ][ 222 ],
   alphaCSR[ 157 ][ 223 ],
   alphaCSR[ 157 ][ 224 ],
   alphaCSR[ 157 ][ 225 ],
   alphaCSR[ 157 ][ 226 ],
   alphaCSR[ 157 ][ 227 ],
   alphaCSR[ 157 ][ 228 ],
   alphaCSR[ 157 ][ 229 ],
   alphaCSR[ 157 ][ 230 ],
   alphaCSR[ 157 ][ 231 ],
   alphaCSR[ 157 ][ 232 ],
   alphaCSR[ 157 ][ 233 ],
   alphaCSR[ 157 ][ 234 ],
   alphaCSR[ 157 ][ 235 ],
   alphaCSR[ 157 ][ 236 ],
   alphaCSR[ 157 ][ 237 ],
   alphaCSR[ 157 ][ 238 ],
   alphaCSR[ 157 ][ 239 ],
   alphaCSR[ 157 ][ 240 ],
   alphaCSR[ 157 ][ 241 ],
   alphaCSR[ 157 ][ 242 ],
   alphaCSR[ 157 ][ 243 ],
   alphaCSR[ 157 ][ 244 ],
   alphaCSR[ 157 ][ 245 ],
   alphaCSR[ 157 ][ 246 ],
   alphaCSR[ 157 ][ 247 ],
   alphaCSR[ 157 ][ 248 ],
   alphaCSR[ 157 ][ 249 ],
   alphaCSR[ 157 ][ 250 ],
   alphaCSR[ 157 ][ 251 ],
   alphaCSR[ 157 ][ 252 ],
   alphaCSR[ 157 ][ 253 ],
   alphaCSR[ 157 ][ 254 ],
   alphaCSR[ 157 ][ 255 ],
   alphaCSR[ 157 ][ 256 ],
   alphaCSR[ 157 ][ 257 ],
   alphaCSR[ 157 ][ 258 ],
   alphaCSR[ 157 ][ 259 ],
   alphaCSR[ 157 ][ 260 ],
   alphaCSR[ 157 ][ 261 ],
   alphaCSR[ 157 ][ 262 ],
   alphaCSR[ 157 ][ 263 ],
   alphaCSR[ 157 ][ 264 ],
   alphaCSR[ 157 ][ 265 ],
   alphaCSR[ 157 ][ 266 ],
   alphaCSR[ 157 ][ 267 ],
   alphaCSR[ 157 ][ 268 ],
   alphaCSR[ 157 ][ 269 ],
   alphaCSR[ 157 ][ 270 ],
   alphaCSR[ 157 ][ 271 ],
   alphaCSR[ 157 ][ 272 ],
   alphaCSR[ 157 ][ 273 ],
   alphaCSR[ 157 ][ 274 ],
   alphaCSR[ 157 ][ 275 ],
   alphaCSR[ 157 ][ 276 ],
   alphaCSR[ 157 ][ 277 ],
   alphaCSR[ 157 ][ 278 ],
   alphaCSR[ 157 ][ 279 ],
   alphaCSR[ 157 ][ 280 ],
   alphaCSR[ 157 ][ 281 ],
   alphaCSR[ 157 ][ 282 ],
   alphaCSR[ 157 ][ 283 ],
   alphaCSR[ 157 ][ 284 ],
   alphaCSR[ 157 ][ 285 ],
   alphaCSR[ 157 ][ 286 ],
   alphaCSR[ 157 ][ 287 ],
   alphaCSR[ 157 ][ 288 ],
   alphaCSR[ 157 ][ 289 ],
   alphaCSR[ 157 ][ 290 ],
   alphaCSR[ 157 ][ 291 ],
   alphaCSR[ 157 ][ 292 ],
   alphaCSR[ 157 ][ 293 ],
   alphaCSR[ 157 ][ 294 ],
   alphaCSR[ 157 ][ 295 ],
   alphaCSR[ 157 ][ 296 ],
   alphaCSR[ 157 ][ 297 ],
   alphaCSR[ 157 ][ 298 ],
   alphaCSR[ 157 ][ 299 ],
   alphaCSR[ 157 ][ 300 ],
   alphaCSR[ 157 ][ 301 ],
   alphaCSR[ 157 ][ 302 ],
   alphaCSR[ 157 ][ 303 ],
   alphaCSR[ 157 ][ 304 ],
   alphaCSR[ 157 ][ 305 ],
   alphaCSR[ 157 ][ 306 ],
   alphaCSR[ 157 ][ 307 ],
   alphaCSR[ 157 ][ 308 ],
   alphaCSR[ 157 ][ 309 ],
   alphaCSR[ 157 ][ 310 ],
   alphaCSR[ 157 ][ 311 ],
   alphaCSR[ 157 ][ 312 ],
   alphaCSR[ 157 ][ 313 ],
   alphaCSR[ 157 ][ 314 ],
   alphaCSR[ 157 ][ 315 ],
   alphaCSR[ 157 ][ 316 ],
   alphaCSR[ 157 ][ 317 ],
   alphaCSR[ 157 ][ 318 ],
   alphaCSR[ 157 ][ 319 ],
   alphaCSR[ 157 ][ 320 ],
   alphaCSR[ 157 ][ 321 ],
   alphaCSR[ 157 ][ 322 ],
   alphaCSR[ 157 ][ 323 ],
   alphaCSR[ 157 ][ 324 ],
   alphaCSR[ 157 ][ 325 ],
   alphaCSR[ 157 ][ 326 ],
   alphaCSR[ 157 ][ 327 ],
   alphaCSR[ 157 ][ 328 ],
   alphaCSR[ 157 ][ 329 ],
   alphaCSR[ 157 ][ 330 ],
   alphaCSR[ 157 ][ 331 ],
   alphaCSR[ 157 ][ 332 ],
   alphaCSR[ 157 ][ 333 ],
   alphaCSR[ 157 ][ 334 ],
   alphaCSR[ 157 ][ 335 ],
   alphaCSR[ 157 ][ 336 ],
   alphaCSR[ 157 ][ 337 ],
   alphaCSR[ 157 ][ 338 ],
   alphaCSR[ 157 ][ 339 ],
   alphaCSR[ 157 ][ 340 ],
   alphaCSR[ 157 ][ 341 ],
   alphaCSR[ 157 ][ 342 ],
   alphaCSR[ 157 ][ 343 ],
   alphaCSR[ 157 ][ 344 ],
   alphaCSR[ 157 ][ 345 ],
   alphaCSR[ 157 ][ 346 ],
   alphaCSR[ 157 ][ 347 ],
   alphaCSR[ 157 ][ 348 ],
   alphaCSR[ 157 ][ 349 ],
   alphaCSR[ 157 ][ 350 ],
   alphaCSR[ 157 ][ 351 ],
   alphaCSR[ 157 ][ 352 ],
   alphaCSR[ 157 ][ 353 ],
   alphaCSR[ 157 ][ 354 ],
   alphaCSR[ 157 ][ 355 ],
   alphaCSR[ 157 ][ 356 ],
   alphaCSR[ 157 ][ 357 ],
   alphaCSR[ 157 ][ 358 ],
   alphaCSR[ 157 ][ 359 ],
   alphaCSR[ 157 ][ 360 ],
   alphaCSR[ 157 ][ 361 ],
   alphaCSR[ 157 ][ 362 ],
   alphaCSR[ 157 ][ 363 ],
   alphaCSR[ 157 ][ 364 ],
   alphaCSR[ 157 ][ 365 ],
   alphaCSR[ 157 ][ 366 ],
   alphaCSR[ 157 ][ 367 ],
   alphaCSR[ 157 ][ 368 ],
   alphaCSR[ 157 ][ 369 ],
   alphaCSR[ 157 ][ 370 ],
   alphaCSR[ 157 ][ 371 ],
   alphaCSR[ 157 ][ 372 ],
   alphaCSR[ 157 ][ 373 ],
   alphaCSR[ 157 ][ 374 ],
   alphaCSR[ 157 ][ 375 ],
   alphaCSR[ 157 ][ 376 ],
   alphaCSR[ 157 ][ 377 ],
   alphaCSR[ 157 ][ 378 ],
   alphaCSR[ 157 ][ 379 ],
   alphaCSR[ 157 ][ 380 ],
   alphaCSR[ 157 ][ 381 ],
   alphaCSR[ 157 ][ 382 ],
   alphaCSR[ 157 ][ 383 ],
   alphaCSR[ 158 ][ 0 ],
   alphaCSR[ 158 ][ 1 ],
   alphaCSR[ 158 ][ 2 ],
   alphaCSR[ 158 ][ 3 ],
   alphaCSR[ 158 ][ 4 ],
   alphaCSR[ 158 ][ 5 ],
   alphaCSR[ 158 ][ 6 ],
   alphaCSR[ 158 ][ 7 ],
   alphaCSR[ 158 ][ 8 ],
   alphaCSR[ 158 ][ 9 ],
   alphaCSR[ 158 ][ 10 ],
   alphaCSR[ 158 ][ 11 ],
   alphaCSR[ 158 ][ 12 ],
   alphaCSR[ 158 ][ 13 ],
   alphaCSR[ 158 ][ 14 ],
   alphaCSR[ 158 ][ 15 ],
   alphaCSR[ 158 ][ 16 ],
   alphaCSR[ 158 ][ 17 ],
   alphaCSR[ 158 ][ 18 ],
   alphaCSR[ 158 ][ 19 ],
   alphaCSR[ 158 ][ 20 ],
   alphaCSR[ 158 ][ 21 ],
   alphaCSR[ 158 ][ 22 ],
   alphaCSR[ 158 ][ 23 ],
   alphaCSR[ 158 ][ 24 ],
   alphaCSR[ 158 ][ 25 ],
   alphaCSR[ 158 ][ 26 ],
   alphaCSR[ 158 ][ 27 ],
   alphaCSR[ 158 ][ 28 ],
   alphaCSR[ 158 ][ 29 ],
   alphaCSR[ 158 ][ 30 ],
   alphaCSR[ 158 ][ 31 ],
   alphaCSR[ 158 ][ 32 ],
   alphaCSR[ 158 ][ 33 ],
   alphaCSR[ 158 ][ 34 ],
   alphaCSR[ 158 ][ 35 ],
   alphaCSR[ 158 ][ 36 ],
   alphaCSR[ 158 ][ 37 ],
   alphaCSR[ 158 ][ 38 ],
   alphaCSR[ 158 ][ 39 ],
   alphaCSR[ 158 ][ 40 ],
   alphaCSR[ 158 ][ 41 ],
   alphaCSR[ 158 ][ 42 ],
   alphaCSR[ 158 ][ 43 ],
   alphaCSR[ 158 ][ 44 ],
   alphaCSR[ 158 ][ 45 ],
   alphaCSR[ 158 ][ 46 ],
   alphaCSR[ 158 ][ 47 ],
   alphaCSR[ 158 ][ 48 ],
   alphaCSR[ 158 ][ 49 ],
   alphaCSR[ 158 ][ 50 ],
   alphaCSR[ 158 ][ 51 ],
   alphaCSR[ 158 ][ 52 ],
   alphaCSR[ 158 ][ 53 ],
   alphaCSR[ 158 ][ 54 ],
   alphaCSR[ 158 ][ 55 ],
   alphaCSR[ 158 ][ 56 ],
   alphaCSR[ 158 ][ 57 ],
   alphaCSR[ 158 ][ 58 ],
   alphaCSR[ 158 ][ 59 ],
   alphaCSR[ 158 ][ 60 ],
   alphaCSR[ 158 ][ 61 ],
   alphaCSR[ 158 ][ 62 ],
   alphaCSR[ 158 ][ 63 ],
   alphaCSR[ 158 ][ 64 ],
   alphaCSR[ 158 ][ 65 ],
   alphaCSR[ 158 ][ 66 ],
   alphaCSR[ 158 ][ 67 ],
   alphaCSR[ 158 ][ 68 ],
   alphaCSR[ 158 ][ 69 ],
   alphaCSR[ 158 ][ 70 ],
   alphaCSR[ 158 ][ 71 ],
   alphaCSR[ 158 ][ 72 ],
   alphaCSR[ 158 ][ 73 ],
   alphaCSR[ 158 ][ 74 ],
   alphaCSR[ 158 ][ 75 ],
   alphaCSR[ 158 ][ 76 ],
   alphaCSR[ 158 ][ 77 ],
   alphaCSR[ 158 ][ 78 ],
   alphaCSR[ 158 ][ 79 ],
   alphaCSR[ 158 ][ 80 ],
   alphaCSR[ 158 ][ 81 ],
   alphaCSR[ 158 ][ 82 ],
   alphaCSR[ 158 ][ 83 ],
   alphaCSR[ 158 ][ 84 ],
   alphaCSR[ 158 ][ 85 ],
   alphaCSR[ 158 ][ 86 ],
   alphaCSR[ 158 ][ 87 ],
   alphaCSR[ 158 ][ 88 ],
   alphaCSR[ 158 ][ 89 ],
   alphaCSR[ 158 ][ 90 ],
   alphaCSR[ 158 ][ 91 ],
   alphaCSR[ 158 ][ 92 ],
   alphaCSR[ 158 ][ 93 ],
   alphaCSR[ 158 ][ 94 ],
   alphaCSR[ 158 ][ 95 ],
   alphaCSR[ 158 ][ 96 ],
   alphaCSR[ 158 ][ 97 ],
   alphaCSR[ 158 ][ 98 ],
   alphaCSR[ 158 ][ 99 ],
   alphaCSR[ 158 ][ 100 ],
   alphaCSR[ 158 ][ 101 ],
   alphaCSR[ 158 ][ 102 ],
   alphaCSR[ 158 ][ 103 ],
   alphaCSR[ 158 ][ 104 ],
   alphaCSR[ 158 ][ 105 ],
   alphaCSR[ 158 ][ 106 ],
   alphaCSR[ 158 ][ 107 ],
   alphaCSR[ 158 ][ 108 ],
   alphaCSR[ 158 ][ 109 ],
   alphaCSR[ 158 ][ 110 ],
   alphaCSR[ 158 ][ 111 ],
   alphaCSR[ 158 ][ 112 ],
   alphaCSR[ 158 ][ 113 ],
   alphaCSR[ 158 ][ 114 ],
   alphaCSR[ 158 ][ 115 ],
   alphaCSR[ 158 ][ 116 ],
   alphaCSR[ 158 ][ 117 ],
   alphaCSR[ 158 ][ 118 ],
   alphaCSR[ 158 ][ 119 ],
   alphaCSR[ 158 ][ 120 ],
   alphaCSR[ 158 ][ 121 ],
   alphaCSR[ 158 ][ 122 ],
   alphaCSR[ 158 ][ 123 ],
   alphaCSR[ 158 ][ 124 ],
   alphaCSR[ 158 ][ 125 ],
   alphaCSR[ 158 ][ 126 ],
   alphaCSR[ 158 ][ 127 ],
   alphaCSR[ 158 ][ 128 ],
   alphaCSR[ 158 ][ 129 ],
   alphaCSR[ 158 ][ 130 ],
   alphaCSR[ 158 ][ 131 ],
   alphaCSR[ 158 ][ 132 ],
   alphaCSR[ 158 ][ 133 ],
   alphaCSR[ 158 ][ 134 ],
   alphaCSR[ 158 ][ 135 ],
   alphaCSR[ 158 ][ 136 ],
   alphaCSR[ 158 ][ 137 ],
   alphaCSR[ 158 ][ 138 ],
   alphaCSR[ 158 ][ 139 ],
   alphaCSR[ 158 ][ 140 ],
   alphaCSR[ 158 ][ 141 ],
   alphaCSR[ 158 ][ 142 ],
   alphaCSR[ 158 ][ 143 ],
   alphaCSR[ 158 ][ 144 ],
   alphaCSR[ 158 ][ 145 ],
   alphaCSR[ 158 ][ 146 ],
   alphaCSR[ 158 ][ 147 ],
   alphaCSR[ 158 ][ 148 ],
   alphaCSR[ 158 ][ 149 ],
   alphaCSR[ 158 ][ 150 ],
   alphaCSR[ 158 ][ 151 ],
   alphaCSR[ 158 ][ 152 ],
   alphaCSR[ 158 ][ 153 ],
   alphaCSR[ 158 ][ 154 ],
   alphaCSR[ 158 ][ 155 ],
   alphaCSR[ 158 ][ 156 ],
   alphaCSR[ 158 ][ 157 ],
   alphaCSR[ 158 ][ 158 ],
   alphaCSR[ 158 ][ 159 ],
   alphaCSR[ 158 ][ 160 ],
   alphaCSR[ 158 ][ 161 ],
   alphaCSR[ 158 ][ 162 ],
   alphaCSR[ 158 ][ 163 ],
   alphaCSR[ 158 ][ 164 ],
   alphaCSR[ 158 ][ 165 ],
   alphaCSR[ 158 ][ 166 ],
   alphaCSR[ 158 ][ 167 ],
   alphaCSR[ 158 ][ 168 ],
   alphaCSR[ 158 ][ 169 ],
   alphaCSR[ 158 ][ 170 ],
   alphaCSR[ 158 ][ 171 ],
   alphaCSR[ 158 ][ 172 ],
   alphaCSR[ 158 ][ 173 ],
   alphaCSR[ 158 ][ 174 ],
   alphaCSR[ 158 ][ 175 ],
   alphaCSR[ 158 ][ 176 ],
   alphaCSR[ 158 ][ 177 ],
   alphaCSR[ 158 ][ 178 ],
   alphaCSR[ 158 ][ 179 ],
   alphaCSR[ 158 ][ 180 ],
   alphaCSR[ 158 ][ 181 ],
   alphaCSR[ 158 ][ 182 ],
   alphaCSR[ 158 ][ 183 ],
   alphaCSR[ 158 ][ 184 ],
   alphaCSR[ 158 ][ 185 ],
   alphaCSR[ 158 ][ 186 ],
   alphaCSR[ 158 ][ 187 ],
   alphaCSR[ 158 ][ 188 ],
   alphaCSR[ 158 ][ 189 ],
   alphaCSR[ 158 ][ 190 ],
   alphaCSR[ 158 ][ 191 ],
   alphaCSR[ 158 ][ 192 ],
   alphaCSR[ 158 ][ 193 ],
   alphaCSR[ 158 ][ 194 ],
   alphaCSR[ 158 ][ 195 ],
   alphaCSR[ 158 ][ 196 ],
   alphaCSR[ 158 ][ 197 ],
   alphaCSR[ 158 ][ 198 ],
   alphaCSR[ 158 ][ 199 ],
   alphaCSR[ 158 ][ 200 ],
   alphaCSR[ 158 ][ 201 ],
   alphaCSR[ 158 ][ 202 ],
   alphaCSR[ 158 ][ 203 ],
   alphaCSR[ 158 ][ 204 ],
   alphaCSR[ 158 ][ 205 ],
   alphaCSR[ 158 ][ 206 ],
   alphaCSR[ 158 ][ 207 ],
   alphaCSR[ 158 ][ 208 ],
   alphaCSR[ 158 ][ 209 ],
   alphaCSR[ 158 ][ 210 ],
   alphaCSR[ 158 ][ 211 ],
   alphaCSR[ 158 ][ 212 ],
   alphaCSR[ 158 ][ 213 ],
   alphaCSR[ 158 ][ 214 ],
   alphaCSR[ 158 ][ 215 ],
   alphaCSR[ 158 ][ 216 ],
   alphaCSR[ 158 ][ 217 ],
   alphaCSR[ 158 ][ 218 ],
   alphaCSR[ 158 ][ 219 ],
   alphaCSR[ 158 ][ 220 ],
   alphaCSR[ 158 ][ 221 ],
   alphaCSR[ 158 ][ 222 ],
   alphaCSR[ 158 ][ 223 ],
   alphaCSR[ 158 ][ 224 ],
   alphaCSR[ 158 ][ 225 ],
   alphaCSR[ 158 ][ 226 ],
   alphaCSR[ 158 ][ 227 ],
   alphaCSR[ 158 ][ 228 ],
   alphaCSR[ 158 ][ 229 ],
   alphaCSR[ 158 ][ 230 ],
   alphaCSR[ 158 ][ 231 ],
   alphaCSR[ 158 ][ 232 ],
   alphaCSR[ 158 ][ 233 ],
   alphaCSR[ 158 ][ 234 ],
   alphaCSR[ 158 ][ 235 ],
   alphaCSR[ 158 ][ 236 ],
   alphaCSR[ 158 ][ 237 ],
   alphaCSR[ 158 ][ 238 ],
   alphaCSR[ 158 ][ 239 ],
   alphaCSR[ 158 ][ 240 ],
   alphaCSR[ 158 ][ 241 ],
   alphaCSR[ 158 ][ 242 ],
   alphaCSR[ 158 ][ 243 ],
   alphaCSR[ 158 ][ 244 ],
   alphaCSR[ 158 ][ 245 ],
   alphaCSR[ 158 ][ 246 ],
   alphaCSR[ 158 ][ 247 ],
   alphaCSR[ 158 ][ 248 ],
   alphaCSR[ 158 ][ 249 ],
   alphaCSR[ 158 ][ 250 ],
   alphaCSR[ 158 ][ 251 ],
   alphaCSR[ 158 ][ 252 ],
   alphaCSR[ 158 ][ 253 ],
   alphaCSR[ 158 ][ 254 ],
   alphaCSR[ 158 ][ 255 ],
   alphaCSR[ 158 ][ 256 ],
   alphaCSR[ 158 ][ 257 ],
   alphaCSR[ 158 ][ 258 ],
   alphaCSR[ 158 ][ 259 ],
   alphaCSR[ 158 ][ 260 ],
   alphaCSR[ 158 ][ 261 ],
   alphaCSR[ 158 ][ 262 ],
   alphaCSR[ 158 ][ 263 ],
   alphaCSR[ 158 ][ 264 ],
   alphaCSR[ 158 ][ 265 ],
   alphaCSR[ 158 ][ 266 ],
   alphaCSR[ 158 ][ 267 ],
   alphaCSR[ 158 ][ 268 ],
   alphaCSR[ 158 ][ 269 ],
   alphaCSR[ 158 ][ 270 ],
   alphaCSR[ 158 ][ 271 ],
   alphaCSR[ 158 ][ 272 ],
   alphaCSR[ 158 ][ 273 ],
   alphaCSR[ 158 ][ 274 ],
   alphaCSR[ 158 ][ 275 ],
   alphaCSR[ 158 ][ 276 ],
   alphaCSR[ 158 ][ 277 ],
   alphaCSR[ 158 ][ 278 ],
   alphaCSR[ 158 ][ 279 ],
   alphaCSR[ 158 ][ 280 ],
   alphaCSR[ 158 ][ 281 ],
   alphaCSR[ 158 ][ 282 ],
   alphaCSR[ 158 ][ 283 ],
   alphaCSR[ 158 ][ 284 ],
   alphaCSR[ 158 ][ 285 ],
   alphaCSR[ 158 ][ 286 ],
   alphaCSR[ 158 ][ 287 ],
   alphaCSR[ 158 ][ 288 ],
   alphaCSR[ 158 ][ 289 ],
   alphaCSR[ 158 ][ 290 ],
   alphaCSR[ 158 ][ 291 ],
   alphaCSR[ 158 ][ 292 ],
   alphaCSR[ 158 ][ 293 ],
   alphaCSR[ 158 ][ 294 ],
   alphaCSR[ 158 ][ 295 ],
   alphaCSR[ 158 ][ 296 ],
   alphaCSR[ 158 ][ 297 ],
   alphaCSR[ 158 ][ 298 ],
   alphaCSR[ 158 ][ 299 ],
   alphaCSR[ 158 ][ 300 ],
   alphaCSR[ 158 ][ 301 ],
   alphaCSR[ 158 ][ 302 ],
   alphaCSR[ 158 ][ 303 ],
   alphaCSR[ 158 ][ 304 ],
   alphaCSR[ 158 ][ 305 ],
   alphaCSR[ 158 ][ 306 ],
   alphaCSR[ 158 ][ 307 ],
   alphaCSR[ 158 ][ 308 ],
   alphaCSR[ 158 ][ 309 ],
   alphaCSR[ 158 ][ 310 ],
   alphaCSR[ 158 ][ 311 ],
   alphaCSR[ 158 ][ 312 ],
   alphaCSR[ 158 ][ 313 ],
   alphaCSR[ 158 ][ 314 ],
   alphaCSR[ 158 ][ 315 ],
   alphaCSR[ 158 ][ 316 ],
   alphaCSR[ 158 ][ 317 ],
   alphaCSR[ 158 ][ 318 ],
   alphaCSR[ 158 ][ 319 ],
   alphaCSR[ 158 ][ 320 ],
   alphaCSR[ 158 ][ 321 ],
   alphaCSR[ 158 ][ 322 ],
   alphaCSR[ 158 ][ 323 ],
   alphaCSR[ 158 ][ 324 ],
   alphaCSR[ 158 ][ 325 ],
   alphaCSR[ 158 ][ 326 ],
   alphaCSR[ 158 ][ 327 ],
   alphaCSR[ 158 ][ 328 ],
   alphaCSR[ 158 ][ 329 ],
   alphaCSR[ 158 ][ 330 ],
   alphaCSR[ 158 ][ 331 ],
   alphaCSR[ 158 ][ 332 ],
   alphaCSR[ 158 ][ 333 ],
   alphaCSR[ 158 ][ 334 ],
   alphaCSR[ 158 ][ 335 ],
   alphaCSR[ 158 ][ 336 ],
   alphaCSR[ 158 ][ 337 ],
   alphaCSR[ 158 ][ 338 ],
   alphaCSR[ 158 ][ 339 ],
   alphaCSR[ 158 ][ 340 ],
   alphaCSR[ 158 ][ 341 ],
   alphaCSR[ 158 ][ 342 ],
   alphaCSR[ 158 ][ 343 ],
   alphaCSR[ 158 ][ 344 ],
   alphaCSR[ 158 ][ 345 ],
   alphaCSR[ 158 ][ 346 ],
   alphaCSR[ 158 ][ 347 ],
   alphaCSR[ 158 ][ 348 ],
   alphaCSR[ 158 ][ 349 ],
   alphaCSR[ 158 ][ 350 ],
   alphaCSR[ 158 ][ 351 ],
   alphaCSR[ 158 ][ 352 ],
   alphaCSR[ 158 ][ 353 ],
   alphaCSR[ 158 ][ 354 ],
   alphaCSR[ 158 ][ 355 ],
   alphaCSR[ 158 ][ 356 ],
   alphaCSR[ 158 ][ 357 ],
   alphaCSR[ 158 ][ 358 ],
   alphaCSR[ 158 ][ 359 ],
   alphaCSR[ 158 ][ 360 ],
   alphaCSR[ 158 ][ 361 ],
   alphaCSR[ 158 ][ 362 ],
   alphaCSR[ 158 ][ 363 ],
   alphaCSR[ 158 ][ 364 ],
   alphaCSR[ 158 ][ 365 ],
   alphaCSR[ 158 ][ 366 ],
   alphaCSR[ 158 ][ 367 ],
   alphaCSR[ 158 ][ 368 ],
   alphaCSR[ 158 ][ 369 ],
   alphaCSR[ 158 ][ 370 ],
   alphaCSR[ 158 ][ 371 ],
   alphaCSR[ 158 ][ 372 ],
   alphaCSR[ 158 ][ 373 ],
   alphaCSR[ 158 ][ 374 ],
   alphaCSR[ 158 ][ 375 ],
   alphaCSR[ 158 ][ 376 ],
   alphaCSR[ 158 ][ 377 ],
   alphaCSR[ 158 ][ 378 ],
   alphaCSR[ 158 ][ 379 ],
   alphaCSR[ 158 ][ 380 ],
   alphaCSR[ 158 ][ 381 ],
   alphaCSR[ 158 ][ 382 ],
   alphaCSR[ 158 ][ 383 ],
   alphaCSR[ 159 ][ 0 ],
   alphaCSR[ 159 ][ 1 ],
   alphaCSR[ 159 ][ 2 ],
   alphaCSR[ 159 ][ 3 ],
   alphaCSR[ 159 ][ 4 ],
   alphaCSR[ 159 ][ 5 ],
   alphaCSR[ 159 ][ 6 ],
   alphaCSR[ 159 ][ 7 ],
   alphaCSR[ 159 ][ 8 ],
   alphaCSR[ 159 ][ 9 ],
   alphaCSR[ 159 ][ 10 ],
   alphaCSR[ 159 ][ 11 ],
   alphaCSR[ 159 ][ 12 ],
   alphaCSR[ 159 ][ 13 ],
   alphaCSR[ 159 ][ 14 ],
   alphaCSR[ 159 ][ 15 ],
   alphaCSR[ 159 ][ 16 ],
   alphaCSR[ 159 ][ 17 ],
   alphaCSR[ 159 ][ 18 ],
   alphaCSR[ 159 ][ 19 ],
   alphaCSR[ 159 ][ 20 ],
   alphaCSR[ 159 ][ 21 ],
   alphaCSR[ 159 ][ 22 ],
   alphaCSR[ 159 ][ 23 ],
   alphaCSR[ 159 ][ 24 ],
   alphaCSR[ 159 ][ 25 ],
   alphaCSR[ 159 ][ 26 ],
   alphaCSR[ 159 ][ 27 ],
   alphaCSR[ 159 ][ 28 ],
   alphaCSR[ 159 ][ 29 ],
   alphaCSR[ 159 ][ 30 ],
   alphaCSR[ 159 ][ 31 ],
   alphaCSR[ 159 ][ 32 ],
   alphaCSR[ 159 ][ 33 ],
   alphaCSR[ 159 ][ 34 ],
   alphaCSR[ 159 ][ 35 ],
   alphaCSR[ 159 ][ 36 ],
   alphaCSR[ 159 ][ 37 ],
   alphaCSR[ 159 ][ 38 ],
   alphaCSR[ 159 ][ 39 ],
   alphaCSR[ 159 ][ 40 ],
   alphaCSR[ 159 ][ 41 ],
   alphaCSR[ 159 ][ 42 ],
   alphaCSR[ 159 ][ 43 ],
   alphaCSR[ 159 ][ 44 ],
   alphaCSR[ 159 ][ 45 ],
   alphaCSR[ 159 ][ 46 ],
   alphaCSR[ 159 ][ 47 ],
   alphaCSR[ 159 ][ 48 ],
   alphaCSR[ 159 ][ 49 ],
   alphaCSR[ 159 ][ 50 ],
   alphaCSR[ 159 ][ 51 ],
   alphaCSR[ 159 ][ 52 ],
   alphaCSR[ 159 ][ 53 ],
   alphaCSR[ 159 ][ 54 ],
   alphaCSR[ 159 ][ 55 ],
   alphaCSR[ 159 ][ 56 ],
   alphaCSR[ 159 ][ 57 ],
   alphaCSR[ 159 ][ 58 ],
   alphaCSR[ 159 ][ 59 ],
   alphaCSR[ 159 ][ 60 ],
   alphaCSR[ 159 ][ 61 ],
   alphaCSR[ 159 ][ 62 ],
   alphaCSR[ 159 ][ 63 ],
   alphaCSR[ 159 ][ 64 ],
   alphaCSR[ 159 ][ 65 ],
   alphaCSR[ 159 ][ 66 ],
   alphaCSR[ 159 ][ 67 ],
   alphaCSR[ 159 ][ 68 ],
   alphaCSR[ 159 ][ 69 ],
   alphaCSR[ 159 ][ 70 ],
   alphaCSR[ 159 ][ 71 ],
   alphaCSR[ 159 ][ 72 ],
   alphaCSR[ 159 ][ 73 ],
   alphaCSR[ 159 ][ 74 ],
   alphaCSR[ 159 ][ 75 ],
   alphaCSR[ 159 ][ 76 ],
   alphaCSR[ 159 ][ 77 ],
   alphaCSR[ 159 ][ 78 ],
   alphaCSR[ 159 ][ 79 ],
   alphaCSR[ 159 ][ 80 ],
   alphaCSR[ 159 ][ 81 ],
   alphaCSR[ 159 ][ 82 ],
   alphaCSR[ 159 ][ 83 ],
   alphaCSR[ 159 ][ 84 ],
   alphaCSR[ 159 ][ 85 ],
   alphaCSR[ 159 ][ 86 ],
   alphaCSR[ 159 ][ 87 ],
   alphaCSR[ 159 ][ 88 ],
   alphaCSR[ 159 ][ 89 ],
   alphaCSR[ 159 ][ 90 ],
   alphaCSR[ 159 ][ 91 ],
   alphaCSR[ 159 ][ 92 ],
   alphaCSR[ 159 ][ 93 ],
   alphaCSR[ 159 ][ 94 ],
   alphaCSR[ 159 ][ 95 ],
   alphaCSR[ 159 ][ 96 ],
   alphaCSR[ 159 ][ 97 ],
   alphaCSR[ 159 ][ 98 ],
   alphaCSR[ 159 ][ 99 ],
   alphaCSR[ 159 ][ 100 ],
   alphaCSR[ 159 ][ 101 ],
   alphaCSR[ 159 ][ 102 ],
   alphaCSR[ 159 ][ 103 ],
   alphaCSR[ 159 ][ 104 ],
   alphaCSR[ 159 ][ 105 ],
   alphaCSR[ 159 ][ 106 ],
   alphaCSR[ 159 ][ 107 ],
   alphaCSR[ 159 ][ 108 ],
   alphaCSR[ 159 ][ 109 ],
   alphaCSR[ 159 ][ 110 ],
   alphaCSR[ 159 ][ 111 ],
   alphaCSR[ 159 ][ 112 ],
   alphaCSR[ 159 ][ 113 ],
   alphaCSR[ 159 ][ 114 ],
   alphaCSR[ 159 ][ 115 ],
   alphaCSR[ 159 ][ 116 ],
   alphaCSR[ 159 ][ 117 ],
   alphaCSR[ 159 ][ 118 ],
   alphaCSR[ 159 ][ 119 ],
   alphaCSR[ 159 ][ 120 ],
   alphaCSR[ 159 ][ 121 ],
   alphaCSR[ 159 ][ 122 ],
   alphaCSR[ 159 ][ 123 ],
   alphaCSR[ 159 ][ 124 ],
   alphaCSR[ 159 ][ 125 ],
   alphaCSR[ 159 ][ 126 ],
   alphaCSR[ 159 ][ 127 ],
   alphaCSR[ 159 ][ 128 ],
   alphaCSR[ 159 ][ 129 ],
   alphaCSR[ 159 ][ 130 ],
   alphaCSR[ 159 ][ 131 ],
   alphaCSR[ 159 ][ 132 ],
   alphaCSR[ 159 ][ 133 ],
   alphaCSR[ 159 ][ 134 ],
   alphaCSR[ 159 ][ 135 ],
   alphaCSR[ 159 ][ 136 ],
   alphaCSR[ 159 ][ 137 ],
   alphaCSR[ 159 ][ 138 ],
   alphaCSR[ 159 ][ 139 ],
   alphaCSR[ 159 ][ 140 ],
   alphaCSR[ 159 ][ 141 ],
   alphaCSR[ 159 ][ 142 ],
   alphaCSR[ 159 ][ 143 ],
   alphaCSR[ 159 ][ 144 ],
   alphaCSR[ 159 ][ 145 ],
   alphaCSR[ 159 ][ 146 ],
   alphaCSR[ 159 ][ 147 ],
   alphaCSR[ 159 ][ 148 ],
   alphaCSR[ 159 ][ 149 ],
   alphaCSR[ 159 ][ 150 ],
   alphaCSR[ 159 ][ 151 ],
   alphaCSR[ 159 ][ 152 ],
   alphaCSR[ 159 ][ 153 ],
   alphaCSR[ 159 ][ 154 ],
   alphaCSR[ 159 ][ 155 ],
   alphaCSR[ 159 ][ 156 ],
   alphaCSR[ 159 ][ 157 ],
   alphaCSR[ 159 ][ 158 ],
   alphaCSR[ 159 ][ 159 ],
   alphaCSR[ 159 ][ 160 ],
   alphaCSR[ 159 ][ 161 ],
   alphaCSR[ 159 ][ 162 ],
   alphaCSR[ 159 ][ 163 ],
   alphaCSR[ 159 ][ 164 ],
   alphaCSR[ 159 ][ 165 ],
   alphaCSR[ 159 ][ 166 ],
   alphaCSR[ 159 ][ 167 ],
   alphaCSR[ 159 ][ 168 ],
   alphaCSR[ 159 ][ 169 ],
   alphaCSR[ 159 ][ 170 ],
   alphaCSR[ 159 ][ 171 ],
   alphaCSR[ 159 ][ 172 ],
   alphaCSR[ 159 ][ 173 ],
   alphaCSR[ 159 ][ 174 ],
   alphaCSR[ 159 ][ 175 ],
   alphaCSR[ 159 ][ 176 ],
   alphaCSR[ 159 ][ 177 ],
   alphaCSR[ 159 ][ 178 ],
   alphaCSR[ 159 ][ 179 ],
   alphaCSR[ 159 ][ 180 ],
   alphaCSR[ 159 ][ 181 ],
   alphaCSR[ 159 ][ 182 ],
   alphaCSR[ 159 ][ 183 ],
   alphaCSR[ 159 ][ 184 ],
   alphaCSR[ 159 ][ 185 ],
   alphaCSR[ 159 ][ 186 ],
   alphaCSR[ 159 ][ 187 ],
   alphaCSR[ 159 ][ 188 ],
   alphaCSR[ 159 ][ 189 ],
   alphaCSR[ 159 ][ 190 ],
   alphaCSR[ 159 ][ 191 ],
   alphaCSR[ 159 ][ 192 ],
   alphaCSR[ 159 ][ 193 ],
   alphaCSR[ 159 ][ 194 ],
   alphaCSR[ 159 ][ 195 ],
   alphaCSR[ 159 ][ 196 ],
   alphaCSR[ 159 ][ 197 ],
   alphaCSR[ 159 ][ 198 ],
   alphaCSR[ 159 ][ 199 ],
   alphaCSR[ 159 ][ 200 ],
   alphaCSR[ 159 ][ 201 ],
   alphaCSR[ 159 ][ 202 ],
   alphaCSR[ 159 ][ 203 ],
   alphaCSR[ 159 ][ 204 ],
   alphaCSR[ 159 ][ 205 ],
   alphaCSR[ 159 ][ 206 ],
   alphaCSR[ 159 ][ 207 ],
   alphaCSR[ 159 ][ 208 ],
   alphaCSR[ 159 ][ 209 ],
   alphaCSR[ 159 ][ 210 ],
   alphaCSR[ 159 ][ 211 ],
   alphaCSR[ 159 ][ 212 ],
   alphaCSR[ 159 ][ 213 ],
   alphaCSR[ 159 ][ 214 ],
   alphaCSR[ 159 ][ 215 ],
   alphaCSR[ 159 ][ 216 ],
   alphaCSR[ 159 ][ 217 ],
   alphaCSR[ 159 ][ 218 ],
   alphaCSR[ 159 ][ 219 ],
   alphaCSR[ 159 ][ 220 ],
   alphaCSR[ 159 ][ 221 ],
   alphaCSR[ 159 ][ 222 ],
   alphaCSR[ 159 ][ 223 ],
   alphaCSR[ 159 ][ 224 ],
   alphaCSR[ 159 ][ 225 ],
   alphaCSR[ 159 ][ 226 ],
   alphaCSR[ 159 ][ 227 ],
   alphaCSR[ 159 ][ 228 ],
   alphaCSR[ 159 ][ 229 ],
   alphaCSR[ 159 ][ 230 ],
   alphaCSR[ 159 ][ 231 ],
   alphaCSR[ 159 ][ 232 ],
   alphaCSR[ 159 ][ 233 ],
   alphaCSR[ 159 ][ 234 ],
   alphaCSR[ 159 ][ 235 ],
   alphaCSR[ 159 ][ 236 ],
   alphaCSR[ 159 ][ 237 ],
   alphaCSR[ 159 ][ 238 ],
   alphaCSR[ 159 ][ 239 ],
   alphaCSR[ 159 ][ 240 ],
   alphaCSR[ 159 ][ 241 ],
   alphaCSR[ 159 ][ 242 ],
   alphaCSR[ 159 ][ 243 ],
   alphaCSR[ 159 ][ 244 ],
   alphaCSR[ 159 ][ 245 ],
   alphaCSR[ 159 ][ 246 ],
   alphaCSR[ 159 ][ 247 ],
   alphaCSR[ 159 ][ 248 ],
   alphaCSR[ 159 ][ 249 ],
   alphaCSR[ 159 ][ 250 ],
   alphaCSR[ 159 ][ 251 ],
   alphaCSR[ 159 ][ 252 ],
   alphaCSR[ 159 ][ 253 ],
   alphaCSR[ 159 ][ 254 ],
   alphaCSR[ 159 ][ 255 ],
   alphaCSR[ 159 ][ 256 ],
   alphaCSR[ 159 ][ 257 ],
   alphaCSR[ 159 ][ 258 ],
   alphaCSR[ 159 ][ 259 ],
   alphaCSR[ 159 ][ 260 ],
   alphaCSR[ 159 ][ 261 ],
   alphaCSR[ 159 ][ 262 ],
   alphaCSR[ 159 ][ 263 ],
   alphaCSR[ 159 ][ 264 ],
   alphaCSR[ 159 ][ 265 ],
   alphaCSR[ 159 ][ 266 ],
   alphaCSR[ 159 ][ 267 ],
   alphaCSR[ 159 ][ 268 ],
   alphaCSR[ 159 ][ 269 ],
   alphaCSR[ 159 ][ 270 ],
   alphaCSR[ 159 ][ 271 ],
   alphaCSR[ 159 ][ 272 ],
   alphaCSR[ 159 ][ 273 ],
   alphaCSR[ 159 ][ 274 ],
   alphaCSR[ 159 ][ 275 ],
   alphaCSR[ 159 ][ 276 ],
   alphaCSR[ 159 ][ 277 ],
   alphaCSR[ 159 ][ 278 ],
   alphaCSR[ 159 ][ 279 ],
   alphaCSR[ 159 ][ 280 ],
   alphaCSR[ 159 ][ 281 ],
   alphaCSR[ 159 ][ 282 ],
   alphaCSR[ 159 ][ 283 ],
   alphaCSR[ 159 ][ 284 ],
   alphaCSR[ 159 ][ 285 ],
   alphaCSR[ 159 ][ 286 ],
   alphaCSR[ 159 ][ 287 ],
   alphaCSR[ 159 ][ 288 ],
   alphaCSR[ 159 ][ 289 ],
   alphaCSR[ 159 ][ 290 ],
   alphaCSR[ 159 ][ 291 ],
   alphaCSR[ 159 ][ 292 ],
   alphaCSR[ 159 ][ 293 ],
   alphaCSR[ 159 ][ 294 ],
   alphaCSR[ 159 ][ 295 ],
   alphaCSR[ 159 ][ 296 ],
   alphaCSR[ 159 ][ 297 ],
   alphaCSR[ 159 ][ 298 ],
   alphaCSR[ 159 ][ 299 ],
   alphaCSR[ 159 ][ 300 ],
   alphaCSR[ 159 ][ 301 ],
   alphaCSR[ 159 ][ 302 ],
   alphaCSR[ 159 ][ 303 ],
   alphaCSR[ 159 ][ 304 ],
   alphaCSR[ 159 ][ 305 ],
   alphaCSR[ 159 ][ 306 ],
   alphaCSR[ 159 ][ 307 ],
   alphaCSR[ 159 ][ 308 ],
   alphaCSR[ 159 ][ 309 ],
   alphaCSR[ 159 ][ 310 ],
   alphaCSR[ 159 ][ 311 ],
   alphaCSR[ 159 ][ 312 ],
   alphaCSR[ 159 ][ 313 ],
   alphaCSR[ 159 ][ 314 ],
   alphaCSR[ 159 ][ 315 ],
   alphaCSR[ 159 ][ 316 ],
   alphaCSR[ 159 ][ 317 ],
   alphaCSR[ 159 ][ 318 ],
   alphaCSR[ 159 ][ 319 ],
   alphaCSR[ 159 ][ 320 ],
   alphaCSR[ 159 ][ 321 ],
   alphaCSR[ 159 ][ 322 ],
   alphaCSR[ 159 ][ 323 ],
   alphaCSR[ 159 ][ 324 ],
   alphaCSR[ 159 ][ 325 ],
   alphaCSR[ 159 ][ 326 ],
   alphaCSR[ 159 ][ 327 ],
   alphaCSR[ 159 ][ 328 ],
   alphaCSR[ 159 ][ 329 ],
   alphaCSR[ 159 ][ 330 ],
   alphaCSR[ 159 ][ 331 ],
   alphaCSR[ 159 ][ 332 ],
   alphaCSR[ 159 ][ 333 ],
   alphaCSR[ 159 ][ 334 ],
   alphaCSR[ 159 ][ 335 ],
   alphaCSR[ 159 ][ 336 ],
   alphaCSR[ 159 ][ 337 ],
   alphaCSR[ 159 ][ 338 ],
   alphaCSR[ 159 ][ 339 ],
   alphaCSR[ 159 ][ 340 ],
   alphaCSR[ 159 ][ 341 ],
   alphaCSR[ 159 ][ 342 ],
   alphaCSR[ 159 ][ 343 ],
   alphaCSR[ 159 ][ 344 ],
   alphaCSR[ 159 ][ 345 ],
   alphaCSR[ 159 ][ 346 ],
   alphaCSR[ 159 ][ 347 ],
   alphaCSR[ 159 ][ 348 ],
   alphaCSR[ 159 ][ 349 ],
   alphaCSR[ 159 ][ 350 ],
   alphaCSR[ 159 ][ 351 ],
   alphaCSR[ 159 ][ 352 ],
   alphaCSR[ 159 ][ 353 ],
   alphaCSR[ 159 ][ 354 ],
   alphaCSR[ 159 ][ 355 ],
   alphaCSR[ 159 ][ 356 ],
   alphaCSR[ 159 ][ 357 ],
   alphaCSR[ 159 ][ 358 ],
   alphaCSR[ 159 ][ 359 ],
   alphaCSR[ 159 ][ 360 ],
   alphaCSR[ 159 ][ 361 ],
   alphaCSR[ 159 ][ 362 ],
   alphaCSR[ 159 ][ 363 ],
   alphaCSR[ 159 ][ 364 ],
   alphaCSR[ 159 ][ 365 ],
   alphaCSR[ 159 ][ 366 ],
   alphaCSR[ 159 ][ 367 ],
   alphaCSR[ 159 ][ 368 ],
   alphaCSR[ 159 ][ 369 ],
   alphaCSR[ 159 ][ 370 ],
   alphaCSR[ 159 ][ 371 ],
   alphaCSR[ 159 ][ 372 ],
   alphaCSR[ 159 ][ 373 ],
   alphaCSR[ 159 ][ 374 ],
   alphaCSR[ 159 ][ 375 ],
   alphaCSR[ 159 ][ 376 ],
   alphaCSR[ 159 ][ 377 ],
   alphaCSR[ 159 ][ 378 ],
   alphaCSR[ 159 ][ 379 ],
   alphaCSR[ 159 ][ 380 ],
   alphaCSR[ 159 ][ 381 ],
   alphaCSR[ 159 ][ 382 ],
   alphaCSR[ 159 ][ 383 ],
   alphaCSR[ 160 ][ 0 ],
   alphaCSR[ 160 ][ 1 ],
   alphaCSR[ 160 ][ 2 ],
   alphaCSR[ 160 ][ 3 ],
   alphaCSR[ 160 ][ 4 ],
   alphaCSR[ 160 ][ 5 ],
   alphaCSR[ 160 ][ 6 ],
   alphaCSR[ 160 ][ 7 ],
   alphaCSR[ 160 ][ 8 ],
   alphaCSR[ 160 ][ 9 ],
   alphaCSR[ 160 ][ 10 ],
   alphaCSR[ 160 ][ 11 ],
   alphaCSR[ 160 ][ 12 ],
   alphaCSR[ 160 ][ 13 ],
   alphaCSR[ 160 ][ 14 ],
   alphaCSR[ 160 ][ 15 ],
   alphaCSR[ 160 ][ 16 ],
   alphaCSR[ 160 ][ 17 ],
   alphaCSR[ 160 ][ 18 ],
   alphaCSR[ 160 ][ 19 ],
   alphaCSR[ 160 ][ 20 ],
   alphaCSR[ 160 ][ 21 ],
   alphaCSR[ 160 ][ 22 ],
   alphaCSR[ 160 ][ 23 ],
   alphaCSR[ 160 ][ 24 ],
   alphaCSR[ 160 ][ 25 ],
   alphaCSR[ 160 ][ 26 ],
   alphaCSR[ 160 ][ 27 ],
   alphaCSR[ 160 ][ 28 ],
   alphaCSR[ 160 ][ 29 ],
   alphaCSR[ 160 ][ 30 ],
   alphaCSR[ 160 ][ 31 ],
   alphaCSR[ 160 ][ 32 ],
   alphaCSR[ 160 ][ 33 ],
   alphaCSR[ 160 ][ 34 ],
   alphaCSR[ 160 ][ 35 ],
   alphaCSR[ 160 ][ 36 ],
   alphaCSR[ 160 ][ 37 ],
   alphaCSR[ 160 ][ 38 ],
   alphaCSR[ 160 ][ 39 ],
   alphaCSR[ 160 ][ 40 ],
   alphaCSR[ 160 ][ 41 ],
   alphaCSR[ 160 ][ 42 ],
   alphaCSR[ 160 ][ 43 ],
   alphaCSR[ 160 ][ 44 ],
   alphaCSR[ 160 ][ 45 ],
   alphaCSR[ 160 ][ 46 ],
   alphaCSR[ 160 ][ 47 ],
   alphaCSR[ 160 ][ 48 ],
   alphaCSR[ 160 ][ 49 ],
   alphaCSR[ 160 ][ 50 ],
   alphaCSR[ 160 ][ 51 ],
   alphaCSR[ 160 ][ 52 ],
   alphaCSR[ 160 ][ 53 ],
   alphaCSR[ 160 ][ 54 ],
   alphaCSR[ 160 ][ 55 ],
   alphaCSR[ 160 ][ 56 ],
   alphaCSR[ 160 ][ 57 ],
   alphaCSR[ 160 ][ 58 ],
   alphaCSR[ 160 ][ 59 ],
   alphaCSR[ 160 ][ 60 ],
   alphaCSR[ 160 ][ 61 ],
   alphaCSR[ 160 ][ 62 ],
   alphaCSR[ 160 ][ 63 ],
   alphaCSR[ 160 ][ 64 ],
   alphaCSR[ 160 ][ 65 ],
   alphaCSR[ 160 ][ 66 ],
   alphaCSR[ 160 ][ 67 ],
   alphaCSR[ 160 ][ 68 ],
   alphaCSR[ 160 ][ 69 ],
   alphaCSR[ 160 ][ 70 ],
   alphaCSR[ 160 ][ 71 ],
   alphaCSR[ 160 ][ 72 ],
   alphaCSR[ 160 ][ 73 ],
   alphaCSR[ 160 ][ 74 ],
   alphaCSR[ 160 ][ 75 ],
   alphaCSR[ 160 ][ 76 ],
   alphaCSR[ 160 ][ 77 ],
   alphaCSR[ 160 ][ 78 ],
   alphaCSR[ 160 ][ 79 ],
   alphaCSR[ 160 ][ 80 ],
   alphaCSR[ 160 ][ 81 ],
   alphaCSR[ 160 ][ 82 ],
   alphaCSR[ 160 ][ 83 ],
   alphaCSR[ 160 ][ 84 ],
   alphaCSR[ 160 ][ 85 ],
   alphaCSR[ 160 ][ 86 ],
   alphaCSR[ 160 ][ 87 ],
   alphaCSR[ 160 ][ 88 ],
   alphaCSR[ 160 ][ 89 ],
   alphaCSR[ 160 ][ 90 ],
   alphaCSR[ 160 ][ 91 ],
   alphaCSR[ 160 ][ 92 ],
   alphaCSR[ 160 ][ 93 ],
   alphaCSR[ 160 ][ 94 ],
   alphaCSR[ 160 ][ 95 ],
   alphaCSR[ 160 ][ 96 ],
   alphaCSR[ 160 ][ 97 ],
   alphaCSR[ 160 ][ 98 ],
   alphaCSR[ 160 ][ 99 ],
   alphaCSR[ 160 ][ 100 ],
   alphaCSR[ 160 ][ 101 ],
   alphaCSR[ 160 ][ 102 ],
   alphaCSR[ 160 ][ 103 ],
   alphaCSR[ 160 ][ 104 ],
   alphaCSR[ 160 ][ 105 ],
   alphaCSR[ 160 ][ 106 ],
   alphaCSR[ 160 ][ 107 ],
   alphaCSR[ 160 ][ 108 ],
   alphaCSR[ 160 ][ 109 ],
   alphaCSR[ 160 ][ 110 ],
   alphaCSR[ 160 ][ 111 ],
   alphaCSR[ 160 ][ 112 ],
   alphaCSR[ 160 ][ 113 ],
   alphaCSR[ 160 ][ 114 ],
   alphaCSR[ 160 ][ 115 ],
   alphaCSR[ 160 ][ 116 ],
   alphaCSR[ 160 ][ 117 ],
   alphaCSR[ 160 ][ 118 ],
   alphaCSR[ 160 ][ 119 ],
   alphaCSR[ 160 ][ 120 ],
   alphaCSR[ 160 ][ 121 ],
   alphaCSR[ 160 ][ 122 ],
   alphaCSR[ 160 ][ 123 ],
   alphaCSR[ 160 ][ 124 ],
   alphaCSR[ 160 ][ 125 ],
   alphaCSR[ 160 ][ 126 ],
   alphaCSR[ 160 ][ 127 ],
   alphaCSR[ 160 ][ 128 ],
   alphaCSR[ 160 ][ 129 ],
   alphaCSR[ 160 ][ 130 ],
   alphaCSR[ 160 ][ 131 ],
   alphaCSR[ 160 ][ 132 ],
   alphaCSR[ 160 ][ 133 ],
   alphaCSR[ 160 ][ 134 ],
   alphaCSR[ 160 ][ 135 ],
   alphaCSR[ 160 ][ 136 ],
   alphaCSR[ 160 ][ 137 ],
   alphaCSR[ 160 ][ 138 ],
   alphaCSR[ 160 ][ 139 ],
   alphaCSR[ 160 ][ 140 ],
   alphaCSR[ 160 ][ 141 ],
   alphaCSR[ 160 ][ 142 ],
   alphaCSR[ 160 ][ 143 ],
   alphaCSR[ 160 ][ 144 ],
   alphaCSR[ 160 ][ 145 ],
   alphaCSR[ 160 ][ 146 ],
   alphaCSR[ 160 ][ 147 ],
   alphaCSR[ 160 ][ 148 ],
   alphaCSR[ 160 ][ 149 ],
   alphaCSR[ 160 ][ 150 ],
   alphaCSR[ 160 ][ 151 ],
   alphaCSR[ 160 ][ 152 ],
   alphaCSR[ 160 ][ 153 ],
   alphaCSR[ 160 ][ 154 ],
   alphaCSR[ 160 ][ 155 ],
   alphaCSR[ 160 ][ 156 ],
   alphaCSR[ 160 ][ 157 ],
   alphaCSR[ 160 ][ 158 ],
   alphaCSR[ 160 ][ 159 ],
   alphaCSR[ 160 ][ 160 ],
   alphaCSR[ 160 ][ 161 ],
   alphaCSR[ 160 ][ 162 ],
   alphaCSR[ 160 ][ 163 ],
   alphaCSR[ 160 ][ 164 ],
   alphaCSR[ 160 ][ 165 ],
   alphaCSR[ 160 ][ 166 ],
   alphaCSR[ 160 ][ 167 ],
   alphaCSR[ 160 ][ 168 ],
   alphaCSR[ 160 ][ 169 ],
   alphaCSR[ 160 ][ 170 ],
   alphaCSR[ 160 ][ 171 ],
   alphaCSR[ 160 ][ 172 ],
   alphaCSR[ 160 ][ 173 ],
   alphaCSR[ 160 ][ 174 ],
   alphaCSR[ 160 ][ 175 ],
   alphaCSR[ 160 ][ 176 ],
   alphaCSR[ 160 ][ 177 ],
   alphaCSR[ 160 ][ 178 ],
   alphaCSR[ 160 ][ 179 ],
   alphaCSR[ 160 ][ 180 ],
   alphaCSR[ 160 ][ 181 ],
   alphaCSR[ 160 ][ 182 ],
   alphaCSR[ 160 ][ 183 ],
   alphaCSR[ 160 ][ 184 ],
   alphaCSR[ 160 ][ 185 ],
   alphaCSR[ 160 ][ 186 ],
   alphaCSR[ 160 ][ 187 ],
   alphaCSR[ 160 ][ 188 ],
   alphaCSR[ 160 ][ 189 ],
   alphaCSR[ 160 ][ 190 ],
   alphaCSR[ 160 ][ 191 ],
   alphaCSR[ 160 ][ 192 ],
   alphaCSR[ 160 ][ 193 ],
   alphaCSR[ 160 ][ 194 ],
   alphaCSR[ 160 ][ 195 ],
   alphaCSR[ 160 ][ 196 ],
   alphaCSR[ 160 ][ 197 ],
   alphaCSR[ 160 ][ 198 ],
   alphaCSR[ 160 ][ 199 ],
   alphaCSR[ 160 ][ 200 ],
   alphaCSR[ 160 ][ 201 ],
   alphaCSR[ 160 ][ 202 ],
   alphaCSR[ 160 ][ 203 ],
   alphaCSR[ 160 ][ 204 ],
   alphaCSR[ 160 ][ 205 ],
   alphaCSR[ 160 ][ 206 ],
   alphaCSR[ 160 ][ 207 ],
   alphaCSR[ 160 ][ 208 ],
   alphaCSR[ 160 ][ 209 ],
   alphaCSR[ 160 ][ 210 ],
   alphaCSR[ 160 ][ 211 ],
   alphaCSR[ 160 ][ 212 ],
   alphaCSR[ 160 ][ 213 ],
   alphaCSR[ 160 ][ 214 ],
   alphaCSR[ 160 ][ 215 ],
   alphaCSR[ 160 ][ 216 ],
   alphaCSR[ 160 ][ 217 ],
   alphaCSR[ 160 ][ 218 ],
   alphaCSR[ 160 ][ 219 ],
   alphaCSR[ 160 ][ 220 ],
   alphaCSR[ 160 ][ 221 ],
   alphaCSR[ 160 ][ 222 ],
   alphaCSR[ 160 ][ 223 ],
   alphaCSR[ 160 ][ 224 ],
   alphaCSR[ 160 ][ 225 ],
   alphaCSR[ 160 ][ 226 ],
   alphaCSR[ 160 ][ 227 ],
   alphaCSR[ 160 ][ 228 ],
   alphaCSR[ 160 ][ 229 ],
   alphaCSR[ 160 ][ 230 ],
   alphaCSR[ 160 ][ 231 ],
   alphaCSR[ 160 ][ 232 ],
   alphaCSR[ 160 ][ 233 ],
   alphaCSR[ 160 ][ 234 ],
   alphaCSR[ 160 ][ 235 ],
   alphaCSR[ 160 ][ 236 ],
   alphaCSR[ 160 ][ 237 ],
   alphaCSR[ 160 ][ 238 ],
   alphaCSR[ 160 ][ 239 ],
   alphaCSR[ 160 ][ 240 ],
   alphaCSR[ 160 ][ 241 ],
   alphaCSR[ 160 ][ 242 ],
   alphaCSR[ 160 ][ 243 ],
   alphaCSR[ 160 ][ 244 ],
   alphaCSR[ 160 ][ 245 ],
   alphaCSR[ 160 ][ 246 ],
   alphaCSR[ 160 ][ 247 ],
   alphaCSR[ 160 ][ 248 ],
   alphaCSR[ 160 ][ 249 ],
   alphaCSR[ 160 ][ 250 ],
   alphaCSR[ 160 ][ 251 ],
   alphaCSR[ 160 ][ 252 ],
   alphaCSR[ 160 ][ 253 ],
   alphaCSR[ 160 ][ 254 ],
   alphaCSR[ 160 ][ 255 ],
   alphaCSR[ 160 ][ 256 ],
   alphaCSR[ 160 ][ 257 ],
   alphaCSR[ 160 ][ 258 ],
   alphaCSR[ 160 ][ 259 ],
   alphaCSR[ 160 ][ 260 ],
   alphaCSR[ 160 ][ 261 ],
   alphaCSR[ 160 ][ 262 ],
   alphaCSR[ 160 ][ 263 ],
   alphaCSR[ 160 ][ 264 ],
   alphaCSR[ 160 ][ 265 ],
   alphaCSR[ 160 ][ 266 ],
   alphaCSR[ 160 ][ 267 ],
   alphaCSR[ 160 ][ 268 ],
   alphaCSR[ 160 ][ 269 ],
   alphaCSR[ 160 ][ 270 ],
   alphaCSR[ 160 ][ 271 ],
   alphaCSR[ 160 ][ 272 ],
   alphaCSR[ 160 ][ 273 ],
   alphaCSR[ 160 ][ 274 ],
   alphaCSR[ 160 ][ 275 ],
   alphaCSR[ 160 ][ 276 ],
   alphaCSR[ 160 ][ 277 ],
   alphaCSR[ 160 ][ 278 ],
   alphaCSR[ 160 ][ 279 ],
   alphaCSR[ 160 ][ 280 ],
   alphaCSR[ 160 ][ 281 ],
   alphaCSR[ 160 ][ 282 ],
   alphaCSR[ 160 ][ 283 ],
   alphaCSR[ 160 ][ 284 ],
   alphaCSR[ 160 ][ 285 ],
   alphaCSR[ 160 ][ 286 ],
   alphaCSR[ 160 ][ 287 ],
   alphaCSR[ 160 ][ 288 ],
   alphaCSR[ 160 ][ 289 ],
   alphaCSR[ 160 ][ 290 ],
   alphaCSR[ 160 ][ 291 ],
   alphaCSR[ 160 ][ 292 ],
   alphaCSR[ 160 ][ 293 ],
   alphaCSR[ 160 ][ 294 ],
   alphaCSR[ 160 ][ 295 ],
   alphaCSR[ 160 ][ 296 ],
   alphaCSR[ 160 ][ 297 ],
   alphaCSR[ 160 ][ 298 ],
   alphaCSR[ 160 ][ 299 ],
   alphaCSR[ 160 ][ 300 ],
   alphaCSR[ 160 ][ 301 ],
   alphaCSR[ 160 ][ 302 ],
   alphaCSR[ 160 ][ 303 ],
   alphaCSR[ 160 ][ 304 ],
   alphaCSR[ 160 ][ 305 ],
   alphaCSR[ 160 ][ 306 ],
   alphaCSR[ 160 ][ 307 ],
   alphaCSR[ 160 ][ 308 ],
   alphaCSR[ 160 ][ 309 ],
   alphaCSR[ 160 ][ 310 ],
   alphaCSR[ 160 ][ 311 ],
   alphaCSR[ 160 ][ 312 ],
   alphaCSR[ 160 ][ 313 ],
   alphaCSR[ 160 ][ 314 ],
   alphaCSR[ 160 ][ 315 ],
   alphaCSR[ 160 ][ 316 ],
   alphaCSR[ 160 ][ 317 ],
   alphaCSR[ 160 ][ 318 ],
   alphaCSR[ 160 ][ 319 ],
   alphaCSR[ 160 ][ 320 ],
   alphaCSR[ 160 ][ 321 ],
   alphaCSR[ 160 ][ 322 ],
   alphaCSR[ 160 ][ 323 ],
   alphaCSR[ 160 ][ 324 ],
   alphaCSR[ 160 ][ 325 ],
   alphaCSR[ 160 ][ 326 ],
   alphaCSR[ 160 ][ 327 ],
   alphaCSR[ 160 ][ 328 ],
   alphaCSR[ 160 ][ 329 ],
   alphaCSR[ 160 ][ 330 ],
   alphaCSR[ 160 ][ 331 ],
   alphaCSR[ 160 ][ 332 ],
   alphaCSR[ 160 ][ 333 ],
   alphaCSR[ 160 ][ 334 ],
   alphaCSR[ 160 ][ 335 ],
   alphaCSR[ 160 ][ 336 ],
   alphaCSR[ 160 ][ 337 ],
   alphaCSR[ 160 ][ 338 ],
   alphaCSR[ 160 ][ 339 ],
   alphaCSR[ 160 ][ 340 ],
   alphaCSR[ 160 ][ 341 ],
   alphaCSR[ 160 ][ 342 ],
   alphaCSR[ 160 ][ 343 ],
   alphaCSR[ 160 ][ 344 ],
   alphaCSR[ 160 ][ 345 ],
   alphaCSR[ 160 ][ 346 ],
   alphaCSR[ 160 ][ 347 ],
   alphaCSR[ 160 ][ 348 ],
   alphaCSR[ 160 ][ 349 ],
   alphaCSR[ 160 ][ 350 ],
   alphaCSR[ 160 ][ 351 ],
   alphaCSR[ 160 ][ 352 ],
   alphaCSR[ 160 ][ 353 ],
   alphaCSR[ 160 ][ 354 ],
   alphaCSR[ 160 ][ 355 ],
   alphaCSR[ 160 ][ 356 ],
   alphaCSR[ 160 ][ 357 ],
   alphaCSR[ 160 ][ 358 ],
   alphaCSR[ 160 ][ 359 ],
   alphaCSR[ 160 ][ 360 ],
   alphaCSR[ 160 ][ 361 ],
   alphaCSR[ 160 ][ 362 ],
   alphaCSR[ 160 ][ 363 ],
   alphaCSR[ 160 ][ 364 ],
   alphaCSR[ 160 ][ 365 ],
   alphaCSR[ 160 ][ 366 ],
   alphaCSR[ 160 ][ 367 ],
   alphaCSR[ 160 ][ 368 ],
   alphaCSR[ 160 ][ 369 ],
   alphaCSR[ 160 ][ 370 ],
   alphaCSR[ 160 ][ 371 ],
   alphaCSR[ 160 ][ 372 ],
   alphaCSR[ 160 ][ 373 ],
   alphaCSR[ 160 ][ 374 ],
   alphaCSR[ 160 ][ 375 ],
   alphaCSR[ 160 ][ 376 ],
   alphaCSR[ 160 ][ 377 ],
   alphaCSR[ 160 ][ 378 ],
   alphaCSR[ 160 ][ 379 ],
   alphaCSR[ 160 ][ 380 ],
   alphaCSR[ 160 ][ 381 ],
   alphaCSR[ 160 ][ 382 ],
   alphaCSR[ 160 ][ 383 ],
   alphaCSR[ 161 ][ 0 ],
   alphaCSR[ 161 ][ 1 ],
   alphaCSR[ 161 ][ 2 ],
   alphaCSR[ 161 ][ 3 ],
   alphaCSR[ 161 ][ 4 ],
   alphaCSR[ 161 ][ 5 ],
   alphaCSR[ 161 ][ 6 ],
   alphaCSR[ 161 ][ 7 ],
   alphaCSR[ 161 ][ 8 ],
   alphaCSR[ 161 ][ 9 ],
   alphaCSR[ 161 ][ 10 ],
   alphaCSR[ 161 ][ 11 ],
   alphaCSR[ 161 ][ 12 ],
   alphaCSR[ 161 ][ 13 ],
   alphaCSR[ 161 ][ 14 ],
   alphaCSR[ 161 ][ 15 ],
   alphaCSR[ 161 ][ 16 ],
   alphaCSR[ 161 ][ 17 ],
   alphaCSR[ 161 ][ 18 ],
   alphaCSR[ 161 ][ 19 ],
   alphaCSR[ 161 ][ 20 ],
   alphaCSR[ 161 ][ 21 ],
   alphaCSR[ 161 ][ 22 ],
   alphaCSR[ 161 ][ 23 ],
   alphaCSR[ 161 ][ 24 ],
   alphaCSR[ 161 ][ 25 ],
   alphaCSR[ 161 ][ 26 ],
   alphaCSR[ 161 ][ 27 ],
   alphaCSR[ 161 ][ 28 ],
   alphaCSR[ 161 ][ 29 ],
   alphaCSR[ 161 ][ 30 ],
   alphaCSR[ 161 ][ 31 ],
   alphaCSR[ 161 ][ 32 ],
   alphaCSR[ 161 ][ 33 ],
   alphaCSR[ 161 ][ 34 ],
   alphaCSR[ 161 ][ 35 ],
   alphaCSR[ 161 ][ 36 ],
   alphaCSR[ 161 ][ 37 ],
   alphaCSR[ 161 ][ 38 ],
   alphaCSR[ 161 ][ 39 ],
   alphaCSR[ 161 ][ 40 ],
   alphaCSR[ 161 ][ 41 ],
   alphaCSR[ 161 ][ 42 ],
   alphaCSR[ 161 ][ 43 ],
   alphaCSR[ 161 ][ 44 ],
   alphaCSR[ 161 ][ 45 ],
   alphaCSR[ 161 ][ 46 ],
   alphaCSR[ 161 ][ 47 ],
   alphaCSR[ 161 ][ 48 ],
   alphaCSR[ 161 ][ 49 ],
   alphaCSR[ 161 ][ 50 ],
   alphaCSR[ 161 ][ 51 ],
   alphaCSR[ 161 ][ 52 ],
   alphaCSR[ 161 ][ 53 ],
   alphaCSR[ 161 ][ 54 ],
   alphaCSR[ 161 ][ 55 ],
   alphaCSR[ 161 ][ 56 ],
   alphaCSR[ 161 ][ 57 ],
   alphaCSR[ 161 ][ 58 ],
   alphaCSR[ 161 ][ 59 ],
   alphaCSR[ 161 ][ 60 ],
   alphaCSR[ 161 ][ 61 ],
   alphaCSR[ 161 ][ 62 ],
   alphaCSR[ 161 ][ 63 ],
   alphaCSR[ 161 ][ 64 ],
   alphaCSR[ 161 ][ 65 ],
   alphaCSR[ 161 ][ 66 ],
   alphaCSR[ 161 ][ 67 ],
   alphaCSR[ 161 ][ 68 ],
   alphaCSR[ 161 ][ 69 ],
   alphaCSR[ 161 ][ 70 ],
   alphaCSR[ 161 ][ 71 ],
   alphaCSR[ 161 ][ 72 ],
   alphaCSR[ 161 ][ 73 ],
   alphaCSR[ 161 ][ 74 ],
   alphaCSR[ 161 ][ 75 ],
   alphaCSR[ 161 ][ 76 ],
   alphaCSR[ 161 ][ 77 ],
   alphaCSR[ 161 ][ 78 ],
   alphaCSR[ 161 ][ 79 ],
   alphaCSR[ 161 ][ 80 ],
   alphaCSR[ 161 ][ 81 ],
   alphaCSR[ 161 ][ 82 ],
   alphaCSR[ 161 ][ 83 ],
   alphaCSR[ 161 ][ 84 ],
   alphaCSR[ 161 ][ 85 ],
   alphaCSR[ 161 ][ 86 ],
   alphaCSR[ 161 ][ 87 ],
   alphaCSR[ 161 ][ 88 ],
   alphaCSR[ 161 ][ 89 ],
   alphaCSR[ 161 ][ 90 ],
   alphaCSR[ 161 ][ 91 ],
   alphaCSR[ 161 ][ 92 ],
   alphaCSR[ 161 ][ 93 ],
   alphaCSR[ 161 ][ 94 ],
   alphaCSR[ 161 ][ 95 ],
   alphaCSR[ 161 ][ 96 ],
   alphaCSR[ 161 ][ 97 ],
   alphaCSR[ 161 ][ 98 ],
   alphaCSR[ 161 ][ 99 ],
   alphaCSR[ 161 ][ 100 ],
   alphaCSR[ 161 ][ 101 ],
   alphaCSR[ 161 ][ 102 ],
   alphaCSR[ 161 ][ 103 ],
   alphaCSR[ 161 ][ 104 ],
   alphaCSR[ 161 ][ 105 ],
   alphaCSR[ 161 ][ 106 ],
   alphaCSR[ 161 ][ 107 ],
   alphaCSR[ 161 ][ 108 ],
   alphaCSR[ 161 ][ 109 ],
   alphaCSR[ 161 ][ 110 ],
   alphaCSR[ 161 ][ 111 ],
   alphaCSR[ 161 ][ 112 ],
   alphaCSR[ 161 ][ 113 ],
   alphaCSR[ 161 ][ 114 ],
   alphaCSR[ 161 ][ 115 ],
   alphaCSR[ 161 ][ 116 ],
   alphaCSR[ 161 ][ 117 ],
   alphaCSR[ 161 ][ 118 ],
   alphaCSR[ 161 ][ 119 ],
   alphaCSR[ 161 ][ 120 ],
   alphaCSR[ 161 ][ 121 ],
   alphaCSR[ 161 ][ 122 ],
   alphaCSR[ 161 ][ 123 ],
   alphaCSR[ 161 ][ 124 ],
   alphaCSR[ 161 ][ 125 ],
   alphaCSR[ 161 ][ 126 ],
   alphaCSR[ 161 ][ 127 ],
   alphaCSR[ 161 ][ 128 ],
   alphaCSR[ 161 ][ 129 ],
   alphaCSR[ 161 ][ 130 ],
   alphaCSR[ 161 ][ 131 ],
   alphaCSR[ 161 ][ 132 ],
   alphaCSR[ 161 ][ 133 ],
   alphaCSR[ 161 ][ 134 ],
   alphaCSR[ 161 ][ 135 ],
   alphaCSR[ 161 ][ 136 ],
   alphaCSR[ 161 ][ 137 ],
   alphaCSR[ 161 ][ 138 ],
   alphaCSR[ 161 ][ 139 ],
   alphaCSR[ 161 ][ 140 ],
   alphaCSR[ 161 ][ 141 ],
   alphaCSR[ 161 ][ 142 ],
   alphaCSR[ 161 ][ 143 ],
   alphaCSR[ 161 ][ 144 ],
   alphaCSR[ 161 ][ 145 ],
   alphaCSR[ 161 ][ 146 ],
   alphaCSR[ 161 ][ 147 ],
   alphaCSR[ 161 ][ 148 ],
   alphaCSR[ 161 ][ 149 ],
   alphaCSR[ 161 ][ 150 ],
   alphaCSR[ 161 ][ 151 ],
   alphaCSR[ 161 ][ 152 ],
   alphaCSR[ 161 ][ 153 ],
   alphaCSR[ 161 ][ 154 ],
   alphaCSR[ 161 ][ 155 ],
   alphaCSR[ 161 ][ 156 ],
   alphaCSR[ 161 ][ 157 ],
   alphaCSR[ 161 ][ 158 ],
   alphaCSR[ 161 ][ 159 ],
   alphaCSR[ 161 ][ 160 ],
   alphaCSR[ 161 ][ 161 ],
   alphaCSR[ 161 ][ 162 ],
   alphaCSR[ 161 ][ 163 ],
   alphaCSR[ 161 ][ 164 ],
   alphaCSR[ 161 ][ 165 ],
   alphaCSR[ 161 ][ 166 ],
   alphaCSR[ 161 ][ 167 ],
   alphaCSR[ 161 ][ 168 ],
   alphaCSR[ 161 ][ 169 ],
   alphaCSR[ 161 ][ 170 ],
   alphaCSR[ 161 ][ 171 ],
   alphaCSR[ 161 ][ 172 ],
   alphaCSR[ 161 ][ 173 ],
   alphaCSR[ 161 ][ 174 ],
   alphaCSR[ 161 ][ 175 ],
   alphaCSR[ 161 ][ 176 ],
   alphaCSR[ 161 ][ 177 ],
   alphaCSR[ 161 ][ 178 ],
   alphaCSR[ 161 ][ 179 ],
   alphaCSR[ 161 ][ 180 ],
   alphaCSR[ 161 ][ 181 ],
   alphaCSR[ 161 ][ 182 ],
   alphaCSR[ 161 ][ 183 ],
   alphaCSR[ 161 ][ 184 ],
   alphaCSR[ 161 ][ 185 ],
   alphaCSR[ 161 ][ 186 ],
   alphaCSR[ 161 ][ 187 ],
   alphaCSR[ 161 ][ 188 ],
   alphaCSR[ 161 ][ 189 ],
   alphaCSR[ 161 ][ 190 ],
   alphaCSR[ 161 ][ 191 ],
   alphaCSR[ 161 ][ 192 ],
   alphaCSR[ 161 ][ 193 ],
   alphaCSR[ 161 ][ 194 ],
   alphaCSR[ 161 ][ 195 ],
   alphaCSR[ 161 ][ 196 ],
   alphaCSR[ 161 ][ 197 ],
   alphaCSR[ 161 ][ 198 ],
   alphaCSR[ 161 ][ 199 ],
   alphaCSR[ 161 ][ 200 ],
   alphaCSR[ 161 ][ 201 ],
   alphaCSR[ 161 ][ 202 ],
   alphaCSR[ 161 ][ 203 ],
   alphaCSR[ 161 ][ 204 ],
   alphaCSR[ 161 ][ 205 ],
   alphaCSR[ 161 ][ 206 ],
   alphaCSR[ 161 ][ 207 ],
   alphaCSR[ 161 ][ 208 ],
   alphaCSR[ 161 ][ 209 ],
   alphaCSR[ 161 ][ 210 ],
   alphaCSR[ 161 ][ 211 ],
   alphaCSR[ 161 ][ 212 ],
   alphaCSR[ 161 ][ 213 ],
   alphaCSR[ 161 ][ 214 ],
   alphaCSR[ 161 ][ 215 ],
   alphaCSR[ 161 ][ 216 ],
   alphaCSR[ 161 ][ 217 ],
   alphaCSR[ 161 ][ 218 ],
   alphaCSR[ 161 ][ 219 ],
   alphaCSR[ 161 ][ 220 ],
   alphaCSR[ 161 ][ 221 ],
   alphaCSR[ 161 ][ 222 ],
   alphaCSR[ 161 ][ 223 ],
   alphaCSR[ 161 ][ 224 ],
   alphaCSR[ 161 ][ 225 ],
   alphaCSR[ 161 ][ 226 ],
   alphaCSR[ 161 ][ 227 ],
   alphaCSR[ 161 ][ 228 ],
   alphaCSR[ 161 ][ 229 ],
   alphaCSR[ 161 ][ 230 ],
   alphaCSR[ 161 ][ 231 ],
   alphaCSR[ 161 ][ 232 ],
   alphaCSR[ 161 ][ 233 ],
   alphaCSR[ 161 ][ 234 ],
   alphaCSR[ 161 ][ 235 ],
   alphaCSR[ 161 ][ 236 ],
   alphaCSR[ 161 ][ 237 ],
   alphaCSR[ 161 ][ 238 ],
   alphaCSR[ 161 ][ 239 ],
   alphaCSR[ 161 ][ 240 ],
   alphaCSR[ 161 ][ 241 ],
   alphaCSR[ 161 ][ 242 ],
   alphaCSR[ 161 ][ 243 ],
   alphaCSR[ 161 ][ 244 ],
   alphaCSR[ 161 ][ 245 ],
   alphaCSR[ 161 ][ 246 ],
   alphaCSR[ 161 ][ 247 ],
   alphaCSR[ 161 ][ 248 ],
   alphaCSR[ 161 ][ 249 ],
   alphaCSR[ 161 ][ 250 ],
   alphaCSR[ 161 ][ 251 ],
   alphaCSR[ 161 ][ 252 ],
   alphaCSR[ 161 ][ 253 ],
   alphaCSR[ 161 ][ 254 ],
   alphaCSR[ 161 ][ 255 ],
   alphaCSR[ 161 ][ 256 ],
   alphaCSR[ 161 ][ 257 ],
   alphaCSR[ 161 ][ 258 ],
   alphaCSR[ 161 ][ 259 ],
   alphaCSR[ 161 ][ 260 ],
   alphaCSR[ 161 ][ 261 ],
   alphaCSR[ 161 ][ 262 ],
   alphaCSR[ 161 ][ 263 ],
   alphaCSR[ 161 ][ 264 ],
   alphaCSR[ 161 ][ 265 ],
   alphaCSR[ 161 ][ 266 ],
   alphaCSR[ 161 ][ 267 ],
   alphaCSR[ 161 ][ 268 ],
   alphaCSR[ 161 ][ 269 ],
   alphaCSR[ 161 ][ 270 ],
   alphaCSR[ 161 ][ 271 ],
   alphaCSR[ 161 ][ 272 ],
   alphaCSR[ 161 ][ 273 ],
   alphaCSR[ 161 ][ 274 ],
   alphaCSR[ 161 ][ 275 ],
   alphaCSR[ 161 ][ 276 ],
   alphaCSR[ 161 ][ 277 ],
   alphaCSR[ 161 ][ 278 ],
   alphaCSR[ 161 ][ 279 ],
   alphaCSR[ 161 ][ 280 ],
   alphaCSR[ 161 ][ 281 ],
   alphaCSR[ 161 ][ 282 ],
   alphaCSR[ 161 ][ 283 ],
   alphaCSR[ 161 ][ 284 ],
   alphaCSR[ 161 ][ 285 ],
   alphaCSR[ 161 ][ 286 ],
   alphaCSR[ 161 ][ 287 ],
   alphaCSR[ 161 ][ 288 ],
   alphaCSR[ 161 ][ 289 ],
   alphaCSR[ 161 ][ 290 ],
   alphaCSR[ 161 ][ 291 ],
   alphaCSR[ 161 ][ 292 ],
   alphaCSR[ 161 ][ 293 ],
   alphaCSR[ 161 ][ 294 ],
   alphaCSR[ 161 ][ 295 ],
   alphaCSR[ 161 ][ 296 ],
   alphaCSR[ 161 ][ 297 ],
   alphaCSR[ 161 ][ 298 ],
   alphaCSR[ 161 ][ 299 ],
   alphaCSR[ 161 ][ 300 ],
   alphaCSR[ 161 ][ 301 ],
   alphaCSR[ 161 ][ 302 ],
   alphaCSR[ 161 ][ 303 ],
   alphaCSR[ 161 ][ 304 ],
   alphaCSR[ 161 ][ 305 ],
   alphaCSR[ 161 ][ 306 ],
   alphaCSR[ 161 ][ 307 ],
   alphaCSR[ 161 ][ 308 ],
   alphaCSR[ 161 ][ 309 ],
   alphaCSR[ 161 ][ 310 ],
   alphaCSR[ 161 ][ 311 ],
   alphaCSR[ 161 ][ 312 ],
   alphaCSR[ 161 ][ 313 ],
   alphaCSR[ 161 ][ 314 ],
   alphaCSR[ 161 ][ 315 ],
   alphaCSR[ 161 ][ 316 ],
   alphaCSR[ 161 ][ 317 ],
   alphaCSR[ 161 ][ 318 ],
   alphaCSR[ 161 ][ 319 ],
   alphaCSR[ 161 ][ 320 ],
   alphaCSR[ 161 ][ 321 ],
   alphaCSR[ 161 ][ 322 ],
   alphaCSR[ 161 ][ 323 ],
   alphaCSR[ 161 ][ 324 ],
   alphaCSR[ 161 ][ 325 ],
   alphaCSR[ 161 ][ 326 ],
   alphaCSR[ 161 ][ 327 ],
   alphaCSR[ 161 ][ 328 ],
   alphaCSR[ 161 ][ 329 ],
   alphaCSR[ 161 ][ 330 ],
   alphaCSR[ 161 ][ 331 ],
   alphaCSR[ 161 ][ 332 ],
   alphaCSR[ 161 ][ 333 ],
   alphaCSR[ 161 ][ 334 ],
   alphaCSR[ 161 ][ 335 ],
   alphaCSR[ 161 ][ 336 ],
   alphaCSR[ 161 ][ 337 ],
   alphaCSR[ 161 ][ 338 ],
   alphaCSR[ 161 ][ 339 ],
   alphaCSR[ 161 ][ 340 ],
   alphaCSR[ 161 ][ 341 ],
   alphaCSR[ 161 ][ 342 ],
   alphaCSR[ 161 ][ 343 ],
   alphaCSR[ 161 ][ 344 ],
   alphaCSR[ 161 ][ 345 ],
   alphaCSR[ 161 ][ 346 ],
   alphaCSR[ 161 ][ 347 ],
   alphaCSR[ 161 ][ 348 ],
   alphaCSR[ 161 ][ 349 ],
   alphaCSR[ 161 ][ 350 ],
   alphaCSR[ 161 ][ 351 ],
   alphaCSR[ 161 ][ 352 ],
   alphaCSR[ 161 ][ 353 ],
   alphaCSR[ 161 ][ 354 ],
   alphaCSR[ 161 ][ 355 ],
   alphaCSR[ 161 ][ 356 ],
   alphaCSR[ 161 ][ 357 ],
   alphaCSR[ 161 ][ 358 ],
   alphaCSR[ 161 ][ 359 ],
   alphaCSR[ 161 ][ 360 ],
   alphaCSR[ 161 ][ 361 ],
   alphaCSR[ 161 ][ 362 ],
   alphaCSR[ 161 ][ 363 ],
   alphaCSR[ 161 ][ 364 ],
   alphaCSR[ 161 ][ 365 ],
   alphaCSR[ 161 ][ 366 ],
   alphaCSR[ 161 ][ 367 ],
   alphaCSR[ 161 ][ 368 ],
   alphaCSR[ 161 ][ 369 ],
   alphaCSR[ 161 ][ 370 ],
   alphaCSR[ 161 ][ 371 ],
   alphaCSR[ 161 ][ 372 ],
   alphaCSR[ 161 ][ 373 ],
   alphaCSR[ 161 ][ 374 ],
   alphaCSR[ 161 ][ 375 ],
   alphaCSR[ 161 ][ 376 ],
   alphaCSR[ 161 ][ 377 ],
   alphaCSR[ 161 ][ 378 ],
   alphaCSR[ 161 ][ 379 ],
   alphaCSR[ 161 ][ 380 ],
   alphaCSR[ 161 ][ 381 ],
   alphaCSR[ 161 ][ 382 ],
   alphaCSR[ 161 ][ 383 ],
   alphaCSR[ 162 ][ 0 ],
   alphaCSR[ 162 ][ 1 ],
   alphaCSR[ 162 ][ 2 ],
   alphaCSR[ 162 ][ 3 ],
   alphaCSR[ 162 ][ 4 ],
   alphaCSR[ 162 ][ 5 ],
   alphaCSR[ 162 ][ 6 ],
   alphaCSR[ 162 ][ 7 ],
   alphaCSR[ 162 ][ 8 ],
   alphaCSR[ 162 ][ 9 ],
   alphaCSR[ 162 ][ 10 ],
   alphaCSR[ 162 ][ 11 ],
   alphaCSR[ 162 ][ 12 ],
   alphaCSR[ 162 ][ 13 ],
   alphaCSR[ 162 ][ 14 ],
   alphaCSR[ 162 ][ 15 ],
   alphaCSR[ 162 ][ 16 ],
   alphaCSR[ 162 ][ 17 ],
   alphaCSR[ 162 ][ 18 ],
   alphaCSR[ 162 ][ 19 ],
   alphaCSR[ 162 ][ 20 ],
   alphaCSR[ 162 ][ 21 ],
   alphaCSR[ 162 ][ 22 ],
   alphaCSR[ 162 ][ 23 ],
   alphaCSR[ 162 ][ 24 ],
   alphaCSR[ 162 ][ 25 ],
   alphaCSR[ 162 ][ 26 ],
   alphaCSR[ 162 ][ 27 ],
   alphaCSR[ 162 ][ 28 ],
   alphaCSR[ 162 ][ 29 ],
   alphaCSR[ 162 ][ 30 ],
   alphaCSR[ 162 ][ 31 ],
   alphaCSR[ 162 ][ 32 ],
   alphaCSR[ 162 ][ 33 ],
   alphaCSR[ 162 ][ 34 ],
   alphaCSR[ 162 ][ 35 ],
   alphaCSR[ 162 ][ 36 ],
   alphaCSR[ 162 ][ 37 ],
   alphaCSR[ 162 ][ 38 ],
   alphaCSR[ 162 ][ 39 ],
   alphaCSR[ 162 ][ 40 ],
   alphaCSR[ 162 ][ 41 ],
   alphaCSR[ 162 ][ 42 ],
   alphaCSR[ 162 ][ 43 ],
   alphaCSR[ 162 ][ 44 ],
   alphaCSR[ 162 ][ 45 ],
   alphaCSR[ 162 ][ 46 ],
   alphaCSR[ 162 ][ 47 ],
   alphaCSR[ 162 ][ 48 ],
   alphaCSR[ 162 ][ 49 ],
   alphaCSR[ 162 ][ 50 ],
   alphaCSR[ 162 ][ 51 ],
   alphaCSR[ 162 ][ 52 ],
   alphaCSR[ 162 ][ 53 ],
   alphaCSR[ 162 ][ 54 ],
   alphaCSR[ 162 ][ 55 ],
   alphaCSR[ 162 ][ 56 ],
   alphaCSR[ 162 ][ 57 ],
   alphaCSR[ 162 ][ 58 ],
   alphaCSR[ 162 ][ 59 ],
   alphaCSR[ 162 ][ 60 ],
   alphaCSR[ 162 ][ 61 ],
   alphaCSR[ 162 ][ 62 ],
   alphaCSR[ 162 ][ 63 ],
   alphaCSR[ 162 ][ 64 ],
   alphaCSR[ 162 ][ 65 ],
   alphaCSR[ 162 ][ 66 ],
   alphaCSR[ 162 ][ 67 ],
   alphaCSR[ 162 ][ 68 ],
   alphaCSR[ 162 ][ 69 ],
   alphaCSR[ 162 ][ 70 ],
   alphaCSR[ 162 ][ 71 ],
   alphaCSR[ 162 ][ 72 ],
   alphaCSR[ 162 ][ 73 ],
   alphaCSR[ 162 ][ 74 ],
   alphaCSR[ 162 ][ 75 ],
   alphaCSR[ 162 ][ 76 ],
   alphaCSR[ 162 ][ 77 ],
   alphaCSR[ 162 ][ 78 ],
   alphaCSR[ 162 ][ 79 ],
   alphaCSR[ 162 ][ 80 ],
   alphaCSR[ 162 ][ 81 ],
   alphaCSR[ 162 ][ 82 ],
   alphaCSR[ 162 ][ 83 ],
   alphaCSR[ 162 ][ 84 ],
   alphaCSR[ 162 ][ 85 ],
   alphaCSR[ 162 ][ 86 ],
   alphaCSR[ 162 ][ 87 ],
   alphaCSR[ 162 ][ 88 ],
   alphaCSR[ 162 ][ 89 ],
   alphaCSR[ 162 ][ 90 ],
   alphaCSR[ 162 ][ 91 ],
   alphaCSR[ 162 ][ 92 ],
   alphaCSR[ 162 ][ 93 ],
   alphaCSR[ 162 ][ 94 ],
   alphaCSR[ 162 ][ 95 ],
   alphaCSR[ 162 ][ 96 ],
   alphaCSR[ 162 ][ 97 ],
   alphaCSR[ 162 ][ 98 ],
   alphaCSR[ 162 ][ 99 ],
   alphaCSR[ 162 ][ 100 ],
   alphaCSR[ 162 ][ 101 ],
   alphaCSR[ 162 ][ 102 ],
   alphaCSR[ 162 ][ 103 ],
   alphaCSR[ 162 ][ 104 ],
   alphaCSR[ 162 ][ 105 ],
   alphaCSR[ 162 ][ 106 ],
   alphaCSR[ 162 ][ 107 ],
   alphaCSR[ 162 ][ 108 ],
   alphaCSR[ 162 ][ 109 ],
   alphaCSR[ 162 ][ 110 ],
   alphaCSR[ 162 ][ 111 ],
   alphaCSR[ 162 ][ 112 ],
   alphaCSR[ 162 ][ 113 ],
   alphaCSR[ 162 ][ 114 ],
   alphaCSR[ 162 ][ 115 ],
   alphaCSR[ 162 ][ 116 ],
   alphaCSR[ 162 ][ 117 ],
   alphaCSR[ 162 ][ 118 ],
   alphaCSR[ 162 ][ 119 ],
   alphaCSR[ 162 ][ 120 ],
   alphaCSR[ 162 ][ 121 ],
   alphaCSR[ 162 ][ 122 ],
   alphaCSR[ 162 ][ 123 ],
   alphaCSR[ 162 ][ 124 ],
   alphaCSR[ 162 ][ 125 ],
   alphaCSR[ 162 ][ 126 ],
   alphaCSR[ 162 ][ 127 ],
   alphaCSR[ 162 ][ 128 ],
   alphaCSR[ 162 ][ 129 ],
   alphaCSR[ 162 ][ 130 ],
   alphaCSR[ 162 ][ 131 ],
   alphaCSR[ 162 ][ 132 ],
   alphaCSR[ 162 ][ 133 ],
   alphaCSR[ 162 ][ 134 ],
   alphaCSR[ 162 ][ 135 ],
   alphaCSR[ 162 ][ 136 ],
   alphaCSR[ 162 ][ 137 ],
   alphaCSR[ 162 ][ 138 ],
   alphaCSR[ 162 ][ 139 ],
   alphaCSR[ 162 ][ 140 ],
   alphaCSR[ 162 ][ 141 ],
   alphaCSR[ 162 ][ 142 ],
   alphaCSR[ 162 ][ 143 ],
   alphaCSR[ 162 ][ 144 ],
   alphaCSR[ 162 ][ 145 ],
   alphaCSR[ 162 ][ 146 ],
   alphaCSR[ 162 ][ 147 ],
   alphaCSR[ 162 ][ 148 ],
   alphaCSR[ 162 ][ 149 ],
   alphaCSR[ 162 ][ 150 ],
   alphaCSR[ 162 ][ 151 ],
   alphaCSR[ 162 ][ 152 ],
   alphaCSR[ 162 ][ 153 ],
   alphaCSR[ 162 ][ 154 ],
   alphaCSR[ 162 ][ 155 ],
   alphaCSR[ 162 ][ 156 ],
   alphaCSR[ 162 ][ 157 ],
   alphaCSR[ 162 ][ 158 ],
   alphaCSR[ 162 ][ 159 ],
   alphaCSR[ 162 ][ 160 ],
   alphaCSR[ 162 ][ 161 ],
   alphaCSR[ 162 ][ 162 ],
   alphaCSR[ 162 ][ 163 ],
   alphaCSR[ 162 ][ 164 ],
   alphaCSR[ 162 ][ 165 ],
   alphaCSR[ 162 ][ 166 ],
   alphaCSR[ 162 ][ 167 ],
   alphaCSR[ 162 ][ 168 ],
   alphaCSR[ 162 ][ 169 ],
   alphaCSR[ 162 ][ 170 ],
   alphaCSR[ 162 ][ 171 ],
   alphaCSR[ 162 ][ 172 ],
   alphaCSR[ 162 ][ 173 ],
   alphaCSR[ 162 ][ 174 ],
   alphaCSR[ 162 ][ 175 ],
   alphaCSR[ 162 ][ 176 ],
   alphaCSR[ 162 ][ 177 ],
   alphaCSR[ 162 ][ 178 ],
   alphaCSR[ 162 ][ 179 ],
   alphaCSR[ 162 ][ 180 ],
   alphaCSR[ 162 ][ 181 ],
   alphaCSR[ 162 ][ 182 ],
   alphaCSR[ 162 ][ 183 ],
   alphaCSR[ 162 ][ 184 ],
   alphaCSR[ 162 ][ 185 ],
   alphaCSR[ 162 ][ 186 ],
   alphaCSR[ 162 ][ 187 ],
   alphaCSR[ 162 ][ 188 ],
   alphaCSR[ 162 ][ 189 ],
   alphaCSR[ 162 ][ 190 ],
   alphaCSR[ 162 ][ 191 ],
   alphaCSR[ 162 ][ 192 ],
   alphaCSR[ 162 ][ 193 ],
   alphaCSR[ 162 ][ 194 ],
   alphaCSR[ 162 ][ 195 ],
   alphaCSR[ 162 ][ 196 ],
   alphaCSR[ 162 ][ 197 ],
   alphaCSR[ 162 ][ 198 ],
   alphaCSR[ 162 ][ 199 ],
   alphaCSR[ 162 ][ 200 ],
   alphaCSR[ 162 ][ 201 ],
   alphaCSR[ 162 ][ 202 ],
   alphaCSR[ 162 ][ 203 ],
   alphaCSR[ 162 ][ 204 ],
   alphaCSR[ 162 ][ 205 ],
   alphaCSR[ 162 ][ 206 ],
   alphaCSR[ 162 ][ 207 ],
   alphaCSR[ 162 ][ 208 ],
   alphaCSR[ 162 ][ 209 ],
   alphaCSR[ 162 ][ 210 ],
   alphaCSR[ 162 ][ 211 ],
   alphaCSR[ 162 ][ 212 ],
   alphaCSR[ 162 ][ 213 ],
   alphaCSR[ 162 ][ 214 ],
   alphaCSR[ 162 ][ 215 ],
   alphaCSR[ 162 ][ 216 ],
   alphaCSR[ 162 ][ 217 ],
   alphaCSR[ 162 ][ 218 ],
   alphaCSR[ 162 ][ 219 ],
   alphaCSR[ 162 ][ 220 ],
   alphaCSR[ 162 ][ 221 ],
   alphaCSR[ 162 ][ 222 ],
   alphaCSR[ 162 ][ 223 ],
   alphaCSR[ 162 ][ 224 ],
   alphaCSR[ 162 ][ 225 ],
   alphaCSR[ 162 ][ 226 ],
   alphaCSR[ 162 ][ 227 ],
   alphaCSR[ 162 ][ 228 ],
   alphaCSR[ 162 ][ 229 ],
   alphaCSR[ 162 ][ 230 ],
   alphaCSR[ 162 ][ 231 ],
   alphaCSR[ 162 ][ 232 ],
   alphaCSR[ 162 ][ 233 ],
   alphaCSR[ 162 ][ 234 ],
   alphaCSR[ 162 ][ 235 ],
   alphaCSR[ 162 ][ 236 ],
   alphaCSR[ 162 ][ 237 ],
   alphaCSR[ 162 ][ 238 ],
   alphaCSR[ 162 ][ 239 ],
   alphaCSR[ 162 ][ 240 ],
   alphaCSR[ 162 ][ 241 ],
   alphaCSR[ 162 ][ 242 ],
   alphaCSR[ 162 ][ 243 ],
   alphaCSR[ 162 ][ 244 ],
   alphaCSR[ 162 ][ 245 ],
   alphaCSR[ 162 ][ 246 ],
   alphaCSR[ 162 ][ 247 ],
   alphaCSR[ 162 ][ 248 ],
   alphaCSR[ 162 ][ 249 ],
   alphaCSR[ 162 ][ 250 ],
   alphaCSR[ 162 ][ 251 ],
   alphaCSR[ 162 ][ 252 ],
   alphaCSR[ 162 ][ 253 ],
   alphaCSR[ 162 ][ 254 ],
   alphaCSR[ 162 ][ 255 ],
   alphaCSR[ 162 ][ 256 ],
   alphaCSR[ 162 ][ 257 ],
   alphaCSR[ 162 ][ 258 ],
   alphaCSR[ 162 ][ 259 ],
   alphaCSR[ 162 ][ 260 ],
   alphaCSR[ 162 ][ 261 ],
   alphaCSR[ 162 ][ 262 ],
   alphaCSR[ 162 ][ 263 ],
   alphaCSR[ 162 ][ 264 ],
   alphaCSR[ 162 ][ 265 ],
   alphaCSR[ 162 ][ 266 ],
   alphaCSR[ 162 ][ 267 ],
   alphaCSR[ 162 ][ 268 ],
   alphaCSR[ 162 ][ 269 ],
   alphaCSR[ 162 ][ 270 ],
   alphaCSR[ 162 ][ 271 ],
   alphaCSR[ 162 ][ 272 ],
   alphaCSR[ 162 ][ 273 ],
   alphaCSR[ 162 ][ 274 ],
   alphaCSR[ 162 ][ 275 ],
   alphaCSR[ 162 ][ 276 ],
   alphaCSR[ 162 ][ 277 ],
   alphaCSR[ 162 ][ 278 ],
   alphaCSR[ 162 ][ 279 ],
   alphaCSR[ 162 ][ 280 ],
   alphaCSR[ 162 ][ 281 ],
   alphaCSR[ 162 ][ 282 ],
   alphaCSR[ 162 ][ 283 ],
   alphaCSR[ 162 ][ 284 ],
   alphaCSR[ 162 ][ 285 ],
   alphaCSR[ 162 ][ 286 ],
   alphaCSR[ 162 ][ 287 ],
   alphaCSR[ 162 ][ 288 ],
   alphaCSR[ 162 ][ 289 ],
   alphaCSR[ 162 ][ 290 ],
   alphaCSR[ 162 ][ 291 ],
   alphaCSR[ 162 ][ 292 ],
   alphaCSR[ 162 ][ 293 ],
   alphaCSR[ 162 ][ 294 ],
   alphaCSR[ 162 ][ 295 ],
   alphaCSR[ 162 ][ 296 ],
   alphaCSR[ 162 ][ 297 ],
   alphaCSR[ 162 ][ 298 ],
   alphaCSR[ 162 ][ 299 ],
   alphaCSR[ 162 ][ 300 ],
   alphaCSR[ 162 ][ 301 ],
   alphaCSR[ 162 ][ 302 ],
   alphaCSR[ 162 ][ 303 ],
   alphaCSR[ 162 ][ 304 ],
   alphaCSR[ 162 ][ 305 ],
   alphaCSR[ 162 ][ 306 ],
   alphaCSR[ 162 ][ 307 ],
   alphaCSR[ 162 ][ 308 ],
   alphaCSR[ 162 ][ 309 ],
   alphaCSR[ 162 ][ 310 ],
   alphaCSR[ 162 ][ 311 ],
   alphaCSR[ 162 ][ 312 ],
   alphaCSR[ 162 ][ 313 ],
   alphaCSR[ 162 ][ 314 ],
   alphaCSR[ 162 ][ 315 ],
   alphaCSR[ 162 ][ 316 ],
   alphaCSR[ 162 ][ 317 ],
   alphaCSR[ 162 ][ 318 ],
   alphaCSR[ 162 ][ 319 ],
   alphaCSR[ 162 ][ 320 ],
   alphaCSR[ 162 ][ 321 ],
   alphaCSR[ 162 ][ 322 ],
   alphaCSR[ 162 ][ 323 ],
   alphaCSR[ 162 ][ 324 ],
   alphaCSR[ 162 ][ 325 ],
   alphaCSR[ 162 ][ 326 ],
   alphaCSR[ 162 ][ 327 ],
   alphaCSR[ 162 ][ 328 ],
   alphaCSR[ 162 ][ 329 ],
   alphaCSR[ 162 ][ 330 ],
   alphaCSR[ 162 ][ 331 ],
   alphaCSR[ 162 ][ 332 ],
   alphaCSR[ 162 ][ 333 ],
   alphaCSR[ 162 ][ 334 ],
   alphaCSR[ 162 ][ 335 ],
   alphaCSR[ 162 ][ 336 ],
   alphaCSR[ 162 ][ 337 ],
   alphaCSR[ 162 ][ 338 ],
   alphaCSR[ 162 ][ 339 ],
   alphaCSR[ 162 ][ 340 ],
   alphaCSR[ 162 ][ 341 ],
   alphaCSR[ 162 ][ 342 ],
   alphaCSR[ 162 ][ 343 ],
   alphaCSR[ 162 ][ 344 ],
   alphaCSR[ 162 ][ 345 ],
   alphaCSR[ 162 ][ 346 ],
   alphaCSR[ 162 ][ 347 ],
   alphaCSR[ 162 ][ 348 ],
   alphaCSR[ 162 ][ 349 ],
   alphaCSR[ 162 ][ 350 ],
   alphaCSR[ 162 ][ 351 ],
   alphaCSR[ 162 ][ 352 ],
   alphaCSR[ 162 ][ 353 ],
   alphaCSR[ 162 ][ 354 ],
   alphaCSR[ 162 ][ 355 ],
   alphaCSR[ 162 ][ 356 ],
   alphaCSR[ 162 ][ 357 ],
   alphaCSR[ 162 ][ 358 ],
   alphaCSR[ 162 ][ 359 ],
   alphaCSR[ 162 ][ 360 ],
   alphaCSR[ 162 ][ 361 ],
   alphaCSR[ 162 ][ 362 ],
   alphaCSR[ 162 ][ 363 ],
   alphaCSR[ 162 ][ 364 ],
   alphaCSR[ 162 ][ 365 ],
   alphaCSR[ 162 ][ 366 ],
   alphaCSR[ 162 ][ 367 ],
   alphaCSR[ 162 ][ 368 ],
   alphaCSR[ 162 ][ 369 ],
   alphaCSR[ 162 ][ 370 ],
   alphaCSR[ 162 ][ 371 ],
   alphaCSR[ 162 ][ 372 ],
   alphaCSR[ 162 ][ 373 ],
   alphaCSR[ 162 ][ 374 ],
   alphaCSR[ 162 ][ 375 ],
   alphaCSR[ 162 ][ 376 ],
   alphaCSR[ 162 ][ 377 ],
   alphaCSR[ 162 ][ 378 ],
   alphaCSR[ 162 ][ 379 ],
   alphaCSR[ 162 ][ 380 ],
   alphaCSR[ 162 ][ 381 ],
   alphaCSR[ 162 ][ 382 ],
   alphaCSR[ 162 ][ 383 ],
   alphaCSR[ 163 ][ 0 ],
   alphaCSR[ 163 ][ 1 ],
   alphaCSR[ 163 ][ 2 ],
   alphaCSR[ 163 ][ 3 ],
   alphaCSR[ 163 ][ 4 ],
   alphaCSR[ 163 ][ 5 ],
   alphaCSR[ 163 ][ 6 ],
   alphaCSR[ 163 ][ 7 ],
   alphaCSR[ 163 ][ 8 ],
   alphaCSR[ 163 ][ 9 ],
   alphaCSR[ 163 ][ 10 ],
   alphaCSR[ 163 ][ 11 ],
   alphaCSR[ 163 ][ 12 ],
   alphaCSR[ 163 ][ 13 ],
   alphaCSR[ 163 ][ 14 ],
   alphaCSR[ 163 ][ 15 ],
   alphaCSR[ 163 ][ 16 ],
   alphaCSR[ 163 ][ 17 ],
   alphaCSR[ 163 ][ 18 ],
   alphaCSR[ 163 ][ 19 ],
   alphaCSR[ 163 ][ 20 ],
   alphaCSR[ 163 ][ 21 ],
   alphaCSR[ 163 ][ 22 ],
   alphaCSR[ 163 ][ 23 ],
   alphaCSR[ 163 ][ 24 ],
   alphaCSR[ 163 ][ 25 ],
   alphaCSR[ 163 ][ 26 ],
   alphaCSR[ 163 ][ 27 ],
   alphaCSR[ 163 ][ 28 ],
   alphaCSR[ 163 ][ 29 ],
   alphaCSR[ 163 ][ 30 ],
   alphaCSR[ 163 ][ 31 ],
   alphaCSR[ 163 ][ 32 ],
   alphaCSR[ 163 ][ 33 ],
   alphaCSR[ 163 ][ 34 ],
   alphaCSR[ 163 ][ 35 ],
   alphaCSR[ 163 ][ 36 ],
   alphaCSR[ 163 ][ 37 ],
   alphaCSR[ 163 ][ 38 ],
   alphaCSR[ 163 ][ 39 ],
   alphaCSR[ 163 ][ 40 ],
   alphaCSR[ 163 ][ 41 ],
   alphaCSR[ 163 ][ 42 ],
   alphaCSR[ 163 ][ 43 ],
   alphaCSR[ 163 ][ 44 ],
   alphaCSR[ 163 ][ 45 ],
   alphaCSR[ 163 ][ 46 ],
   alphaCSR[ 163 ][ 47 ],
   alphaCSR[ 163 ][ 48 ],
   alphaCSR[ 163 ][ 49 ],
   alphaCSR[ 163 ][ 50 ],
   alphaCSR[ 163 ][ 51 ],
   alphaCSR[ 163 ][ 52 ],
   alphaCSR[ 163 ][ 53 ],
   alphaCSR[ 163 ][ 54 ],
   alphaCSR[ 163 ][ 55 ],
   alphaCSR[ 163 ][ 56 ],
   alphaCSR[ 163 ][ 57 ],
   alphaCSR[ 163 ][ 58 ],
   alphaCSR[ 163 ][ 59 ],
   alphaCSR[ 163 ][ 60 ],
   alphaCSR[ 163 ][ 61 ],
   alphaCSR[ 163 ][ 62 ],
   alphaCSR[ 163 ][ 63 ],
   alphaCSR[ 163 ][ 64 ],
   alphaCSR[ 163 ][ 65 ],
   alphaCSR[ 163 ][ 66 ],
   alphaCSR[ 163 ][ 67 ],
   alphaCSR[ 163 ][ 68 ],
   alphaCSR[ 163 ][ 69 ],
   alphaCSR[ 163 ][ 70 ],
   alphaCSR[ 163 ][ 71 ],
   alphaCSR[ 163 ][ 72 ],
   alphaCSR[ 163 ][ 73 ],
   alphaCSR[ 163 ][ 74 ],
   alphaCSR[ 163 ][ 75 ],
   alphaCSR[ 163 ][ 76 ],
   alphaCSR[ 163 ][ 77 ],
   alphaCSR[ 163 ][ 78 ],
   alphaCSR[ 163 ][ 79 ],
   alphaCSR[ 163 ][ 80 ],
   alphaCSR[ 163 ][ 81 ],
   alphaCSR[ 163 ][ 82 ],
   alphaCSR[ 163 ][ 83 ],
   alphaCSR[ 163 ][ 84 ],
   alphaCSR[ 163 ][ 85 ],
   alphaCSR[ 163 ][ 86 ],
   alphaCSR[ 163 ][ 87 ],
   alphaCSR[ 163 ][ 88 ],
   alphaCSR[ 163 ][ 89 ],
   alphaCSR[ 163 ][ 90 ],
   alphaCSR[ 163 ][ 91 ],
   alphaCSR[ 163 ][ 92 ],
   alphaCSR[ 163 ][ 93 ],
   alphaCSR[ 163 ][ 94 ],
   alphaCSR[ 163 ][ 95 ],
   alphaCSR[ 163 ][ 96 ],
   alphaCSR[ 163 ][ 97 ],
   alphaCSR[ 163 ][ 98 ],
   alphaCSR[ 163 ][ 99 ],
   alphaCSR[ 163 ][ 100 ],
   alphaCSR[ 163 ][ 101 ],
   alphaCSR[ 163 ][ 102 ],
   alphaCSR[ 163 ][ 103 ],
   alphaCSR[ 163 ][ 104 ],
   alphaCSR[ 163 ][ 105 ],
   alphaCSR[ 163 ][ 106 ],
   alphaCSR[ 163 ][ 107 ],
   alphaCSR[ 163 ][ 108 ],
   alphaCSR[ 163 ][ 109 ],
   alphaCSR[ 163 ][ 110 ],
   alphaCSR[ 163 ][ 111 ],
   alphaCSR[ 163 ][ 112 ],
   alphaCSR[ 163 ][ 113 ],
   alphaCSR[ 163 ][ 114 ],
   alphaCSR[ 163 ][ 115 ],
   alphaCSR[ 163 ][ 116 ],
   alphaCSR[ 163 ][ 117 ],
   alphaCSR[ 163 ][ 118 ],
   alphaCSR[ 163 ][ 119 ],
   alphaCSR[ 163 ][ 120 ],
   alphaCSR[ 163 ][ 121 ],
   alphaCSR[ 163 ][ 122 ],
   alphaCSR[ 163 ][ 123 ],
   alphaCSR[ 163 ][ 124 ],
   alphaCSR[ 163 ][ 125 ],
   alphaCSR[ 163 ][ 126 ],
   alphaCSR[ 163 ][ 127 ],
   alphaCSR[ 163 ][ 128 ],
   alphaCSR[ 163 ][ 129 ],
   alphaCSR[ 163 ][ 130 ],
   alphaCSR[ 163 ][ 131 ],
   alphaCSR[ 163 ][ 132 ],
   alphaCSR[ 163 ][ 133 ],
   alphaCSR[ 163 ][ 134 ],
   alphaCSR[ 163 ][ 135 ],
   alphaCSR[ 163 ][ 136 ],
   alphaCSR[ 163 ][ 137 ],
   alphaCSR[ 163 ][ 138 ],
   alphaCSR[ 163 ][ 139 ],
   alphaCSR[ 163 ][ 140 ],
   alphaCSR[ 163 ][ 141 ],
   alphaCSR[ 163 ][ 142 ],
   alphaCSR[ 163 ][ 143 ],
   alphaCSR[ 163 ][ 144 ],
   alphaCSR[ 163 ][ 145 ],
   alphaCSR[ 163 ][ 146 ],
   alphaCSR[ 163 ][ 147 ],
   alphaCSR[ 163 ][ 148 ],
   alphaCSR[ 163 ][ 149 ],
   alphaCSR[ 163 ][ 150 ],
   alphaCSR[ 163 ][ 151 ],
   alphaCSR[ 163 ][ 152 ],
   alphaCSR[ 163 ][ 153 ],
   alphaCSR[ 163 ][ 154 ],
   alphaCSR[ 163 ][ 155 ],
   alphaCSR[ 163 ][ 156 ],
   alphaCSR[ 163 ][ 157 ],
   alphaCSR[ 163 ][ 158 ],
   alphaCSR[ 163 ][ 159 ],
   alphaCSR[ 163 ][ 160 ],
   alphaCSR[ 163 ][ 161 ],
   alphaCSR[ 163 ][ 162 ],
   alphaCSR[ 163 ][ 163 ],
   alphaCSR[ 163 ][ 164 ],
   alphaCSR[ 163 ][ 165 ],
   alphaCSR[ 163 ][ 166 ],
   alphaCSR[ 163 ][ 167 ],
   alphaCSR[ 163 ][ 168 ],
   alphaCSR[ 163 ][ 169 ],
   alphaCSR[ 163 ][ 170 ],
   alphaCSR[ 163 ][ 171 ],
   alphaCSR[ 163 ][ 172 ],
   alphaCSR[ 163 ][ 173 ],
   alphaCSR[ 163 ][ 174 ],
   alphaCSR[ 163 ][ 175 ],
   alphaCSR[ 163 ][ 176 ],
   alphaCSR[ 163 ][ 177 ],
   alphaCSR[ 163 ][ 178 ],
   alphaCSR[ 163 ][ 179 ],
   alphaCSR[ 163 ][ 180 ],
   alphaCSR[ 163 ][ 181 ],
   alphaCSR[ 163 ][ 182 ],
   alphaCSR[ 163 ][ 183 ],
   alphaCSR[ 163 ][ 184 ],
   alphaCSR[ 163 ][ 185 ],
   alphaCSR[ 163 ][ 186 ],
   alphaCSR[ 163 ][ 187 ],
   alphaCSR[ 163 ][ 188 ],
   alphaCSR[ 163 ][ 189 ],
   alphaCSR[ 163 ][ 190 ],
   alphaCSR[ 163 ][ 191 ],
   alphaCSR[ 163 ][ 192 ],
   alphaCSR[ 163 ][ 193 ],
   alphaCSR[ 163 ][ 194 ],
   alphaCSR[ 163 ][ 195 ],
   alphaCSR[ 163 ][ 196 ],
   alphaCSR[ 163 ][ 197 ],
   alphaCSR[ 163 ][ 198 ],
   alphaCSR[ 163 ][ 199 ],
   alphaCSR[ 163 ][ 200 ],
   alphaCSR[ 163 ][ 201 ],
   alphaCSR[ 163 ][ 202 ],
   alphaCSR[ 163 ][ 203 ],
   alphaCSR[ 163 ][ 204 ],
   alphaCSR[ 163 ][ 205 ],
   alphaCSR[ 163 ][ 206 ],
   alphaCSR[ 163 ][ 207 ],
   alphaCSR[ 163 ][ 208 ],
   alphaCSR[ 163 ][ 209 ],
   alphaCSR[ 163 ][ 210 ],
   alphaCSR[ 163 ][ 211 ],
   alphaCSR[ 163 ][ 212 ],
   alphaCSR[ 163 ][ 213 ],
   alphaCSR[ 163 ][ 214 ],
   alphaCSR[ 163 ][ 215 ],
   alphaCSR[ 163 ][ 216 ],
   alphaCSR[ 163 ][ 217 ],
   alphaCSR[ 163 ][ 218 ],
   alphaCSR[ 163 ][ 219 ],
   alphaCSR[ 163 ][ 220 ],
   alphaCSR[ 163 ][ 221 ],
   alphaCSR[ 163 ][ 222 ],
   alphaCSR[ 163 ][ 223 ],
   alphaCSR[ 163 ][ 224 ],
   alphaCSR[ 163 ][ 225 ],
   alphaCSR[ 163 ][ 226 ],
   alphaCSR[ 163 ][ 227 ],
   alphaCSR[ 163 ][ 228 ],
   alphaCSR[ 163 ][ 229 ],
   alphaCSR[ 163 ][ 230 ],
   alphaCSR[ 163 ][ 231 ],
   alphaCSR[ 163 ][ 232 ],
   alphaCSR[ 163 ][ 233 ],
   alphaCSR[ 163 ][ 234 ],
   alphaCSR[ 163 ][ 235 ],
   alphaCSR[ 163 ][ 236 ],
   alphaCSR[ 163 ][ 237 ],
   alphaCSR[ 163 ][ 238 ],
   alphaCSR[ 163 ][ 239 ],
   alphaCSR[ 163 ][ 240 ],
   alphaCSR[ 163 ][ 241 ],
   alphaCSR[ 163 ][ 242 ],
   alphaCSR[ 163 ][ 243 ],
   alphaCSR[ 163 ][ 244 ],
   alphaCSR[ 163 ][ 245 ],
   alphaCSR[ 163 ][ 246 ],
   alphaCSR[ 163 ][ 247 ],
   alphaCSR[ 163 ][ 248 ],
   alphaCSR[ 163 ][ 249 ],
   alphaCSR[ 163 ][ 250 ],
   alphaCSR[ 163 ][ 251 ],
   alphaCSR[ 163 ][ 252 ],
   alphaCSR[ 163 ][ 253 ],
   alphaCSR[ 163 ][ 254 ],
   alphaCSR[ 163 ][ 255 ],
   alphaCSR[ 163 ][ 256 ],
   alphaCSR[ 163 ][ 257 ],
   alphaCSR[ 163 ][ 258 ],
   alphaCSR[ 163 ][ 259 ],
   alphaCSR[ 163 ][ 260 ],
   alphaCSR[ 163 ][ 261 ],
   alphaCSR[ 163 ][ 262 ],
   alphaCSR[ 163 ][ 263 ],
   alphaCSR[ 163 ][ 264 ],
   alphaCSR[ 163 ][ 265 ],
   alphaCSR[ 163 ][ 266 ],
   alphaCSR[ 163 ][ 267 ],
   alphaCSR[ 163 ][ 268 ],
   alphaCSR[ 163 ][ 269 ],
   alphaCSR[ 163 ][ 270 ],
   alphaCSR[ 163 ][ 271 ],
   alphaCSR[ 163 ][ 272 ],
   alphaCSR[ 163 ][ 273 ],
   alphaCSR[ 163 ][ 274 ],
   alphaCSR[ 163 ][ 275 ],
   alphaCSR[ 163 ][ 276 ],
   alphaCSR[ 163 ][ 277 ],
   alphaCSR[ 163 ][ 278 ],
   alphaCSR[ 163 ][ 279 ],
   alphaCSR[ 163 ][ 280 ],
   alphaCSR[ 163 ][ 281 ],
   alphaCSR[ 163 ][ 282 ],
   alphaCSR[ 163 ][ 283 ],
   alphaCSR[ 163 ][ 284 ],
   alphaCSR[ 163 ][ 285 ],
   alphaCSR[ 163 ][ 286 ],
   alphaCSR[ 163 ][ 287 ],
   alphaCSR[ 163 ][ 288 ],
   alphaCSR[ 163 ][ 289 ],
   alphaCSR[ 163 ][ 290 ],
   alphaCSR[ 163 ][ 291 ],
   alphaCSR[ 163 ][ 292 ],
   alphaCSR[ 163 ][ 293 ],
   alphaCSR[ 163 ][ 294 ],
   alphaCSR[ 163 ][ 295 ],
   alphaCSR[ 163 ][ 296 ],
   alphaCSR[ 163 ][ 297 ],
   alphaCSR[ 163 ][ 298 ],
   alphaCSR[ 163 ][ 299 ],
   alphaCSR[ 163 ][ 300 ],
   alphaCSR[ 163 ][ 301 ],
   alphaCSR[ 163 ][ 302 ],
   alphaCSR[ 163 ][ 303 ],
   alphaCSR[ 163 ][ 304 ],
   alphaCSR[ 163 ][ 305 ],
   alphaCSR[ 163 ][ 306 ],
   alphaCSR[ 163 ][ 307 ],
   alphaCSR[ 163 ][ 308 ],
   alphaCSR[ 163 ][ 309 ],
   alphaCSR[ 163 ][ 310 ],
   alphaCSR[ 163 ][ 311 ],
   alphaCSR[ 163 ][ 312 ],
   alphaCSR[ 163 ][ 313 ],
   alphaCSR[ 163 ][ 314 ],
   alphaCSR[ 163 ][ 315 ],
   alphaCSR[ 163 ][ 316 ],
   alphaCSR[ 163 ][ 317 ],
   alphaCSR[ 163 ][ 318 ],
   alphaCSR[ 163 ][ 319 ],
   alphaCSR[ 163 ][ 320 ],
   alphaCSR[ 163 ][ 321 ],
   alphaCSR[ 163 ][ 322 ],
   alphaCSR[ 163 ][ 323 ],
   alphaCSR[ 163 ][ 324 ],
   alphaCSR[ 163 ][ 325 ],
   alphaCSR[ 163 ][ 326 ],
   alphaCSR[ 163 ][ 327 ],
   alphaCSR[ 163 ][ 328 ],
   alphaCSR[ 163 ][ 329 ],
   alphaCSR[ 163 ][ 330 ],
   alphaCSR[ 163 ][ 331 ],
   alphaCSR[ 163 ][ 332 ],
   alphaCSR[ 163 ][ 333 ],
   alphaCSR[ 163 ][ 334 ],
   alphaCSR[ 163 ][ 335 ],
   alphaCSR[ 163 ][ 336 ],
   alphaCSR[ 163 ][ 337 ],
   alphaCSR[ 163 ][ 338 ],
   alphaCSR[ 163 ][ 339 ],
   alphaCSR[ 163 ][ 340 ],
   alphaCSR[ 163 ][ 341 ],
   alphaCSR[ 163 ][ 342 ],
   alphaCSR[ 163 ][ 343 ],
   alphaCSR[ 163 ][ 344 ],
   alphaCSR[ 163 ][ 345 ],
   alphaCSR[ 163 ][ 346 ],
   alphaCSR[ 163 ][ 347 ],
   alphaCSR[ 163 ][ 348 ],
   alphaCSR[ 163 ][ 349 ],
   alphaCSR[ 163 ][ 350 ],
   alphaCSR[ 163 ][ 351 ],
   alphaCSR[ 163 ][ 352 ],
   alphaCSR[ 163 ][ 353 ],
   alphaCSR[ 163 ][ 354 ],
   alphaCSR[ 163 ][ 355 ],
   alphaCSR[ 163 ][ 356 ],
   alphaCSR[ 163 ][ 357 ],
   alphaCSR[ 163 ][ 358 ],
   alphaCSR[ 163 ][ 359 ],
   alphaCSR[ 163 ][ 360 ],
   alphaCSR[ 163 ][ 361 ],
   alphaCSR[ 163 ][ 362 ],
   alphaCSR[ 163 ][ 363 ],
   alphaCSR[ 163 ][ 364 ],
   alphaCSR[ 163 ][ 365 ],
   alphaCSR[ 163 ][ 366 ],
   alphaCSR[ 163 ][ 367 ],
   alphaCSR[ 163 ][ 368 ],
   alphaCSR[ 163 ][ 369 ],
   alphaCSR[ 163 ][ 370 ],
   alphaCSR[ 163 ][ 371 ],
   alphaCSR[ 163 ][ 372 ],
   alphaCSR[ 163 ][ 373 ],
   alphaCSR[ 163 ][ 374 ],
   alphaCSR[ 163 ][ 375 ],
   alphaCSR[ 163 ][ 376 ],
   alphaCSR[ 163 ][ 377 ],
   alphaCSR[ 163 ][ 378 ],
   alphaCSR[ 163 ][ 379 ],
   alphaCSR[ 163 ][ 380 ],
   alphaCSR[ 163 ][ 381 ],
   alphaCSR[ 163 ][ 382 ],
   alphaCSR[ 163 ][ 383 ],
   alphaCSR[ 164 ][ 0 ],
   alphaCSR[ 164 ][ 1 ],
   alphaCSR[ 164 ][ 2 ],
   alphaCSR[ 164 ][ 3 ],
   alphaCSR[ 164 ][ 4 ],
   alphaCSR[ 164 ][ 5 ],
   alphaCSR[ 164 ][ 6 ],
   alphaCSR[ 164 ][ 7 ],
   alphaCSR[ 164 ][ 8 ],
   alphaCSR[ 164 ][ 9 ],
   alphaCSR[ 164 ][ 10 ],
   alphaCSR[ 164 ][ 11 ],
   alphaCSR[ 164 ][ 12 ],
   alphaCSR[ 164 ][ 13 ],
   alphaCSR[ 164 ][ 14 ],
   alphaCSR[ 164 ][ 15 ],
   alphaCSR[ 164 ][ 16 ],
   alphaCSR[ 164 ][ 17 ],
   alphaCSR[ 164 ][ 18 ],
   alphaCSR[ 164 ][ 19 ],
   alphaCSR[ 164 ][ 20 ],
   alphaCSR[ 164 ][ 21 ],
   alphaCSR[ 164 ][ 22 ],
   alphaCSR[ 164 ][ 23 ],
   alphaCSR[ 164 ][ 24 ],
   alphaCSR[ 164 ][ 25 ],
   alphaCSR[ 164 ][ 26 ],
   alphaCSR[ 164 ][ 27 ],
   alphaCSR[ 164 ][ 28 ],
   alphaCSR[ 164 ][ 29 ],
   alphaCSR[ 164 ][ 30 ],
   alphaCSR[ 164 ][ 31 ],
   alphaCSR[ 164 ][ 32 ],
   alphaCSR[ 164 ][ 33 ],
   alphaCSR[ 164 ][ 34 ],
   alphaCSR[ 164 ][ 35 ],
   alphaCSR[ 164 ][ 36 ],
   alphaCSR[ 164 ][ 37 ],
   alphaCSR[ 164 ][ 38 ],
   alphaCSR[ 164 ][ 39 ],
   alphaCSR[ 164 ][ 40 ],
   alphaCSR[ 164 ][ 41 ],
   alphaCSR[ 164 ][ 42 ],
   alphaCSR[ 164 ][ 43 ],
   alphaCSR[ 164 ][ 44 ],
   alphaCSR[ 164 ][ 45 ],
   alphaCSR[ 164 ][ 46 ],
   alphaCSR[ 164 ][ 47 ],
   alphaCSR[ 164 ][ 48 ],
   alphaCSR[ 164 ][ 49 ],
   alphaCSR[ 164 ][ 50 ],
   alphaCSR[ 164 ][ 51 ],
   alphaCSR[ 164 ][ 52 ],
   alphaCSR[ 164 ][ 53 ],
   alphaCSR[ 164 ][ 54 ],
   alphaCSR[ 164 ][ 55 ],
   alphaCSR[ 164 ][ 56 ],
   alphaCSR[ 164 ][ 57 ],
   alphaCSR[ 164 ][ 58 ],
   alphaCSR[ 164 ][ 59 ],
   alphaCSR[ 164 ][ 60 ],
   alphaCSR[ 164 ][ 61 ],
   alphaCSR[ 164 ][ 62 ],
   alphaCSR[ 164 ][ 63 ],
   alphaCSR[ 164 ][ 64 ],
   alphaCSR[ 164 ][ 65 ],
   alphaCSR[ 164 ][ 66 ],
   alphaCSR[ 164 ][ 67 ],
   alphaCSR[ 164 ][ 68 ],
   alphaCSR[ 164 ][ 69 ],
   alphaCSR[ 164 ][ 70 ],
   alphaCSR[ 164 ][ 71 ],
   alphaCSR[ 164 ][ 72 ],
   alphaCSR[ 164 ][ 73 ],
   alphaCSR[ 164 ][ 74 ],
   alphaCSR[ 164 ][ 75 ],
   alphaCSR[ 164 ][ 76 ],
   alphaCSR[ 164 ][ 77 ],
   alphaCSR[ 164 ][ 78 ],
   alphaCSR[ 164 ][ 79 ],
   alphaCSR[ 164 ][ 80 ],
   alphaCSR[ 164 ][ 81 ],
   alphaCSR[ 164 ][ 82 ],
   alphaCSR[ 164 ][ 83 ],
   alphaCSR[ 164 ][ 84 ],
   alphaCSR[ 164 ][ 85 ],
   alphaCSR[ 164 ][ 86 ],
   alphaCSR[ 164 ][ 87 ],
   alphaCSR[ 164 ][ 88 ],
   alphaCSR[ 164 ][ 89 ],
   alphaCSR[ 164 ][ 90 ],
   alphaCSR[ 164 ][ 91 ],
   alphaCSR[ 164 ][ 92 ],
   alphaCSR[ 164 ][ 93 ],
   alphaCSR[ 164 ][ 94 ],
   alphaCSR[ 164 ][ 95 ],
   alphaCSR[ 164 ][ 96 ],
   alphaCSR[ 164 ][ 97 ],
   alphaCSR[ 164 ][ 98 ],
   alphaCSR[ 164 ][ 99 ],
   alphaCSR[ 164 ][ 100 ],
   alphaCSR[ 164 ][ 101 ],
   alphaCSR[ 164 ][ 102 ],
   alphaCSR[ 164 ][ 103 ],
   alphaCSR[ 164 ][ 104 ],
   alphaCSR[ 164 ][ 105 ],
   alphaCSR[ 164 ][ 106 ],
   alphaCSR[ 164 ][ 107 ],
   alphaCSR[ 164 ][ 108 ],
   alphaCSR[ 164 ][ 109 ],
   alphaCSR[ 164 ][ 110 ],
   alphaCSR[ 164 ][ 111 ],
   alphaCSR[ 164 ][ 112 ],
   alphaCSR[ 164 ][ 113 ],
   alphaCSR[ 164 ][ 114 ],
   alphaCSR[ 164 ][ 115 ],
   alphaCSR[ 164 ][ 116 ],
   alphaCSR[ 164 ][ 117 ],
   alphaCSR[ 164 ][ 118 ],
   alphaCSR[ 164 ][ 119 ],
   alphaCSR[ 164 ][ 120 ],
   alphaCSR[ 164 ][ 121 ],
   alphaCSR[ 164 ][ 122 ],
   alphaCSR[ 164 ][ 123 ],
   alphaCSR[ 164 ][ 124 ],
   alphaCSR[ 164 ][ 125 ],
   alphaCSR[ 164 ][ 126 ],
   alphaCSR[ 164 ][ 127 ],
   alphaCSR[ 164 ][ 128 ],
   alphaCSR[ 164 ][ 129 ],
   alphaCSR[ 164 ][ 130 ],
   alphaCSR[ 164 ][ 131 ],
   alphaCSR[ 164 ][ 132 ],
   alphaCSR[ 164 ][ 133 ],
   alphaCSR[ 164 ][ 134 ],
   alphaCSR[ 164 ][ 135 ],
   alphaCSR[ 164 ][ 136 ],
   alphaCSR[ 164 ][ 137 ],
   alphaCSR[ 164 ][ 138 ],
   alphaCSR[ 164 ][ 139 ],
   alphaCSR[ 164 ][ 140 ],
   alphaCSR[ 164 ][ 141 ],
   alphaCSR[ 164 ][ 142 ],
   alphaCSR[ 164 ][ 143 ],
   alphaCSR[ 164 ][ 144 ],
   alphaCSR[ 164 ][ 145 ],
   alphaCSR[ 164 ][ 146 ],
   alphaCSR[ 164 ][ 147 ],
   alphaCSR[ 164 ][ 148 ],
   alphaCSR[ 164 ][ 149 ],
   alphaCSR[ 164 ][ 150 ],
   alphaCSR[ 164 ][ 151 ],
   alphaCSR[ 164 ][ 152 ],
   alphaCSR[ 164 ][ 153 ],
   alphaCSR[ 164 ][ 154 ],
   alphaCSR[ 164 ][ 155 ],
   alphaCSR[ 164 ][ 156 ],
   alphaCSR[ 164 ][ 157 ],
   alphaCSR[ 164 ][ 158 ],
   alphaCSR[ 164 ][ 159 ],
   alphaCSR[ 164 ][ 160 ],
   alphaCSR[ 164 ][ 161 ],
   alphaCSR[ 164 ][ 162 ],
   alphaCSR[ 164 ][ 163 ],
   alphaCSR[ 164 ][ 164 ],
   alphaCSR[ 164 ][ 165 ],
   alphaCSR[ 164 ][ 166 ],
   alphaCSR[ 164 ][ 167 ],
   alphaCSR[ 164 ][ 168 ],
   alphaCSR[ 164 ][ 169 ],
   alphaCSR[ 164 ][ 170 ],
   alphaCSR[ 164 ][ 171 ],
   alphaCSR[ 164 ][ 172 ],
   alphaCSR[ 164 ][ 173 ],
   alphaCSR[ 164 ][ 174 ],
   alphaCSR[ 164 ][ 175 ],
   alphaCSR[ 164 ][ 176 ],
   alphaCSR[ 164 ][ 177 ],
   alphaCSR[ 164 ][ 178 ],
   alphaCSR[ 164 ][ 179 ],
   alphaCSR[ 164 ][ 180 ],
   alphaCSR[ 164 ][ 181 ],
   alphaCSR[ 164 ][ 182 ],
   alphaCSR[ 164 ][ 183 ],
   alphaCSR[ 164 ][ 184 ],
   alphaCSR[ 164 ][ 185 ],
   alphaCSR[ 164 ][ 186 ],
   alphaCSR[ 164 ][ 187 ],
   alphaCSR[ 164 ][ 188 ],
   alphaCSR[ 164 ][ 189 ],
   alphaCSR[ 164 ][ 190 ],
   alphaCSR[ 164 ][ 191 ],
   alphaCSR[ 164 ][ 192 ],
   alphaCSR[ 164 ][ 193 ],
   alphaCSR[ 164 ][ 194 ],
   alphaCSR[ 164 ][ 195 ],
   alphaCSR[ 164 ][ 196 ],
   alphaCSR[ 164 ][ 197 ],
   alphaCSR[ 164 ][ 198 ],
   alphaCSR[ 164 ][ 199 ],
   alphaCSR[ 164 ][ 200 ],
   alphaCSR[ 164 ][ 201 ],
   alphaCSR[ 164 ][ 202 ],
   alphaCSR[ 164 ][ 203 ],
   alphaCSR[ 164 ][ 204 ],
   alphaCSR[ 164 ][ 205 ],
   alphaCSR[ 164 ][ 206 ],
   alphaCSR[ 164 ][ 207 ],
   alphaCSR[ 164 ][ 208 ],
   alphaCSR[ 164 ][ 209 ],
   alphaCSR[ 164 ][ 210 ],
   alphaCSR[ 164 ][ 211 ],
   alphaCSR[ 164 ][ 212 ],
   alphaCSR[ 164 ][ 213 ],
   alphaCSR[ 164 ][ 214 ],
   alphaCSR[ 164 ][ 215 ],
   alphaCSR[ 164 ][ 216 ],
   alphaCSR[ 164 ][ 217 ],
   alphaCSR[ 164 ][ 218 ],
   alphaCSR[ 164 ][ 219 ],
   alphaCSR[ 164 ][ 220 ],
   alphaCSR[ 164 ][ 221 ],
   alphaCSR[ 164 ][ 222 ],
   alphaCSR[ 164 ][ 223 ],
   alphaCSR[ 164 ][ 224 ],
   alphaCSR[ 164 ][ 225 ],
   alphaCSR[ 164 ][ 226 ],
   alphaCSR[ 164 ][ 227 ],
   alphaCSR[ 164 ][ 228 ],
   alphaCSR[ 164 ][ 229 ],
   alphaCSR[ 164 ][ 230 ],
   alphaCSR[ 164 ][ 231 ],
   alphaCSR[ 164 ][ 232 ],
   alphaCSR[ 164 ][ 233 ],
   alphaCSR[ 164 ][ 234 ],
   alphaCSR[ 164 ][ 235 ],
   alphaCSR[ 164 ][ 236 ],
   alphaCSR[ 164 ][ 237 ],
   alphaCSR[ 164 ][ 238 ],
   alphaCSR[ 164 ][ 239 ],
   alphaCSR[ 164 ][ 240 ],
   alphaCSR[ 164 ][ 241 ],
   alphaCSR[ 164 ][ 242 ],
   alphaCSR[ 164 ][ 243 ],
   alphaCSR[ 164 ][ 244 ],
   alphaCSR[ 164 ][ 245 ],
   alphaCSR[ 164 ][ 246 ],
   alphaCSR[ 164 ][ 247 ],
   alphaCSR[ 164 ][ 248 ],
   alphaCSR[ 164 ][ 249 ],
   alphaCSR[ 164 ][ 250 ],
   alphaCSR[ 164 ][ 251 ],
   alphaCSR[ 164 ][ 252 ],
   alphaCSR[ 164 ][ 253 ],
   alphaCSR[ 164 ][ 254 ],
   alphaCSR[ 164 ][ 255 ],
   alphaCSR[ 164 ][ 256 ],
   alphaCSR[ 164 ][ 257 ],
   alphaCSR[ 164 ][ 258 ],
   alphaCSR[ 164 ][ 259 ],
   alphaCSR[ 164 ][ 260 ],
   alphaCSR[ 164 ][ 261 ],
   alphaCSR[ 164 ][ 262 ],
   alphaCSR[ 164 ][ 263 ],
   alphaCSR[ 164 ][ 264 ],
   alphaCSR[ 164 ][ 265 ],
   alphaCSR[ 164 ][ 266 ],
   alphaCSR[ 164 ][ 267 ],
   alphaCSR[ 164 ][ 268 ],
   alphaCSR[ 164 ][ 269 ],
   alphaCSR[ 164 ][ 270 ],
   alphaCSR[ 164 ][ 271 ],
   alphaCSR[ 164 ][ 272 ],
   alphaCSR[ 164 ][ 273 ],
   alphaCSR[ 164 ][ 274 ],
   alphaCSR[ 164 ][ 275 ],
   alphaCSR[ 164 ][ 276 ],
   alphaCSR[ 164 ][ 277 ],
   alphaCSR[ 164 ][ 278 ],
   alphaCSR[ 164 ][ 279 ],
   alphaCSR[ 164 ][ 280 ],
   alphaCSR[ 164 ][ 281 ],
   alphaCSR[ 164 ][ 282 ],
   alphaCSR[ 164 ][ 283 ],
   alphaCSR[ 164 ][ 284 ],
   alphaCSR[ 164 ][ 285 ],
   alphaCSR[ 164 ][ 286 ],
   alphaCSR[ 164 ][ 287 ],
   alphaCSR[ 164 ][ 288 ],
   alphaCSR[ 164 ][ 289 ],
   alphaCSR[ 164 ][ 290 ],
   alphaCSR[ 164 ][ 291 ],
   alphaCSR[ 164 ][ 292 ],
   alphaCSR[ 164 ][ 293 ],
   alphaCSR[ 164 ][ 294 ],
   alphaCSR[ 164 ][ 295 ],
   alphaCSR[ 164 ][ 296 ],
   alphaCSR[ 164 ][ 297 ],
   alphaCSR[ 164 ][ 298 ],
   alphaCSR[ 164 ][ 299 ],
   alphaCSR[ 164 ][ 300 ],
   alphaCSR[ 164 ][ 301 ],
   alphaCSR[ 164 ][ 302 ],
   alphaCSR[ 164 ][ 303 ],
   alphaCSR[ 164 ][ 304 ],
   alphaCSR[ 164 ][ 305 ],
   alphaCSR[ 164 ][ 306 ],
   alphaCSR[ 164 ][ 307 ],
   alphaCSR[ 164 ][ 308 ],
   alphaCSR[ 164 ][ 309 ],
   alphaCSR[ 164 ][ 310 ],
   alphaCSR[ 164 ][ 311 ],
   alphaCSR[ 164 ][ 312 ],
   alphaCSR[ 164 ][ 313 ],
   alphaCSR[ 164 ][ 314 ],
   alphaCSR[ 164 ][ 315 ],
   alphaCSR[ 164 ][ 316 ],
   alphaCSR[ 164 ][ 317 ],
   alphaCSR[ 164 ][ 318 ],
   alphaCSR[ 164 ][ 319 ],
   alphaCSR[ 164 ][ 320 ],
   alphaCSR[ 164 ][ 321 ],
   alphaCSR[ 164 ][ 322 ],
   alphaCSR[ 164 ][ 323 ],
   alphaCSR[ 164 ][ 324 ],
   alphaCSR[ 164 ][ 325 ],
   alphaCSR[ 164 ][ 326 ],
   alphaCSR[ 164 ][ 327 ],
   alphaCSR[ 164 ][ 328 ],
   alphaCSR[ 164 ][ 329 ],
   alphaCSR[ 164 ][ 330 ],
   alphaCSR[ 164 ][ 331 ],
   alphaCSR[ 164 ][ 332 ],
   alphaCSR[ 164 ][ 333 ],
   alphaCSR[ 164 ][ 334 ],
   alphaCSR[ 164 ][ 335 ],
   alphaCSR[ 164 ][ 336 ],
   alphaCSR[ 164 ][ 337 ],
   alphaCSR[ 164 ][ 338 ],
   alphaCSR[ 164 ][ 339 ],
   alphaCSR[ 164 ][ 340 ],
   alphaCSR[ 164 ][ 341 ],
   alphaCSR[ 164 ][ 342 ],
   alphaCSR[ 164 ][ 343 ],
   alphaCSR[ 164 ][ 344 ],
   alphaCSR[ 164 ][ 345 ],
   alphaCSR[ 164 ][ 346 ],
   alphaCSR[ 164 ][ 347 ],
   alphaCSR[ 164 ][ 348 ],
   alphaCSR[ 164 ][ 349 ],
   alphaCSR[ 164 ][ 350 ],
   alphaCSR[ 164 ][ 351 ],
   alphaCSR[ 164 ][ 352 ],
   alphaCSR[ 164 ][ 353 ],
   alphaCSR[ 164 ][ 354 ],
   alphaCSR[ 164 ][ 355 ],
   alphaCSR[ 164 ][ 356 ],
   alphaCSR[ 164 ][ 357 ],
   alphaCSR[ 164 ][ 358 ],
   alphaCSR[ 164 ][ 359 ],
   alphaCSR[ 164 ][ 360 ],
   alphaCSR[ 164 ][ 361 ],
   alphaCSR[ 164 ][ 362 ],
   alphaCSR[ 164 ][ 363 ],
   alphaCSR[ 164 ][ 364 ],
   alphaCSR[ 164 ][ 365 ],
   alphaCSR[ 164 ][ 366 ],
   alphaCSR[ 164 ][ 367 ],
   alphaCSR[ 164 ][ 368 ],
   alphaCSR[ 164 ][ 369 ],
   alphaCSR[ 164 ][ 370 ],
   alphaCSR[ 164 ][ 371 ],
   alphaCSR[ 164 ][ 372 ],
   alphaCSR[ 164 ][ 373 ],
   alphaCSR[ 164 ][ 374 ],
   alphaCSR[ 164 ][ 375 ],
   alphaCSR[ 164 ][ 376 ],
   alphaCSR[ 164 ][ 377 ],
   alphaCSR[ 164 ][ 378 ],
   alphaCSR[ 164 ][ 379 ],
   alphaCSR[ 164 ][ 380 ],
   alphaCSR[ 164 ][ 381 ],
   alphaCSR[ 164 ][ 382 ],
   alphaCSR[ 164 ][ 383 ],
   alphaCSR[ 165 ][ 0 ],
   alphaCSR[ 165 ][ 1 ],
   alphaCSR[ 165 ][ 2 ],
   alphaCSR[ 165 ][ 3 ],
   alphaCSR[ 165 ][ 4 ],
   alphaCSR[ 165 ][ 5 ],
   alphaCSR[ 165 ][ 6 ],
   alphaCSR[ 165 ][ 7 ],
   alphaCSR[ 165 ][ 8 ],
   alphaCSR[ 165 ][ 9 ],
   alphaCSR[ 165 ][ 10 ],
   alphaCSR[ 165 ][ 11 ],
   alphaCSR[ 165 ][ 12 ],
   alphaCSR[ 165 ][ 13 ],
   alphaCSR[ 165 ][ 14 ],
   alphaCSR[ 165 ][ 15 ],
   alphaCSR[ 165 ][ 16 ],
   alphaCSR[ 165 ][ 17 ],
   alphaCSR[ 165 ][ 18 ],
   alphaCSR[ 165 ][ 19 ],
   alphaCSR[ 165 ][ 20 ],
   alphaCSR[ 165 ][ 21 ],
   alphaCSR[ 165 ][ 22 ],
   alphaCSR[ 165 ][ 23 ],
   alphaCSR[ 165 ][ 24 ],
   alphaCSR[ 165 ][ 25 ],
   alphaCSR[ 165 ][ 26 ],
   alphaCSR[ 165 ][ 27 ],
   alphaCSR[ 165 ][ 28 ],
   alphaCSR[ 165 ][ 29 ],
   alphaCSR[ 165 ][ 30 ],
   alphaCSR[ 165 ][ 31 ],
   alphaCSR[ 165 ][ 32 ],
   alphaCSR[ 165 ][ 33 ],
   alphaCSR[ 165 ][ 34 ],
   alphaCSR[ 165 ][ 35 ],
   alphaCSR[ 165 ][ 36 ],
   alphaCSR[ 165 ][ 37 ],
   alphaCSR[ 165 ][ 38 ],
   alphaCSR[ 165 ][ 39 ],
   alphaCSR[ 165 ][ 40 ],
   alphaCSR[ 165 ][ 41 ],
   alphaCSR[ 165 ][ 42 ],
   alphaCSR[ 165 ][ 43 ],
   alphaCSR[ 165 ][ 44 ],
   alphaCSR[ 165 ][ 45 ],
   alphaCSR[ 165 ][ 46 ],
   alphaCSR[ 165 ][ 47 ],
   alphaCSR[ 165 ][ 48 ],
   alphaCSR[ 165 ][ 49 ],
   alphaCSR[ 165 ][ 50 ],
   alphaCSR[ 165 ][ 51 ],
   alphaCSR[ 165 ][ 52 ],
   alphaCSR[ 165 ][ 53 ],
   alphaCSR[ 165 ][ 54 ],
   alphaCSR[ 165 ][ 55 ],
   alphaCSR[ 165 ][ 56 ],
   alphaCSR[ 165 ][ 57 ],
   alphaCSR[ 165 ][ 58 ],
   alphaCSR[ 165 ][ 59 ],
   alphaCSR[ 165 ][ 60 ],
   alphaCSR[ 165 ][ 61 ],
   alphaCSR[ 165 ][ 62 ],
   alphaCSR[ 165 ][ 63 ],
   alphaCSR[ 165 ][ 64 ],
   alphaCSR[ 165 ][ 65 ],
   alphaCSR[ 165 ][ 66 ],
   alphaCSR[ 165 ][ 67 ],
   alphaCSR[ 165 ][ 68 ],
   alphaCSR[ 165 ][ 69 ],
   alphaCSR[ 165 ][ 70 ],
   alphaCSR[ 165 ][ 71 ],
   alphaCSR[ 165 ][ 72 ],
   alphaCSR[ 165 ][ 73 ],
   alphaCSR[ 165 ][ 74 ],
   alphaCSR[ 165 ][ 75 ],
   alphaCSR[ 165 ][ 76 ],
   alphaCSR[ 165 ][ 77 ],
   alphaCSR[ 165 ][ 78 ],
   alphaCSR[ 165 ][ 79 ],
   alphaCSR[ 165 ][ 80 ],
   alphaCSR[ 165 ][ 81 ],
   alphaCSR[ 165 ][ 82 ],
   alphaCSR[ 165 ][ 83 ],
   alphaCSR[ 165 ][ 84 ],
   alphaCSR[ 165 ][ 85 ],
   alphaCSR[ 165 ][ 86 ],
   alphaCSR[ 165 ][ 87 ],
   alphaCSR[ 165 ][ 88 ],
   alphaCSR[ 165 ][ 89 ],
   alphaCSR[ 165 ][ 90 ],
   alphaCSR[ 165 ][ 91 ],
   alphaCSR[ 165 ][ 92 ],
   alphaCSR[ 165 ][ 93 ],
   alphaCSR[ 165 ][ 94 ],
   alphaCSR[ 165 ][ 95 ],
   alphaCSR[ 165 ][ 96 ],
   alphaCSR[ 165 ][ 97 ],
   alphaCSR[ 165 ][ 98 ],
   alphaCSR[ 165 ][ 99 ],
   alphaCSR[ 165 ][ 100 ],
   alphaCSR[ 165 ][ 101 ],
   alphaCSR[ 165 ][ 102 ],
   alphaCSR[ 165 ][ 103 ],
   alphaCSR[ 165 ][ 104 ],
   alphaCSR[ 165 ][ 105 ],
   alphaCSR[ 165 ][ 106 ],
   alphaCSR[ 165 ][ 107 ],
   alphaCSR[ 165 ][ 108 ],
   alphaCSR[ 165 ][ 109 ],
   alphaCSR[ 165 ][ 110 ],
   alphaCSR[ 165 ][ 111 ],
   alphaCSR[ 165 ][ 112 ],
   alphaCSR[ 165 ][ 113 ],
   alphaCSR[ 165 ][ 114 ],
   alphaCSR[ 165 ][ 115 ],
   alphaCSR[ 165 ][ 116 ],
   alphaCSR[ 165 ][ 117 ],
   alphaCSR[ 165 ][ 118 ],
   alphaCSR[ 165 ][ 119 ],
   alphaCSR[ 165 ][ 120 ],
   alphaCSR[ 165 ][ 121 ],
   alphaCSR[ 165 ][ 122 ],
   alphaCSR[ 165 ][ 123 ],
   alphaCSR[ 165 ][ 124 ],
   alphaCSR[ 165 ][ 125 ],
   alphaCSR[ 165 ][ 126 ],
   alphaCSR[ 165 ][ 127 ],
   alphaCSR[ 165 ][ 128 ],
   alphaCSR[ 165 ][ 129 ],
   alphaCSR[ 165 ][ 130 ],
   alphaCSR[ 165 ][ 131 ],
   alphaCSR[ 165 ][ 132 ],
   alphaCSR[ 165 ][ 133 ],
   alphaCSR[ 165 ][ 134 ],
   alphaCSR[ 165 ][ 135 ],
   alphaCSR[ 165 ][ 136 ],
   alphaCSR[ 165 ][ 137 ],
   alphaCSR[ 165 ][ 138 ],
   alphaCSR[ 165 ][ 139 ],
   alphaCSR[ 165 ][ 140 ],
   alphaCSR[ 165 ][ 141 ],
   alphaCSR[ 165 ][ 142 ],
   alphaCSR[ 165 ][ 143 ],
   alphaCSR[ 165 ][ 144 ],
   alphaCSR[ 165 ][ 145 ],
   alphaCSR[ 165 ][ 146 ],
   alphaCSR[ 165 ][ 147 ],
   alphaCSR[ 165 ][ 148 ],
   alphaCSR[ 165 ][ 149 ],
   alphaCSR[ 165 ][ 150 ],
   alphaCSR[ 165 ][ 151 ],
   alphaCSR[ 165 ][ 152 ],
   alphaCSR[ 165 ][ 153 ],
   alphaCSR[ 165 ][ 154 ],
   alphaCSR[ 165 ][ 155 ],
   alphaCSR[ 165 ][ 156 ],
   alphaCSR[ 165 ][ 157 ],
   alphaCSR[ 165 ][ 158 ],
   alphaCSR[ 165 ][ 159 ],
   alphaCSR[ 165 ][ 160 ],
   alphaCSR[ 165 ][ 161 ],
   alphaCSR[ 165 ][ 162 ],
   alphaCSR[ 165 ][ 163 ],
   alphaCSR[ 165 ][ 164 ],
   alphaCSR[ 165 ][ 165 ],
   alphaCSR[ 165 ][ 166 ],
   alphaCSR[ 165 ][ 167 ],
   alphaCSR[ 165 ][ 168 ],
   alphaCSR[ 165 ][ 169 ],
   alphaCSR[ 165 ][ 170 ],
   alphaCSR[ 165 ][ 171 ],
   alphaCSR[ 165 ][ 172 ],
   alphaCSR[ 165 ][ 173 ],
   alphaCSR[ 165 ][ 174 ],
   alphaCSR[ 165 ][ 175 ],
   alphaCSR[ 165 ][ 176 ],
   alphaCSR[ 165 ][ 177 ],
   alphaCSR[ 165 ][ 178 ],
   alphaCSR[ 165 ][ 179 ],
   alphaCSR[ 165 ][ 180 ],
   alphaCSR[ 165 ][ 181 ],
   alphaCSR[ 165 ][ 182 ],
   alphaCSR[ 165 ][ 183 ],
   alphaCSR[ 165 ][ 184 ],
   alphaCSR[ 165 ][ 185 ],
   alphaCSR[ 165 ][ 186 ],
   alphaCSR[ 165 ][ 187 ],
   alphaCSR[ 165 ][ 188 ],
   alphaCSR[ 165 ][ 189 ],
   alphaCSR[ 165 ][ 190 ],
   alphaCSR[ 165 ][ 191 ],
   alphaCSR[ 165 ][ 192 ],
   alphaCSR[ 165 ][ 193 ],
   alphaCSR[ 165 ][ 194 ],
   alphaCSR[ 165 ][ 195 ],
   alphaCSR[ 165 ][ 196 ],
   alphaCSR[ 165 ][ 197 ],
   alphaCSR[ 165 ][ 198 ],
   alphaCSR[ 165 ][ 199 ],
   alphaCSR[ 165 ][ 200 ],
   alphaCSR[ 165 ][ 201 ],
   alphaCSR[ 165 ][ 202 ],
   alphaCSR[ 165 ][ 203 ],
   alphaCSR[ 165 ][ 204 ],
   alphaCSR[ 165 ][ 205 ],
   alphaCSR[ 165 ][ 206 ],
   alphaCSR[ 165 ][ 207 ],
   alphaCSR[ 165 ][ 208 ],
   alphaCSR[ 165 ][ 209 ],
   alphaCSR[ 165 ][ 210 ],
   alphaCSR[ 165 ][ 211 ],
   alphaCSR[ 165 ][ 212 ],
   alphaCSR[ 165 ][ 213 ],
   alphaCSR[ 165 ][ 214 ],
   alphaCSR[ 165 ][ 215 ],
   alphaCSR[ 165 ][ 216 ],
   alphaCSR[ 165 ][ 217 ],
   alphaCSR[ 165 ][ 218 ],
   alphaCSR[ 165 ][ 219 ],
   alphaCSR[ 165 ][ 220 ],
   alphaCSR[ 165 ][ 221 ],
   alphaCSR[ 165 ][ 222 ],
   alphaCSR[ 165 ][ 223 ],
   alphaCSR[ 165 ][ 224 ],
   alphaCSR[ 165 ][ 225 ],
   alphaCSR[ 165 ][ 226 ],
   alphaCSR[ 165 ][ 227 ],
   alphaCSR[ 165 ][ 228 ],
   alphaCSR[ 165 ][ 229 ],
   alphaCSR[ 165 ][ 230 ],
   alphaCSR[ 165 ][ 231 ],
   alphaCSR[ 165 ][ 232 ],
   alphaCSR[ 165 ][ 233 ],
   alphaCSR[ 165 ][ 234 ],
   alphaCSR[ 165 ][ 235 ],
   alphaCSR[ 165 ][ 236 ],
   alphaCSR[ 165 ][ 237 ],
   alphaCSR[ 165 ][ 238 ],
   alphaCSR[ 165 ][ 239 ],
   alphaCSR[ 165 ][ 240 ],
   alphaCSR[ 165 ][ 241 ],
   alphaCSR[ 165 ][ 242 ],
   alphaCSR[ 165 ][ 243 ],
   alphaCSR[ 165 ][ 244 ],
   alphaCSR[ 165 ][ 245 ],
   alphaCSR[ 165 ][ 246 ],
   alphaCSR[ 165 ][ 247 ],
   alphaCSR[ 165 ][ 248 ],
   alphaCSR[ 165 ][ 249 ],
   alphaCSR[ 165 ][ 250 ],
   alphaCSR[ 165 ][ 251 ],
   alphaCSR[ 165 ][ 252 ],
   alphaCSR[ 165 ][ 253 ],
   alphaCSR[ 165 ][ 254 ],
   alphaCSR[ 165 ][ 255 ],
   alphaCSR[ 165 ][ 256 ],
   alphaCSR[ 165 ][ 257 ],
   alphaCSR[ 165 ][ 258 ],
   alphaCSR[ 165 ][ 259 ],
   alphaCSR[ 165 ][ 260 ],
   alphaCSR[ 165 ][ 261 ],
   alphaCSR[ 165 ][ 262 ],
   alphaCSR[ 165 ][ 263 ],
   alphaCSR[ 165 ][ 264 ],
   alphaCSR[ 165 ][ 265 ],
   alphaCSR[ 165 ][ 266 ],
   alphaCSR[ 165 ][ 267 ],
   alphaCSR[ 165 ][ 268 ],
   alphaCSR[ 165 ][ 269 ],
   alphaCSR[ 165 ][ 270 ],
   alphaCSR[ 165 ][ 271 ],
   alphaCSR[ 165 ][ 272 ],
   alphaCSR[ 165 ][ 273 ],
   alphaCSR[ 165 ][ 274 ],
   alphaCSR[ 165 ][ 275 ],
   alphaCSR[ 165 ][ 276 ],
   alphaCSR[ 165 ][ 277 ],
   alphaCSR[ 165 ][ 278 ],
   alphaCSR[ 165 ][ 279 ],
   alphaCSR[ 165 ][ 280 ],
   alphaCSR[ 165 ][ 281 ],
   alphaCSR[ 165 ][ 282 ],
   alphaCSR[ 165 ][ 283 ],
   alphaCSR[ 165 ][ 284 ],
   alphaCSR[ 165 ][ 285 ],
   alphaCSR[ 165 ][ 286 ],
   alphaCSR[ 165 ][ 287 ],
   alphaCSR[ 165 ][ 288 ],
   alphaCSR[ 165 ][ 289 ],
   alphaCSR[ 165 ][ 290 ],
   alphaCSR[ 165 ][ 291 ],
   alphaCSR[ 165 ][ 292 ],
   alphaCSR[ 165 ][ 293 ],
   alphaCSR[ 165 ][ 294 ],
   alphaCSR[ 165 ][ 295 ],
   alphaCSR[ 165 ][ 296 ],
   alphaCSR[ 165 ][ 297 ],
   alphaCSR[ 165 ][ 298 ],
   alphaCSR[ 165 ][ 299 ],
   alphaCSR[ 165 ][ 300 ],
   alphaCSR[ 165 ][ 301 ],
   alphaCSR[ 165 ][ 302 ],
   alphaCSR[ 165 ][ 303 ],
   alphaCSR[ 165 ][ 304 ],
   alphaCSR[ 165 ][ 305 ],
   alphaCSR[ 165 ][ 306 ],
   alphaCSR[ 165 ][ 307 ],
   alphaCSR[ 165 ][ 308 ],
   alphaCSR[ 165 ][ 309 ],
   alphaCSR[ 165 ][ 310 ],
   alphaCSR[ 165 ][ 311 ],
   alphaCSR[ 165 ][ 312 ],
   alphaCSR[ 165 ][ 313 ],
   alphaCSR[ 165 ][ 314 ],
   alphaCSR[ 165 ][ 315 ],
   alphaCSR[ 165 ][ 316 ],
   alphaCSR[ 165 ][ 317 ],
   alphaCSR[ 165 ][ 318 ],
   alphaCSR[ 165 ][ 319 ],
   alphaCSR[ 165 ][ 320 ],
   alphaCSR[ 165 ][ 321 ],
   alphaCSR[ 165 ][ 322 ],
   alphaCSR[ 165 ][ 323 ],
   alphaCSR[ 165 ][ 324 ],
   alphaCSR[ 165 ][ 325 ],
   alphaCSR[ 165 ][ 326 ],
   alphaCSR[ 165 ][ 327 ],
   alphaCSR[ 165 ][ 328 ],
   alphaCSR[ 165 ][ 329 ],
   alphaCSR[ 165 ][ 330 ],
   alphaCSR[ 165 ][ 331 ],
   alphaCSR[ 165 ][ 332 ],
   alphaCSR[ 165 ][ 333 ],
   alphaCSR[ 165 ][ 334 ],
   alphaCSR[ 165 ][ 335 ],
   alphaCSR[ 165 ][ 336 ],
   alphaCSR[ 165 ][ 337 ],
   alphaCSR[ 165 ][ 338 ],
   alphaCSR[ 165 ][ 339 ],
   alphaCSR[ 165 ][ 340 ],
   alphaCSR[ 165 ][ 341 ],
   alphaCSR[ 165 ][ 342 ],
   alphaCSR[ 165 ][ 343 ],
   alphaCSR[ 165 ][ 344 ],
   alphaCSR[ 165 ][ 345 ],
   alphaCSR[ 165 ][ 346 ],
   alphaCSR[ 165 ][ 347 ],
   alphaCSR[ 165 ][ 348 ],
   alphaCSR[ 165 ][ 349 ],
   alphaCSR[ 165 ][ 350 ],
   alphaCSR[ 165 ][ 351 ],
   alphaCSR[ 165 ][ 352 ],
   alphaCSR[ 165 ][ 353 ],
   alphaCSR[ 165 ][ 354 ],
   alphaCSR[ 165 ][ 355 ],
   alphaCSR[ 165 ][ 356 ],
   alphaCSR[ 165 ][ 357 ],
   alphaCSR[ 165 ][ 358 ],
   alphaCSR[ 165 ][ 359 ],
   alphaCSR[ 165 ][ 360 ],
   alphaCSR[ 165 ][ 361 ],
   alphaCSR[ 165 ][ 362 ],
   alphaCSR[ 165 ][ 363 ],
   alphaCSR[ 165 ][ 364 ],
   alphaCSR[ 165 ][ 365 ],
   alphaCSR[ 165 ][ 366 ],
   alphaCSR[ 165 ][ 367 ],
   alphaCSR[ 165 ][ 368 ],
   alphaCSR[ 165 ][ 369 ],
   alphaCSR[ 165 ][ 370 ],
   alphaCSR[ 165 ][ 371 ],
   alphaCSR[ 165 ][ 372 ],
   alphaCSR[ 165 ][ 373 ],
   alphaCSR[ 165 ][ 374 ],
   alphaCSR[ 165 ][ 375 ],
   alphaCSR[ 165 ][ 376 ],
   alphaCSR[ 165 ][ 377 ],
   alphaCSR[ 165 ][ 378 ],
   alphaCSR[ 165 ][ 379 ],
   alphaCSR[ 165 ][ 380 ],
   alphaCSR[ 165 ][ 381 ],
   alphaCSR[ 165 ][ 382 ],
   alphaCSR[ 165 ][ 383 ],
   alphaCSR[ 166 ][ 0 ],
   alphaCSR[ 166 ][ 1 ],
   alphaCSR[ 166 ][ 2 ],
   alphaCSR[ 166 ][ 3 ],
   alphaCSR[ 166 ][ 4 ],
   alphaCSR[ 166 ][ 5 ],
   alphaCSR[ 166 ][ 6 ],
   alphaCSR[ 166 ][ 7 ],
   alphaCSR[ 166 ][ 8 ],
   alphaCSR[ 166 ][ 9 ],
   alphaCSR[ 166 ][ 10 ],
   alphaCSR[ 166 ][ 11 ],
   alphaCSR[ 166 ][ 12 ],
   alphaCSR[ 166 ][ 13 ],
   alphaCSR[ 166 ][ 14 ],
   alphaCSR[ 166 ][ 15 ],
   alphaCSR[ 166 ][ 16 ],
   alphaCSR[ 166 ][ 17 ],
   alphaCSR[ 166 ][ 18 ],
   alphaCSR[ 166 ][ 19 ],
   alphaCSR[ 166 ][ 20 ],
   alphaCSR[ 166 ][ 21 ],
   alphaCSR[ 166 ][ 22 ],
   alphaCSR[ 166 ][ 23 ],
   alphaCSR[ 166 ][ 24 ],
   alphaCSR[ 166 ][ 25 ],
   alphaCSR[ 166 ][ 26 ],
   alphaCSR[ 166 ][ 27 ],
   alphaCSR[ 166 ][ 28 ],
   alphaCSR[ 166 ][ 29 ],
   alphaCSR[ 166 ][ 30 ],
   alphaCSR[ 166 ][ 31 ],
   alphaCSR[ 166 ][ 32 ],
   alphaCSR[ 166 ][ 33 ],
   alphaCSR[ 166 ][ 34 ],
   alphaCSR[ 166 ][ 35 ],
   alphaCSR[ 166 ][ 36 ],
   alphaCSR[ 166 ][ 37 ],
   alphaCSR[ 166 ][ 38 ],
   alphaCSR[ 166 ][ 39 ],
   alphaCSR[ 166 ][ 40 ],
   alphaCSR[ 166 ][ 41 ],
   alphaCSR[ 166 ][ 42 ],
   alphaCSR[ 166 ][ 43 ],
   alphaCSR[ 166 ][ 44 ],
   alphaCSR[ 166 ][ 45 ],
   alphaCSR[ 166 ][ 46 ],
   alphaCSR[ 166 ][ 47 ],
   alphaCSR[ 166 ][ 48 ],
   alphaCSR[ 166 ][ 49 ],
   alphaCSR[ 166 ][ 50 ],
   alphaCSR[ 166 ][ 51 ],
   alphaCSR[ 166 ][ 52 ],
   alphaCSR[ 166 ][ 53 ],
   alphaCSR[ 166 ][ 54 ],
   alphaCSR[ 166 ][ 55 ],
   alphaCSR[ 166 ][ 56 ],
   alphaCSR[ 166 ][ 57 ],
   alphaCSR[ 166 ][ 58 ],
   alphaCSR[ 166 ][ 59 ],
   alphaCSR[ 166 ][ 60 ],
   alphaCSR[ 166 ][ 61 ],
   alphaCSR[ 166 ][ 62 ],
   alphaCSR[ 166 ][ 63 ],
   alphaCSR[ 166 ][ 64 ],
   alphaCSR[ 166 ][ 65 ],
   alphaCSR[ 166 ][ 66 ],
   alphaCSR[ 166 ][ 67 ],
   alphaCSR[ 166 ][ 68 ],
   alphaCSR[ 166 ][ 69 ],
   alphaCSR[ 166 ][ 70 ],
   alphaCSR[ 166 ][ 71 ],
   alphaCSR[ 166 ][ 72 ],
   alphaCSR[ 166 ][ 73 ],
   alphaCSR[ 166 ][ 74 ],
   alphaCSR[ 166 ][ 75 ],
   alphaCSR[ 166 ][ 76 ],
   alphaCSR[ 166 ][ 77 ],
   alphaCSR[ 166 ][ 78 ],
   alphaCSR[ 166 ][ 79 ],
   alphaCSR[ 166 ][ 80 ],
   alphaCSR[ 166 ][ 81 ],
   alphaCSR[ 166 ][ 82 ],
   alphaCSR[ 166 ][ 83 ],
   alphaCSR[ 166 ][ 84 ],
   alphaCSR[ 166 ][ 85 ],
   alphaCSR[ 166 ][ 86 ],
   alphaCSR[ 166 ][ 87 ],
   alphaCSR[ 166 ][ 88 ],
   alphaCSR[ 166 ][ 89 ],
   alphaCSR[ 166 ][ 90 ],
   alphaCSR[ 166 ][ 91 ],
   alphaCSR[ 166 ][ 92 ],
   alphaCSR[ 166 ][ 93 ],
   alphaCSR[ 166 ][ 94 ],
   alphaCSR[ 166 ][ 95 ],
   alphaCSR[ 166 ][ 96 ],
   alphaCSR[ 166 ][ 97 ],
   alphaCSR[ 166 ][ 98 ],
   alphaCSR[ 166 ][ 99 ],
   alphaCSR[ 166 ][ 100 ],
   alphaCSR[ 166 ][ 101 ],
   alphaCSR[ 166 ][ 102 ],
   alphaCSR[ 166 ][ 103 ],
   alphaCSR[ 166 ][ 104 ],
   alphaCSR[ 166 ][ 105 ],
   alphaCSR[ 166 ][ 106 ],
   alphaCSR[ 166 ][ 107 ],
   alphaCSR[ 166 ][ 108 ],
   alphaCSR[ 166 ][ 109 ],
   alphaCSR[ 166 ][ 110 ],
   alphaCSR[ 166 ][ 111 ],
   alphaCSR[ 166 ][ 112 ],
   alphaCSR[ 166 ][ 113 ],
   alphaCSR[ 166 ][ 114 ],
   alphaCSR[ 166 ][ 115 ],
   alphaCSR[ 166 ][ 116 ],
   alphaCSR[ 166 ][ 117 ],
   alphaCSR[ 166 ][ 118 ],
   alphaCSR[ 166 ][ 119 ],
   alphaCSR[ 166 ][ 120 ],
   alphaCSR[ 166 ][ 121 ],
   alphaCSR[ 166 ][ 122 ],
   alphaCSR[ 166 ][ 123 ],
   alphaCSR[ 166 ][ 124 ],
   alphaCSR[ 166 ][ 125 ],
   alphaCSR[ 166 ][ 126 ],
   alphaCSR[ 166 ][ 127 ],
   alphaCSR[ 166 ][ 128 ],
   alphaCSR[ 166 ][ 129 ],
   alphaCSR[ 166 ][ 130 ],
   alphaCSR[ 166 ][ 131 ],
   alphaCSR[ 166 ][ 132 ],
   alphaCSR[ 166 ][ 133 ],
   alphaCSR[ 166 ][ 134 ],
   alphaCSR[ 166 ][ 135 ],
   alphaCSR[ 166 ][ 136 ],
   alphaCSR[ 166 ][ 137 ],
   alphaCSR[ 166 ][ 138 ],
   alphaCSR[ 166 ][ 139 ],
   alphaCSR[ 166 ][ 140 ],
   alphaCSR[ 166 ][ 141 ],
   alphaCSR[ 166 ][ 142 ],
   alphaCSR[ 166 ][ 143 ],
   alphaCSR[ 166 ][ 144 ],
   alphaCSR[ 166 ][ 145 ],
   alphaCSR[ 166 ][ 146 ],
   alphaCSR[ 166 ][ 147 ],
   alphaCSR[ 166 ][ 148 ],
   alphaCSR[ 166 ][ 149 ],
   alphaCSR[ 166 ][ 150 ],
   alphaCSR[ 166 ][ 151 ],
   alphaCSR[ 166 ][ 152 ],
   alphaCSR[ 166 ][ 153 ],
   alphaCSR[ 166 ][ 154 ],
   alphaCSR[ 166 ][ 155 ],
   alphaCSR[ 166 ][ 156 ],
   alphaCSR[ 166 ][ 157 ],
   alphaCSR[ 166 ][ 158 ],
   alphaCSR[ 166 ][ 159 ],
   alphaCSR[ 166 ][ 160 ],
   alphaCSR[ 166 ][ 161 ],
   alphaCSR[ 166 ][ 162 ],
   alphaCSR[ 166 ][ 163 ],
   alphaCSR[ 166 ][ 164 ],
   alphaCSR[ 166 ][ 165 ],
   alphaCSR[ 166 ][ 166 ],
   alphaCSR[ 166 ][ 167 ],
   alphaCSR[ 166 ][ 168 ],
   alphaCSR[ 166 ][ 169 ],
   alphaCSR[ 166 ][ 170 ],
   alphaCSR[ 166 ][ 171 ],
   alphaCSR[ 166 ][ 172 ],
   alphaCSR[ 166 ][ 173 ],
   alphaCSR[ 166 ][ 174 ],
   alphaCSR[ 166 ][ 175 ],
   alphaCSR[ 166 ][ 176 ],
   alphaCSR[ 166 ][ 177 ],
   alphaCSR[ 166 ][ 178 ],
   alphaCSR[ 166 ][ 179 ],
   alphaCSR[ 166 ][ 180 ],
   alphaCSR[ 166 ][ 181 ],
   alphaCSR[ 166 ][ 182 ],
   alphaCSR[ 166 ][ 183 ],
   alphaCSR[ 166 ][ 184 ],
   alphaCSR[ 166 ][ 185 ],
   alphaCSR[ 166 ][ 186 ],
   alphaCSR[ 166 ][ 187 ],
   alphaCSR[ 166 ][ 188 ],
   alphaCSR[ 166 ][ 189 ],
   alphaCSR[ 166 ][ 190 ],
   alphaCSR[ 166 ][ 191 ],
   alphaCSR[ 166 ][ 192 ],
   alphaCSR[ 166 ][ 193 ],
   alphaCSR[ 166 ][ 194 ],
   alphaCSR[ 166 ][ 195 ],
   alphaCSR[ 166 ][ 196 ],
   alphaCSR[ 166 ][ 197 ],
   alphaCSR[ 166 ][ 198 ],
   alphaCSR[ 166 ][ 199 ],
   alphaCSR[ 166 ][ 200 ],
   alphaCSR[ 166 ][ 201 ],
   alphaCSR[ 166 ][ 202 ],
   alphaCSR[ 166 ][ 203 ],
   alphaCSR[ 166 ][ 204 ],
   alphaCSR[ 166 ][ 205 ],
   alphaCSR[ 166 ][ 206 ],
   alphaCSR[ 166 ][ 207 ],
   alphaCSR[ 166 ][ 208 ],
   alphaCSR[ 166 ][ 209 ],
   alphaCSR[ 166 ][ 210 ],
   alphaCSR[ 166 ][ 211 ],
   alphaCSR[ 166 ][ 212 ],
   alphaCSR[ 166 ][ 213 ],
   alphaCSR[ 166 ][ 214 ],
   alphaCSR[ 166 ][ 215 ],
   alphaCSR[ 166 ][ 216 ],
   alphaCSR[ 166 ][ 217 ],
   alphaCSR[ 166 ][ 218 ],
   alphaCSR[ 166 ][ 219 ],
   alphaCSR[ 166 ][ 220 ],
   alphaCSR[ 166 ][ 221 ],
   alphaCSR[ 166 ][ 222 ],
   alphaCSR[ 166 ][ 223 ],
   alphaCSR[ 166 ][ 224 ],
   alphaCSR[ 166 ][ 225 ],
   alphaCSR[ 166 ][ 226 ],
   alphaCSR[ 166 ][ 227 ],
   alphaCSR[ 166 ][ 228 ],
   alphaCSR[ 166 ][ 229 ],
   alphaCSR[ 166 ][ 230 ],
   alphaCSR[ 166 ][ 231 ],
   alphaCSR[ 166 ][ 232 ],
   alphaCSR[ 166 ][ 233 ],
   alphaCSR[ 166 ][ 234 ],
   alphaCSR[ 166 ][ 235 ],
   alphaCSR[ 166 ][ 236 ],
   alphaCSR[ 166 ][ 237 ],
   alphaCSR[ 166 ][ 238 ],
   alphaCSR[ 166 ][ 239 ],
   alphaCSR[ 166 ][ 240 ],
   alphaCSR[ 166 ][ 241 ],
   alphaCSR[ 166 ][ 242 ],
   alphaCSR[ 166 ][ 243 ],
   alphaCSR[ 166 ][ 244 ],
   alphaCSR[ 166 ][ 245 ],
   alphaCSR[ 166 ][ 246 ],
   alphaCSR[ 166 ][ 247 ],
   alphaCSR[ 166 ][ 248 ],
   alphaCSR[ 166 ][ 249 ],
   alphaCSR[ 166 ][ 250 ],
   alphaCSR[ 166 ][ 251 ],
   alphaCSR[ 166 ][ 252 ],
   alphaCSR[ 166 ][ 253 ],
   alphaCSR[ 166 ][ 254 ],
   alphaCSR[ 166 ][ 255 ],
   alphaCSR[ 166 ][ 256 ],
   alphaCSR[ 166 ][ 257 ],
   alphaCSR[ 166 ][ 258 ],
   alphaCSR[ 166 ][ 259 ],
   alphaCSR[ 166 ][ 260 ],
   alphaCSR[ 166 ][ 261 ],
   alphaCSR[ 166 ][ 262 ],
   alphaCSR[ 166 ][ 263 ],
   alphaCSR[ 166 ][ 264 ],
   alphaCSR[ 166 ][ 265 ],
   alphaCSR[ 166 ][ 266 ],
   alphaCSR[ 166 ][ 267 ],
   alphaCSR[ 166 ][ 268 ],
   alphaCSR[ 166 ][ 269 ],
   alphaCSR[ 166 ][ 270 ],
   alphaCSR[ 166 ][ 271 ],
   alphaCSR[ 166 ][ 272 ],
   alphaCSR[ 166 ][ 273 ],
   alphaCSR[ 166 ][ 274 ],
   alphaCSR[ 166 ][ 275 ],
   alphaCSR[ 166 ][ 276 ],
   alphaCSR[ 166 ][ 277 ],
   alphaCSR[ 166 ][ 278 ],
   alphaCSR[ 166 ][ 279 ],
   alphaCSR[ 166 ][ 280 ],
   alphaCSR[ 166 ][ 281 ],
   alphaCSR[ 166 ][ 282 ],
   alphaCSR[ 166 ][ 283 ],
   alphaCSR[ 166 ][ 284 ],
   alphaCSR[ 166 ][ 285 ],
   alphaCSR[ 166 ][ 286 ],
   alphaCSR[ 166 ][ 287 ],
   alphaCSR[ 166 ][ 288 ],
   alphaCSR[ 166 ][ 289 ],
   alphaCSR[ 166 ][ 290 ],
   alphaCSR[ 166 ][ 291 ],
   alphaCSR[ 166 ][ 292 ],
   alphaCSR[ 166 ][ 293 ],
   alphaCSR[ 166 ][ 294 ],
   alphaCSR[ 166 ][ 295 ],
   alphaCSR[ 166 ][ 296 ],
   alphaCSR[ 166 ][ 297 ],
   alphaCSR[ 166 ][ 298 ],
   alphaCSR[ 166 ][ 299 ],
   alphaCSR[ 166 ][ 300 ],
   alphaCSR[ 166 ][ 301 ],
   alphaCSR[ 166 ][ 302 ],
   alphaCSR[ 166 ][ 303 ],
   alphaCSR[ 166 ][ 304 ],
   alphaCSR[ 166 ][ 305 ],
   alphaCSR[ 166 ][ 306 ],
   alphaCSR[ 166 ][ 307 ],
   alphaCSR[ 166 ][ 308 ],
   alphaCSR[ 166 ][ 309 ],
   alphaCSR[ 166 ][ 310 ],
   alphaCSR[ 166 ][ 311 ],
   alphaCSR[ 166 ][ 312 ],
   alphaCSR[ 166 ][ 313 ],
   alphaCSR[ 166 ][ 314 ],
   alphaCSR[ 166 ][ 315 ],
   alphaCSR[ 166 ][ 316 ],
   alphaCSR[ 166 ][ 317 ],
   alphaCSR[ 166 ][ 318 ],
   alphaCSR[ 166 ][ 319 ],
   alphaCSR[ 166 ][ 320 ],
   alphaCSR[ 166 ][ 321 ],
   alphaCSR[ 166 ][ 322 ],
   alphaCSR[ 166 ][ 323 ],
   alphaCSR[ 166 ][ 324 ],
   alphaCSR[ 166 ][ 325 ],
   alphaCSR[ 166 ][ 326 ],
   alphaCSR[ 166 ][ 327 ],
   alphaCSR[ 166 ][ 328 ],
   alphaCSR[ 166 ][ 329 ],
   alphaCSR[ 166 ][ 330 ],
   alphaCSR[ 166 ][ 331 ],
   alphaCSR[ 166 ][ 332 ],
   alphaCSR[ 166 ][ 333 ],
   alphaCSR[ 166 ][ 334 ],
   alphaCSR[ 166 ][ 335 ],
   alphaCSR[ 166 ][ 336 ],
   alphaCSR[ 166 ][ 337 ],
   alphaCSR[ 166 ][ 338 ],
   alphaCSR[ 166 ][ 339 ],
   alphaCSR[ 166 ][ 340 ],
   alphaCSR[ 166 ][ 341 ],
   alphaCSR[ 166 ][ 342 ],
   alphaCSR[ 166 ][ 343 ],
   alphaCSR[ 166 ][ 344 ],
   alphaCSR[ 166 ][ 345 ],
   alphaCSR[ 166 ][ 346 ],
   alphaCSR[ 166 ][ 347 ],
   alphaCSR[ 166 ][ 348 ],
   alphaCSR[ 166 ][ 349 ],
   alphaCSR[ 166 ][ 350 ],
   alphaCSR[ 166 ][ 351 ],
   alphaCSR[ 166 ][ 352 ],
   alphaCSR[ 166 ][ 353 ],
   alphaCSR[ 166 ][ 354 ],
   alphaCSR[ 166 ][ 355 ],
   alphaCSR[ 166 ][ 356 ],
   alphaCSR[ 166 ][ 357 ],
   alphaCSR[ 166 ][ 358 ],
   alphaCSR[ 166 ][ 359 ],
   alphaCSR[ 166 ][ 360 ],
   alphaCSR[ 166 ][ 361 ],
   alphaCSR[ 166 ][ 362 ],
   alphaCSR[ 166 ][ 363 ],
   alphaCSR[ 166 ][ 364 ],
   alphaCSR[ 166 ][ 365 ],
   alphaCSR[ 166 ][ 366 ],
   alphaCSR[ 166 ][ 367 ],
   alphaCSR[ 166 ][ 368 ],
   alphaCSR[ 166 ][ 369 ],
   alphaCSR[ 166 ][ 370 ],
   alphaCSR[ 166 ][ 371 ],
   alphaCSR[ 166 ][ 372 ],
   alphaCSR[ 166 ][ 373 ],
   alphaCSR[ 166 ][ 374 ],
   alphaCSR[ 166 ][ 375 ],
   alphaCSR[ 166 ][ 376 ],
   alphaCSR[ 166 ][ 377 ],
   alphaCSR[ 166 ][ 378 ],
   alphaCSR[ 166 ][ 379 ],
   alphaCSR[ 166 ][ 380 ],
   alphaCSR[ 166 ][ 381 ],
   alphaCSR[ 166 ][ 382 ],
   alphaCSR[ 166 ][ 383 ],
   alphaCSR[ 167 ][ 0 ],
   alphaCSR[ 167 ][ 1 ],
   alphaCSR[ 167 ][ 2 ],
   alphaCSR[ 167 ][ 3 ],
   alphaCSR[ 167 ][ 4 ],
   alphaCSR[ 167 ][ 5 ],
   alphaCSR[ 167 ][ 6 ],
   alphaCSR[ 167 ][ 7 ],
   alphaCSR[ 167 ][ 8 ],
   alphaCSR[ 167 ][ 9 ],
   alphaCSR[ 167 ][ 10 ],
   alphaCSR[ 167 ][ 11 ],
   alphaCSR[ 167 ][ 12 ],
   alphaCSR[ 167 ][ 13 ],
   alphaCSR[ 167 ][ 14 ],
   alphaCSR[ 167 ][ 15 ],
   alphaCSR[ 167 ][ 16 ],
   alphaCSR[ 167 ][ 17 ],
   alphaCSR[ 167 ][ 18 ],
   alphaCSR[ 167 ][ 19 ],
   alphaCSR[ 167 ][ 20 ],
   alphaCSR[ 167 ][ 21 ],
   alphaCSR[ 167 ][ 22 ],
   alphaCSR[ 167 ][ 23 ],
   alphaCSR[ 167 ][ 24 ],
   alphaCSR[ 167 ][ 25 ],
   alphaCSR[ 167 ][ 26 ],
   alphaCSR[ 167 ][ 27 ],
   alphaCSR[ 167 ][ 28 ],
   alphaCSR[ 167 ][ 29 ],
   alphaCSR[ 167 ][ 30 ],
   alphaCSR[ 167 ][ 31 ],
   alphaCSR[ 167 ][ 32 ],
   alphaCSR[ 167 ][ 33 ],
   alphaCSR[ 167 ][ 34 ],
   alphaCSR[ 167 ][ 35 ],
   alphaCSR[ 167 ][ 36 ],
   alphaCSR[ 167 ][ 37 ],
   alphaCSR[ 167 ][ 38 ],
   alphaCSR[ 167 ][ 39 ],
   alphaCSR[ 167 ][ 40 ],
   alphaCSR[ 167 ][ 41 ],
   alphaCSR[ 167 ][ 42 ],
   alphaCSR[ 167 ][ 43 ],
   alphaCSR[ 167 ][ 44 ],
   alphaCSR[ 167 ][ 45 ],
   alphaCSR[ 167 ][ 46 ],
   alphaCSR[ 167 ][ 47 ],
   alphaCSR[ 167 ][ 48 ],
   alphaCSR[ 167 ][ 49 ],
   alphaCSR[ 167 ][ 50 ],
   alphaCSR[ 167 ][ 51 ],
   alphaCSR[ 167 ][ 52 ],
   alphaCSR[ 167 ][ 53 ],
   alphaCSR[ 167 ][ 54 ],
   alphaCSR[ 167 ][ 55 ],
   alphaCSR[ 167 ][ 56 ],
   alphaCSR[ 167 ][ 57 ],
   alphaCSR[ 167 ][ 58 ],
   alphaCSR[ 167 ][ 59 ],
   alphaCSR[ 167 ][ 60 ],
   alphaCSR[ 167 ][ 61 ],
   alphaCSR[ 167 ][ 62 ],
   alphaCSR[ 167 ][ 63 ],
   alphaCSR[ 167 ][ 64 ],
   alphaCSR[ 167 ][ 65 ],
   alphaCSR[ 167 ][ 66 ],
   alphaCSR[ 167 ][ 67 ],
   alphaCSR[ 167 ][ 68 ],
   alphaCSR[ 167 ][ 69 ],
   alphaCSR[ 167 ][ 70 ],
   alphaCSR[ 167 ][ 71 ],
   alphaCSR[ 167 ][ 72 ],
   alphaCSR[ 167 ][ 73 ],
   alphaCSR[ 167 ][ 74 ],
   alphaCSR[ 167 ][ 75 ],
   alphaCSR[ 167 ][ 76 ],
   alphaCSR[ 167 ][ 77 ],
   alphaCSR[ 167 ][ 78 ],
   alphaCSR[ 167 ][ 79 ],
   alphaCSR[ 167 ][ 80 ],
   alphaCSR[ 167 ][ 81 ],
   alphaCSR[ 167 ][ 82 ],
   alphaCSR[ 167 ][ 83 ],
   alphaCSR[ 167 ][ 84 ],
   alphaCSR[ 167 ][ 85 ],
   alphaCSR[ 167 ][ 86 ],
   alphaCSR[ 167 ][ 87 ],
   alphaCSR[ 167 ][ 88 ],
   alphaCSR[ 167 ][ 89 ],
   alphaCSR[ 167 ][ 90 ],
   alphaCSR[ 167 ][ 91 ],
   alphaCSR[ 167 ][ 92 ],
   alphaCSR[ 167 ][ 93 ],
   alphaCSR[ 167 ][ 94 ],
   alphaCSR[ 167 ][ 95 ],
   alphaCSR[ 167 ][ 96 ],
   alphaCSR[ 167 ][ 97 ],
   alphaCSR[ 167 ][ 98 ],
   alphaCSR[ 167 ][ 99 ],
   alphaCSR[ 167 ][ 100 ],
   alphaCSR[ 167 ][ 101 ],
   alphaCSR[ 167 ][ 102 ],
   alphaCSR[ 167 ][ 103 ],
   alphaCSR[ 167 ][ 104 ],
   alphaCSR[ 167 ][ 105 ],
   alphaCSR[ 167 ][ 106 ],
   alphaCSR[ 167 ][ 107 ],
   alphaCSR[ 167 ][ 108 ],
   alphaCSR[ 167 ][ 109 ],
   alphaCSR[ 167 ][ 110 ],
   alphaCSR[ 167 ][ 111 ],
   alphaCSR[ 167 ][ 112 ],
   alphaCSR[ 167 ][ 113 ],
   alphaCSR[ 167 ][ 114 ],
   alphaCSR[ 167 ][ 115 ],
   alphaCSR[ 167 ][ 116 ],
   alphaCSR[ 167 ][ 117 ],
   alphaCSR[ 167 ][ 118 ],
   alphaCSR[ 167 ][ 119 ],
   alphaCSR[ 167 ][ 120 ],
   alphaCSR[ 167 ][ 121 ],
   alphaCSR[ 167 ][ 122 ],
   alphaCSR[ 167 ][ 123 ],
   alphaCSR[ 167 ][ 124 ],
   alphaCSR[ 167 ][ 125 ],
   alphaCSR[ 167 ][ 126 ],
   alphaCSR[ 167 ][ 127 ],
   alphaCSR[ 167 ][ 128 ],
   alphaCSR[ 167 ][ 129 ],
   alphaCSR[ 167 ][ 130 ],
   alphaCSR[ 167 ][ 131 ],
   alphaCSR[ 167 ][ 132 ],
   alphaCSR[ 167 ][ 133 ],
   alphaCSR[ 167 ][ 134 ],
   alphaCSR[ 167 ][ 135 ],
   alphaCSR[ 167 ][ 136 ],
   alphaCSR[ 167 ][ 137 ],
   alphaCSR[ 167 ][ 138 ],
   alphaCSR[ 167 ][ 139 ],
   alphaCSR[ 167 ][ 140 ],
   alphaCSR[ 167 ][ 141 ],
   alphaCSR[ 167 ][ 142 ],
   alphaCSR[ 167 ][ 143 ],
   alphaCSR[ 167 ][ 144 ],
   alphaCSR[ 167 ][ 145 ],
   alphaCSR[ 167 ][ 146 ],
   alphaCSR[ 167 ][ 147 ],
   alphaCSR[ 167 ][ 148 ],
   alphaCSR[ 167 ][ 149 ],
   alphaCSR[ 167 ][ 150 ],
   alphaCSR[ 167 ][ 151 ],
   alphaCSR[ 167 ][ 152 ],
   alphaCSR[ 167 ][ 153 ],
   alphaCSR[ 167 ][ 154 ],
   alphaCSR[ 167 ][ 155 ],
   alphaCSR[ 167 ][ 156 ],
   alphaCSR[ 167 ][ 157 ],
   alphaCSR[ 167 ][ 158 ],
   alphaCSR[ 167 ][ 159 ],
   alphaCSR[ 167 ][ 160 ],
   alphaCSR[ 167 ][ 161 ],
   alphaCSR[ 167 ][ 162 ],
   alphaCSR[ 167 ][ 163 ],
   alphaCSR[ 167 ][ 164 ],
   alphaCSR[ 167 ][ 165 ],
   alphaCSR[ 167 ][ 166 ],
   alphaCSR[ 167 ][ 167 ],
   alphaCSR[ 167 ][ 168 ],
   alphaCSR[ 167 ][ 169 ],
   alphaCSR[ 167 ][ 170 ],
   alphaCSR[ 167 ][ 171 ],
   alphaCSR[ 167 ][ 172 ],
   alphaCSR[ 167 ][ 173 ],
   alphaCSR[ 167 ][ 174 ],
   alphaCSR[ 167 ][ 175 ],
   alphaCSR[ 167 ][ 176 ],
   alphaCSR[ 167 ][ 177 ],
   alphaCSR[ 167 ][ 178 ],
   alphaCSR[ 167 ][ 179 ],
   alphaCSR[ 167 ][ 180 ],
   alphaCSR[ 167 ][ 181 ],
   alphaCSR[ 167 ][ 182 ],
   alphaCSR[ 167 ][ 183 ],
   alphaCSR[ 167 ][ 184 ],
   alphaCSR[ 167 ][ 185 ],
   alphaCSR[ 167 ][ 186 ],
   alphaCSR[ 167 ][ 187 ],
   alphaCSR[ 167 ][ 188 ],
   alphaCSR[ 167 ][ 189 ],
   alphaCSR[ 167 ][ 190 ],
   alphaCSR[ 167 ][ 191 ],
   alphaCSR[ 167 ][ 192 ],
   alphaCSR[ 167 ][ 193 ],
   alphaCSR[ 167 ][ 194 ],
   alphaCSR[ 167 ][ 195 ],
   alphaCSR[ 167 ][ 196 ],
   alphaCSR[ 167 ][ 197 ],
   alphaCSR[ 167 ][ 198 ],
   alphaCSR[ 167 ][ 199 ],
   alphaCSR[ 167 ][ 200 ],
   alphaCSR[ 167 ][ 201 ],
   alphaCSR[ 167 ][ 202 ],
   alphaCSR[ 167 ][ 203 ],
   alphaCSR[ 167 ][ 204 ],
   alphaCSR[ 167 ][ 205 ],
   alphaCSR[ 167 ][ 206 ],
   alphaCSR[ 167 ][ 207 ],
   alphaCSR[ 167 ][ 208 ],
   alphaCSR[ 167 ][ 209 ],
   alphaCSR[ 167 ][ 210 ],
   alphaCSR[ 167 ][ 211 ],
   alphaCSR[ 167 ][ 212 ],
   alphaCSR[ 167 ][ 213 ],
   alphaCSR[ 167 ][ 214 ],
   alphaCSR[ 167 ][ 215 ],
   alphaCSR[ 167 ][ 216 ],
   alphaCSR[ 167 ][ 217 ],
   alphaCSR[ 167 ][ 218 ],
   alphaCSR[ 167 ][ 219 ],
   alphaCSR[ 167 ][ 220 ],
   alphaCSR[ 167 ][ 221 ],
   alphaCSR[ 167 ][ 222 ],
   alphaCSR[ 167 ][ 223 ],
   alphaCSR[ 167 ][ 224 ],
   alphaCSR[ 167 ][ 225 ],
   alphaCSR[ 167 ][ 226 ],
   alphaCSR[ 167 ][ 227 ],
   alphaCSR[ 167 ][ 228 ],
   alphaCSR[ 167 ][ 229 ],
   alphaCSR[ 167 ][ 230 ],
   alphaCSR[ 167 ][ 231 ],
   alphaCSR[ 167 ][ 232 ],
   alphaCSR[ 167 ][ 233 ],
   alphaCSR[ 167 ][ 234 ],
   alphaCSR[ 167 ][ 235 ],
   alphaCSR[ 167 ][ 236 ],
   alphaCSR[ 167 ][ 237 ],
   alphaCSR[ 167 ][ 238 ],
   alphaCSR[ 167 ][ 239 ],
   alphaCSR[ 167 ][ 240 ],
   alphaCSR[ 167 ][ 241 ],
   alphaCSR[ 167 ][ 242 ],
   alphaCSR[ 167 ][ 243 ],
   alphaCSR[ 167 ][ 244 ],
   alphaCSR[ 167 ][ 245 ],
   alphaCSR[ 167 ][ 246 ],
   alphaCSR[ 167 ][ 247 ],
   alphaCSR[ 167 ][ 248 ],
   alphaCSR[ 167 ][ 249 ],
   alphaCSR[ 167 ][ 250 ],
   alphaCSR[ 167 ][ 251 ],
   alphaCSR[ 167 ][ 252 ],
   alphaCSR[ 167 ][ 253 ],
   alphaCSR[ 167 ][ 254 ],
   alphaCSR[ 167 ][ 255 ],
   alphaCSR[ 167 ][ 256 ],
   alphaCSR[ 167 ][ 257 ],
   alphaCSR[ 167 ][ 258 ],
   alphaCSR[ 167 ][ 259 ],
   alphaCSR[ 167 ][ 260 ],
   alphaCSR[ 167 ][ 261 ],
   alphaCSR[ 167 ][ 262 ],
   alphaCSR[ 167 ][ 263 ],
   alphaCSR[ 167 ][ 264 ],
   alphaCSR[ 167 ][ 265 ],
   alphaCSR[ 167 ][ 266 ],
   alphaCSR[ 167 ][ 267 ],
   alphaCSR[ 167 ][ 268 ],
   alphaCSR[ 167 ][ 269 ],
   alphaCSR[ 167 ][ 270 ],
   alphaCSR[ 167 ][ 271 ],
   alphaCSR[ 167 ][ 272 ],
   alphaCSR[ 167 ][ 273 ],
   alphaCSR[ 167 ][ 274 ],
   alphaCSR[ 167 ][ 275 ],
   alphaCSR[ 167 ][ 276 ],
   alphaCSR[ 167 ][ 277 ],
   alphaCSR[ 167 ][ 278 ],
   alphaCSR[ 167 ][ 279 ],
   alphaCSR[ 167 ][ 280 ],
   alphaCSR[ 167 ][ 281 ],
   alphaCSR[ 167 ][ 282 ],
   alphaCSR[ 167 ][ 283 ],
   alphaCSR[ 167 ][ 284 ],
   alphaCSR[ 167 ][ 285 ],
   alphaCSR[ 167 ][ 286 ],
   alphaCSR[ 167 ][ 287 ],
   alphaCSR[ 167 ][ 288 ],
   alphaCSR[ 167 ][ 289 ],
   alphaCSR[ 167 ][ 290 ],
   alphaCSR[ 167 ][ 291 ],
   alphaCSR[ 167 ][ 292 ],
   alphaCSR[ 167 ][ 293 ],
   alphaCSR[ 167 ][ 294 ],
   alphaCSR[ 167 ][ 295 ],
   alphaCSR[ 167 ][ 296 ],
   alphaCSR[ 167 ][ 297 ],
   alphaCSR[ 167 ][ 298 ],
   alphaCSR[ 167 ][ 299 ],
   alphaCSR[ 167 ][ 300 ],
   alphaCSR[ 167 ][ 301 ],
   alphaCSR[ 167 ][ 302 ],
   alphaCSR[ 167 ][ 303 ],
   alphaCSR[ 167 ][ 304 ],
   alphaCSR[ 167 ][ 305 ],
   alphaCSR[ 167 ][ 306 ],
   alphaCSR[ 167 ][ 307 ],
   alphaCSR[ 167 ][ 308 ],
   alphaCSR[ 167 ][ 309 ],
   alphaCSR[ 167 ][ 310 ],
   alphaCSR[ 167 ][ 311 ],
   alphaCSR[ 167 ][ 312 ],
   alphaCSR[ 167 ][ 313 ],
   alphaCSR[ 167 ][ 314 ],
   alphaCSR[ 167 ][ 315 ],
   alphaCSR[ 167 ][ 316 ],
   alphaCSR[ 167 ][ 317 ],
   alphaCSR[ 167 ][ 318 ],
   alphaCSR[ 167 ][ 319 ],
   alphaCSR[ 167 ][ 320 ],
   alphaCSR[ 167 ][ 321 ],
   alphaCSR[ 167 ][ 322 ],
   alphaCSR[ 167 ][ 323 ],
   alphaCSR[ 167 ][ 324 ],
   alphaCSR[ 167 ][ 325 ],
   alphaCSR[ 167 ][ 326 ],
   alphaCSR[ 167 ][ 327 ],
   alphaCSR[ 167 ][ 328 ],
   alphaCSR[ 167 ][ 329 ],
   alphaCSR[ 167 ][ 330 ],
   alphaCSR[ 167 ][ 331 ],
   alphaCSR[ 167 ][ 332 ],
   alphaCSR[ 167 ][ 333 ],
   alphaCSR[ 167 ][ 334 ],
   alphaCSR[ 167 ][ 335 ],
   alphaCSR[ 167 ][ 336 ],
   alphaCSR[ 167 ][ 337 ],
   alphaCSR[ 167 ][ 338 ],
   alphaCSR[ 167 ][ 339 ],
   alphaCSR[ 167 ][ 340 ],
   alphaCSR[ 167 ][ 341 ],
   alphaCSR[ 167 ][ 342 ],
   alphaCSR[ 167 ][ 343 ],
   alphaCSR[ 167 ][ 344 ],
   alphaCSR[ 167 ][ 345 ],
   alphaCSR[ 167 ][ 346 ],
   alphaCSR[ 167 ][ 347 ],
   alphaCSR[ 167 ][ 348 ],
   alphaCSR[ 167 ][ 349 ],
   alphaCSR[ 167 ][ 350 ],
   alphaCSR[ 167 ][ 351 ],
   alphaCSR[ 167 ][ 352 ],
   alphaCSR[ 167 ][ 353 ],
   alphaCSR[ 167 ][ 354 ],
   alphaCSR[ 167 ][ 355 ],
   alphaCSR[ 167 ][ 356 ],
   alphaCSR[ 167 ][ 357 ],
   alphaCSR[ 167 ][ 358 ],
   alphaCSR[ 167 ][ 359 ],
   alphaCSR[ 167 ][ 360 ],
   alphaCSR[ 167 ][ 361 ],
   alphaCSR[ 167 ][ 362 ],
   alphaCSR[ 167 ][ 363 ],
   alphaCSR[ 167 ][ 364 ],
   alphaCSR[ 167 ][ 365 ],
   alphaCSR[ 167 ][ 366 ],
   alphaCSR[ 167 ][ 367 ],
   alphaCSR[ 167 ][ 368 ],
   alphaCSR[ 167 ][ 369 ],
   alphaCSR[ 167 ][ 370 ],
   alphaCSR[ 167 ][ 371 ],
   alphaCSR[ 167 ][ 372 ],
   alphaCSR[ 167 ][ 373 ],
   alphaCSR[ 167 ][ 374 ],
   alphaCSR[ 167 ][ 375 ],
   alphaCSR[ 167 ][ 376 ],
   alphaCSR[ 167 ][ 377 ],
   alphaCSR[ 167 ][ 378 ],
   alphaCSR[ 167 ][ 379 ],
   alphaCSR[ 167 ][ 380 ],
   alphaCSR[ 167 ][ 381 ],
   alphaCSR[ 167 ][ 382 ],
   alphaCSR[ 167 ][ 383 ],
   alphaCSR[ 168 ][ 0 ],
   alphaCSR[ 168 ][ 1 ],
   alphaCSR[ 168 ][ 2 ],
   alphaCSR[ 168 ][ 3 ],
   alphaCSR[ 168 ][ 4 ],
   alphaCSR[ 168 ][ 5 ],
   alphaCSR[ 168 ][ 6 ],
   alphaCSR[ 168 ][ 7 ],
   alphaCSR[ 168 ][ 8 ],
   alphaCSR[ 168 ][ 9 ],
   alphaCSR[ 168 ][ 10 ],
   alphaCSR[ 168 ][ 11 ],
   alphaCSR[ 168 ][ 12 ],
   alphaCSR[ 168 ][ 13 ],
   alphaCSR[ 168 ][ 14 ],
   alphaCSR[ 168 ][ 15 ],
   alphaCSR[ 168 ][ 16 ],
   alphaCSR[ 168 ][ 17 ],
   alphaCSR[ 168 ][ 18 ],
   alphaCSR[ 168 ][ 19 ],
   alphaCSR[ 168 ][ 20 ],
   alphaCSR[ 168 ][ 21 ],
   alphaCSR[ 168 ][ 22 ],
   alphaCSR[ 168 ][ 23 ],
   alphaCSR[ 168 ][ 24 ],
   alphaCSR[ 168 ][ 25 ],
   alphaCSR[ 168 ][ 26 ],
   alphaCSR[ 168 ][ 27 ],
   alphaCSR[ 168 ][ 28 ],
   alphaCSR[ 168 ][ 29 ],
   alphaCSR[ 168 ][ 30 ],
   alphaCSR[ 168 ][ 31 ],
   alphaCSR[ 168 ][ 32 ],
   alphaCSR[ 168 ][ 33 ],
   alphaCSR[ 168 ][ 34 ],
   alphaCSR[ 168 ][ 35 ],
   alphaCSR[ 168 ][ 36 ],
   alphaCSR[ 168 ][ 37 ],
   alphaCSR[ 168 ][ 38 ],
   alphaCSR[ 168 ][ 39 ],
   alphaCSR[ 168 ][ 40 ],
   alphaCSR[ 168 ][ 41 ],
   alphaCSR[ 168 ][ 42 ],
   alphaCSR[ 168 ][ 43 ],
   alphaCSR[ 168 ][ 44 ],
   alphaCSR[ 168 ][ 45 ],
   alphaCSR[ 168 ][ 46 ],
   alphaCSR[ 168 ][ 47 ],
   alphaCSR[ 168 ][ 48 ],
   alphaCSR[ 168 ][ 49 ],
   alphaCSR[ 168 ][ 50 ],
   alphaCSR[ 168 ][ 51 ],
   alphaCSR[ 168 ][ 52 ],
   alphaCSR[ 168 ][ 53 ],
   alphaCSR[ 168 ][ 54 ],
   alphaCSR[ 168 ][ 55 ],
   alphaCSR[ 168 ][ 56 ],
   alphaCSR[ 168 ][ 57 ],
   alphaCSR[ 168 ][ 58 ],
   alphaCSR[ 168 ][ 59 ],
   alphaCSR[ 168 ][ 60 ],
   alphaCSR[ 168 ][ 61 ],
   alphaCSR[ 168 ][ 62 ],
   alphaCSR[ 168 ][ 63 ],
   alphaCSR[ 168 ][ 64 ],
   alphaCSR[ 168 ][ 65 ],
   alphaCSR[ 168 ][ 66 ],
   alphaCSR[ 168 ][ 67 ],
   alphaCSR[ 168 ][ 68 ],
   alphaCSR[ 168 ][ 69 ],
   alphaCSR[ 168 ][ 70 ],
   alphaCSR[ 168 ][ 71 ],
   alphaCSR[ 168 ][ 72 ],
   alphaCSR[ 168 ][ 73 ],
   alphaCSR[ 168 ][ 74 ],
   alphaCSR[ 168 ][ 75 ],
   alphaCSR[ 168 ][ 76 ],
   alphaCSR[ 168 ][ 77 ],
   alphaCSR[ 168 ][ 78 ],
   alphaCSR[ 168 ][ 79 ],
   alphaCSR[ 168 ][ 80 ],
   alphaCSR[ 168 ][ 81 ],
   alphaCSR[ 168 ][ 82 ],
   alphaCSR[ 168 ][ 83 ],
   alphaCSR[ 168 ][ 84 ],
   alphaCSR[ 168 ][ 85 ],
   alphaCSR[ 168 ][ 86 ],
   alphaCSR[ 168 ][ 87 ],
   alphaCSR[ 168 ][ 88 ],
   alphaCSR[ 168 ][ 89 ],
   alphaCSR[ 168 ][ 90 ],
   alphaCSR[ 168 ][ 91 ],
   alphaCSR[ 168 ][ 92 ],
   alphaCSR[ 168 ][ 93 ],
   alphaCSR[ 168 ][ 94 ],
   alphaCSR[ 168 ][ 95 ],
   alphaCSR[ 168 ][ 96 ],
   alphaCSR[ 168 ][ 97 ],
   alphaCSR[ 168 ][ 98 ],
   alphaCSR[ 168 ][ 99 ],
   alphaCSR[ 168 ][ 100 ],
   alphaCSR[ 168 ][ 101 ],
   alphaCSR[ 168 ][ 102 ],
   alphaCSR[ 168 ][ 103 ],
   alphaCSR[ 168 ][ 104 ],
   alphaCSR[ 168 ][ 105 ],
   alphaCSR[ 168 ][ 106 ],
   alphaCSR[ 168 ][ 107 ],
   alphaCSR[ 168 ][ 108 ],
   alphaCSR[ 168 ][ 109 ],
   alphaCSR[ 168 ][ 110 ],
   alphaCSR[ 168 ][ 111 ],
   alphaCSR[ 168 ][ 112 ],
   alphaCSR[ 168 ][ 113 ],
   alphaCSR[ 168 ][ 114 ],
   alphaCSR[ 168 ][ 115 ],
   alphaCSR[ 168 ][ 116 ],
   alphaCSR[ 168 ][ 117 ],
   alphaCSR[ 168 ][ 118 ],
   alphaCSR[ 168 ][ 119 ],
   alphaCSR[ 168 ][ 120 ],
   alphaCSR[ 168 ][ 121 ],
   alphaCSR[ 168 ][ 122 ],
   alphaCSR[ 168 ][ 123 ],
   alphaCSR[ 168 ][ 124 ],
   alphaCSR[ 168 ][ 125 ],
   alphaCSR[ 168 ][ 126 ],
   alphaCSR[ 168 ][ 127 ],
   alphaCSR[ 168 ][ 128 ],
   alphaCSR[ 168 ][ 129 ],
   alphaCSR[ 168 ][ 130 ],
   alphaCSR[ 168 ][ 131 ],
   alphaCSR[ 168 ][ 132 ],
   alphaCSR[ 168 ][ 133 ],
   alphaCSR[ 168 ][ 134 ],
   alphaCSR[ 168 ][ 135 ],
   alphaCSR[ 168 ][ 136 ],
   alphaCSR[ 168 ][ 137 ],
   alphaCSR[ 168 ][ 138 ],
   alphaCSR[ 168 ][ 139 ],
   alphaCSR[ 168 ][ 140 ],
   alphaCSR[ 168 ][ 141 ],
   alphaCSR[ 168 ][ 142 ],
   alphaCSR[ 168 ][ 143 ],
   alphaCSR[ 168 ][ 144 ],
   alphaCSR[ 168 ][ 145 ],
   alphaCSR[ 168 ][ 146 ],
   alphaCSR[ 168 ][ 147 ],
   alphaCSR[ 168 ][ 148 ],
   alphaCSR[ 168 ][ 149 ],
   alphaCSR[ 168 ][ 150 ],
   alphaCSR[ 168 ][ 151 ],
   alphaCSR[ 168 ][ 152 ],
   alphaCSR[ 168 ][ 153 ],
   alphaCSR[ 168 ][ 154 ],
   alphaCSR[ 168 ][ 155 ],
   alphaCSR[ 168 ][ 156 ],
   alphaCSR[ 168 ][ 157 ],
   alphaCSR[ 168 ][ 158 ],
   alphaCSR[ 168 ][ 159 ],
   alphaCSR[ 168 ][ 160 ],
   alphaCSR[ 168 ][ 161 ],
   alphaCSR[ 168 ][ 162 ],
   alphaCSR[ 168 ][ 163 ],
   alphaCSR[ 168 ][ 164 ],
   alphaCSR[ 168 ][ 165 ],
   alphaCSR[ 168 ][ 166 ],
   alphaCSR[ 168 ][ 167 ],
   alphaCSR[ 168 ][ 168 ],
   alphaCSR[ 168 ][ 169 ],
   alphaCSR[ 168 ][ 170 ],
   alphaCSR[ 168 ][ 171 ],
   alphaCSR[ 168 ][ 172 ],
   alphaCSR[ 168 ][ 173 ],
   alphaCSR[ 168 ][ 174 ],
   alphaCSR[ 168 ][ 175 ],
   alphaCSR[ 168 ][ 176 ],
   alphaCSR[ 168 ][ 177 ],
   alphaCSR[ 168 ][ 178 ],
   alphaCSR[ 168 ][ 179 ],
   alphaCSR[ 168 ][ 180 ],
   alphaCSR[ 168 ][ 181 ],
   alphaCSR[ 168 ][ 182 ],
   alphaCSR[ 168 ][ 183 ],
   alphaCSR[ 168 ][ 184 ],
   alphaCSR[ 168 ][ 185 ],
   alphaCSR[ 168 ][ 186 ],
   alphaCSR[ 168 ][ 187 ],
   alphaCSR[ 168 ][ 188 ],
   alphaCSR[ 168 ][ 189 ],
   alphaCSR[ 168 ][ 190 ],
   alphaCSR[ 168 ][ 191 ],
   alphaCSR[ 168 ][ 192 ],
   alphaCSR[ 168 ][ 193 ],
   alphaCSR[ 168 ][ 194 ],
   alphaCSR[ 168 ][ 195 ],
   alphaCSR[ 168 ][ 196 ],
   alphaCSR[ 168 ][ 197 ],
   alphaCSR[ 168 ][ 198 ],
   alphaCSR[ 168 ][ 199 ],
   alphaCSR[ 168 ][ 200 ],
   alphaCSR[ 168 ][ 201 ],
   alphaCSR[ 168 ][ 202 ],
   alphaCSR[ 168 ][ 203 ],
   alphaCSR[ 168 ][ 204 ],
   alphaCSR[ 168 ][ 205 ],
   alphaCSR[ 168 ][ 206 ],
   alphaCSR[ 168 ][ 207 ],
   alphaCSR[ 168 ][ 208 ],
   alphaCSR[ 168 ][ 209 ],
   alphaCSR[ 168 ][ 210 ],
   alphaCSR[ 168 ][ 211 ],
   alphaCSR[ 168 ][ 212 ],
   alphaCSR[ 168 ][ 213 ],
   alphaCSR[ 168 ][ 214 ],
   alphaCSR[ 168 ][ 215 ],
   alphaCSR[ 168 ][ 216 ],
   alphaCSR[ 168 ][ 217 ],
   alphaCSR[ 168 ][ 218 ],
   alphaCSR[ 168 ][ 219 ],
   alphaCSR[ 168 ][ 220 ],
   alphaCSR[ 168 ][ 221 ],
   alphaCSR[ 168 ][ 222 ],
   alphaCSR[ 168 ][ 223 ],
   alphaCSR[ 168 ][ 224 ],
   alphaCSR[ 168 ][ 225 ],
   alphaCSR[ 168 ][ 226 ],
   alphaCSR[ 168 ][ 227 ],
   alphaCSR[ 168 ][ 228 ],
   alphaCSR[ 168 ][ 229 ],
   alphaCSR[ 168 ][ 230 ],
   alphaCSR[ 168 ][ 231 ],
   alphaCSR[ 168 ][ 232 ],
   alphaCSR[ 168 ][ 233 ],
   alphaCSR[ 168 ][ 234 ],
   alphaCSR[ 168 ][ 235 ],
   alphaCSR[ 168 ][ 236 ],
   alphaCSR[ 168 ][ 237 ],
   alphaCSR[ 168 ][ 238 ],
   alphaCSR[ 168 ][ 239 ],
   alphaCSR[ 168 ][ 240 ],
   alphaCSR[ 168 ][ 241 ],
   alphaCSR[ 168 ][ 242 ],
   alphaCSR[ 168 ][ 243 ],
   alphaCSR[ 168 ][ 244 ],
   alphaCSR[ 168 ][ 245 ],
   alphaCSR[ 168 ][ 246 ],
   alphaCSR[ 168 ][ 247 ],
   alphaCSR[ 168 ][ 248 ],
   alphaCSR[ 168 ][ 249 ],
   alphaCSR[ 168 ][ 250 ],
   alphaCSR[ 168 ][ 251 ],
   alphaCSR[ 168 ][ 252 ],
   alphaCSR[ 168 ][ 253 ],
   alphaCSR[ 168 ][ 254 ],
   alphaCSR[ 168 ][ 255 ],
   alphaCSR[ 168 ][ 256 ],
   alphaCSR[ 168 ][ 257 ],
   alphaCSR[ 168 ][ 258 ],
   alphaCSR[ 168 ][ 259 ],
   alphaCSR[ 168 ][ 260 ],
   alphaCSR[ 168 ][ 261 ],
   alphaCSR[ 168 ][ 262 ],
   alphaCSR[ 168 ][ 263 ],
   alphaCSR[ 168 ][ 264 ],
   alphaCSR[ 168 ][ 265 ],
   alphaCSR[ 168 ][ 266 ],
   alphaCSR[ 168 ][ 267 ],
   alphaCSR[ 168 ][ 268 ],
   alphaCSR[ 168 ][ 269 ],
   alphaCSR[ 168 ][ 270 ],
   alphaCSR[ 168 ][ 271 ],
   alphaCSR[ 168 ][ 272 ],
   alphaCSR[ 168 ][ 273 ],
   alphaCSR[ 168 ][ 274 ],
   alphaCSR[ 168 ][ 275 ],
   alphaCSR[ 168 ][ 276 ],
   alphaCSR[ 168 ][ 277 ],
   alphaCSR[ 168 ][ 278 ],
   alphaCSR[ 168 ][ 279 ],
   alphaCSR[ 168 ][ 280 ],
   alphaCSR[ 168 ][ 281 ],
   alphaCSR[ 168 ][ 282 ],
   alphaCSR[ 168 ][ 283 ],
   alphaCSR[ 168 ][ 284 ],
   alphaCSR[ 168 ][ 285 ],
   alphaCSR[ 168 ][ 286 ],
   alphaCSR[ 168 ][ 287 ],
   alphaCSR[ 168 ][ 288 ],
   alphaCSR[ 168 ][ 289 ],
   alphaCSR[ 168 ][ 290 ],
   alphaCSR[ 168 ][ 291 ],
   alphaCSR[ 168 ][ 292 ],
   alphaCSR[ 168 ][ 293 ],
   alphaCSR[ 168 ][ 294 ],
   alphaCSR[ 168 ][ 295 ],
   alphaCSR[ 168 ][ 296 ],
   alphaCSR[ 168 ][ 297 ],
   alphaCSR[ 168 ][ 298 ],
   alphaCSR[ 168 ][ 299 ],
   alphaCSR[ 168 ][ 300 ],
   alphaCSR[ 168 ][ 301 ],
   alphaCSR[ 168 ][ 302 ],
   alphaCSR[ 168 ][ 303 ],
   alphaCSR[ 168 ][ 304 ],
   alphaCSR[ 168 ][ 305 ],
   alphaCSR[ 168 ][ 306 ],
   alphaCSR[ 168 ][ 307 ],
   alphaCSR[ 168 ][ 308 ],
   alphaCSR[ 168 ][ 309 ],
   alphaCSR[ 168 ][ 310 ],
   alphaCSR[ 168 ][ 311 ],
   alphaCSR[ 168 ][ 312 ],
   alphaCSR[ 168 ][ 313 ],
   alphaCSR[ 168 ][ 314 ],
   alphaCSR[ 168 ][ 315 ],
   alphaCSR[ 168 ][ 316 ],
   alphaCSR[ 168 ][ 317 ],
   alphaCSR[ 168 ][ 318 ],
   alphaCSR[ 168 ][ 319 ],
   alphaCSR[ 168 ][ 320 ],
   alphaCSR[ 168 ][ 321 ],
   alphaCSR[ 168 ][ 322 ],
   alphaCSR[ 168 ][ 323 ],
   alphaCSR[ 168 ][ 324 ],
   alphaCSR[ 168 ][ 325 ],
   alphaCSR[ 168 ][ 326 ],
   alphaCSR[ 168 ][ 327 ],
   alphaCSR[ 168 ][ 328 ],
   alphaCSR[ 168 ][ 329 ],
   alphaCSR[ 168 ][ 330 ],
   alphaCSR[ 168 ][ 331 ],
   alphaCSR[ 168 ][ 332 ],
   alphaCSR[ 168 ][ 333 ],
   alphaCSR[ 168 ][ 334 ],
   alphaCSR[ 168 ][ 335 ],
   alphaCSR[ 168 ][ 336 ],
   alphaCSR[ 168 ][ 337 ],
   alphaCSR[ 168 ][ 338 ],
   alphaCSR[ 168 ][ 339 ],
   alphaCSR[ 168 ][ 340 ],
   alphaCSR[ 168 ][ 341 ],
   alphaCSR[ 168 ][ 342 ],
   alphaCSR[ 168 ][ 343 ],
   alphaCSR[ 168 ][ 344 ],
   alphaCSR[ 168 ][ 345 ],
   alphaCSR[ 168 ][ 346 ],
   alphaCSR[ 168 ][ 347 ],
   alphaCSR[ 168 ][ 348 ],
   alphaCSR[ 168 ][ 349 ],
   alphaCSR[ 168 ][ 350 ],
   alphaCSR[ 168 ][ 351 ],
   alphaCSR[ 168 ][ 352 ],
   alphaCSR[ 168 ][ 353 ],
   alphaCSR[ 168 ][ 354 ],
   alphaCSR[ 168 ][ 355 ],
   alphaCSR[ 168 ][ 356 ],
   alphaCSR[ 168 ][ 357 ],
   alphaCSR[ 168 ][ 358 ],
   alphaCSR[ 168 ][ 359 ],
   alphaCSR[ 168 ][ 360 ],
   alphaCSR[ 168 ][ 361 ],
   alphaCSR[ 168 ][ 362 ],
   alphaCSR[ 168 ][ 363 ],
   alphaCSR[ 168 ][ 364 ],
   alphaCSR[ 168 ][ 365 ],
   alphaCSR[ 168 ][ 366 ],
   alphaCSR[ 168 ][ 367 ],
   alphaCSR[ 168 ][ 368 ],
   alphaCSR[ 168 ][ 369 ],
   alphaCSR[ 168 ][ 370 ],
   alphaCSR[ 168 ][ 371 ],
   alphaCSR[ 168 ][ 372 ],
   alphaCSR[ 168 ][ 373 ],
   alphaCSR[ 168 ][ 374 ],
   alphaCSR[ 168 ][ 375 ],
   alphaCSR[ 168 ][ 376 ],
   alphaCSR[ 168 ][ 377 ],
   alphaCSR[ 168 ][ 378 ],
   alphaCSR[ 168 ][ 379 ],
   alphaCSR[ 168 ][ 380 ],
   alphaCSR[ 168 ][ 381 ],
   alphaCSR[ 168 ][ 382 ],
   alphaCSR[ 168 ][ 383 ],
   alphaCSR[ 169 ][ 0 ],
   alphaCSR[ 169 ][ 1 ],
   alphaCSR[ 169 ][ 2 ],
   alphaCSR[ 169 ][ 3 ],
   alphaCSR[ 169 ][ 4 ],
   alphaCSR[ 169 ][ 5 ],
   alphaCSR[ 169 ][ 6 ],
   alphaCSR[ 169 ][ 7 ],
   alphaCSR[ 169 ][ 8 ],
   alphaCSR[ 169 ][ 9 ],
   alphaCSR[ 169 ][ 10 ],
   alphaCSR[ 169 ][ 11 ],
   alphaCSR[ 169 ][ 12 ],
   alphaCSR[ 169 ][ 13 ],
   alphaCSR[ 169 ][ 14 ],
   alphaCSR[ 169 ][ 15 ],
   alphaCSR[ 169 ][ 16 ],
   alphaCSR[ 169 ][ 17 ],
   alphaCSR[ 169 ][ 18 ],
   alphaCSR[ 169 ][ 19 ],
   alphaCSR[ 169 ][ 20 ],
   alphaCSR[ 169 ][ 21 ],
   alphaCSR[ 169 ][ 22 ],
   alphaCSR[ 169 ][ 23 ],
   alphaCSR[ 169 ][ 24 ],
   alphaCSR[ 169 ][ 25 ],
   alphaCSR[ 169 ][ 26 ],
   alphaCSR[ 169 ][ 27 ],
   alphaCSR[ 169 ][ 28 ],
   alphaCSR[ 169 ][ 29 ],
   alphaCSR[ 169 ][ 30 ],
   alphaCSR[ 169 ][ 31 ],
   alphaCSR[ 169 ][ 32 ],
   alphaCSR[ 169 ][ 33 ],
   alphaCSR[ 169 ][ 34 ],
   alphaCSR[ 169 ][ 35 ],
   alphaCSR[ 169 ][ 36 ],
   alphaCSR[ 169 ][ 37 ],
   alphaCSR[ 169 ][ 38 ],
   alphaCSR[ 169 ][ 39 ],
   alphaCSR[ 169 ][ 40 ],
   alphaCSR[ 169 ][ 41 ],
   alphaCSR[ 169 ][ 42 ],
   alphaCSR[ 169 ][ 43 ],
   alphaCSR[ 169 ][ 44 ],
   alphaCSR[ 169 ][ 45 ],
   alphaCSR[ 169 ][ 46 ],
   alphaCSR[ 169 ][ 47 ],
   alphaCSR[ 169 ][ 48 ],
   alphaCSR[ 169 ][ 49 ],
   alphaCSR[ 169 ][ 50 ],
   alphaCSR[ 169 ][ 51 ],
   alphaCSR[ 169 ][ 52 ],
   alphaCSR[ 169 ][ 53 ],
   alphaCSR[ 169 ][ 54 ],
   alphaCSR[ 169 ][ 55 ],
   alphaCSR[ 169 ][ 56 ],
   alphaCSR[ 169 ][ 57 ],
   alphaCSR[ 169 ][ 58 ],
   alphaCSR[ 169 ][ 59 ],
   alphaCSR[ 169 ][ 60 ],
   alphaCSR[ 169 ][ 61 ],
   alphaCSR[ 169 ][ 62 ],
   alphaCSR[ 169 ][ 63 ],
   alphaCSR[ 169 ][ 64 ],
   alphaCSR[ 169 ][ 65 ],
   alphaCSR[ 169 ][ 66 ],
   alphaCSR[ 169 ][ 67 ],
   alphaCSR[ 169 ][ 68 ],
   alphaCSR[ 169 ][ 69 ],
   alphaCSR[ 169 ][ 70 ],
   alphaCSR[ 169 ][ 71 ],
   alphaCSR[ 169 ][ 72 ],
   alphaCSR[ 169 ][ 73 ],
   alphaCSR[ 169 ][ 74 ],
   alphaCSR[ 169 ][ 75 ],
   alphaCSR[ 169 ][ 76 ],
   alphaCSR[ 169 ][ 77 ],
   alphaCSR[ 169 ][ 78 ],
   alphaCSR[ 169 ][ 79 ],
   alphaCSR[ 169 ][ 80 ],
   alphaCSR[ 169 ][ 81 ],
   alphaCSR[ 169 ][ 82 ],
   alphaCSR[ 169 ][ 83 ],
   alphaCSR[ 169 ][ 84 ],
   alphaCSR[ 169 ][ 85 ],
   alphaCSR[ 169 ][ 86 ],
   alphaCSR[ 169 ][ 87 ],
   alphaCSR[ 169 ][ 88 ],
   alphaCSR[ 169 ][ 89 ],
   alphaCSR[ 169 ][ 90 ],
   alphaCSR[ 169 ][ 91 ],
   alphaCSR[ 169 ][ 92 ],
   alphaCSR[ 169 ][ 93 ],
   alphaCSR[ 169 ][ 94 ],
   alphaCSR[ 169 ][ 95 ],
   alphaCSR[ 169 ][ 96 ],
   alphaCSR[ 169 ][ 97 ],
   alphaCSR[ 169 ][ 98 ],
   alphaCSR[ 169 ][ 99 ],
   alphaCSR[ 169 ][ 100 ],
   alphaCSR[ 169 ][ 101 ],
   alphaCSR[ 169 ][ 102 ],
   alphaCSR[ 169 ][ 103 ],
   alphaCSR[ 169 ][ 104 ],
   alphaCSR[ 169 ][ 105 ],
   alphaCSR[ 169 ][ 106 ],
   alphaCSR[ 169 ][ 107 ],
   alphaCSR[ 169 ][ 108 ],
   alphaCSR[ 169 ][ 109 ],
   alphaCSR[ 169 ][ 110 ],
   alphaCSR[ 169 ][ 111 ],
   alphaCSR[ 169 ][ 112 ],
   alphaCSR[ 169 ][ 113 ],
   alphaCSR[ 169 ][ 114 ],
   alphaCSR[ 169 ][ 115 ],
   alphaCSR[ 169 ][ 116 ],
   alphaCSR[ 169 ][ 117 ],
   alphaCSR[ 169 ][ 118 ],
   alphaCSR[ 169 ][ 119 ],
   alphaCSR[ 169 ][ 120 ],
   alphaCSR[ 169 ][ 121 ],
   alphaCSR[ 169 ][ 122 ],
   alphaCSR[ 169 ][ 123 ],
   alphaCSR[ 169 ][ 124 ],
   alphaCSR[ 169 ][ 125 ],
   alphaCSR[ 169 ][ 126 ],
   alphaCSR[ 169 ][ 127 ],
   alphaCSR[ 169 ][ 128 ],
   alphaCSR[ 169 ][ 129 ],
   alphaCSR[ 169 ][ 130 ],
   alphaCSR[ 169 ][ 131 ],
   alphaCSR[ 169 ][ 132 ],
   alphaCSR[ 169 ][ 133 ],
   alphaCSR[ 169 ][ 134 ],
   alphaCSR[ 169 ][ 135 ],
   alphaCSR[ 169 ][ 136 ],
   alphaCSR[ 169 ][ 137 ],
   alphaCSR[ 169 ][ 138 ],
   alphaCSR[ 169 ][ 139 ],
   alphaCSR[ 169 ][ 140 ],
   alphaCSR[ 169 ][ 141 ],
   alphaCSR[ 169 ][ 142 ],
   alphaCSR[ 169 ][ 143 ],
   alphaCSR[ 169 ][ 144 ],
   alphaCSR[ 169 ][ 145 ],
   alphaCSR[ 169 ][ 146 ],
   alphaCSR[ 169 ][ 147 ],
   alphaCSR[ 169 ][ 148 ],
   alphaCSR[ 169 ][ 149 ],
   alphaCSR[ 169 ][ 150 ],
   alphaCSR[ 169 ][ 151 ],
   alphaCSR[ 169 ][ 152 ],
   alphaCSR[ 169 ][ 153 ],
   alphaCSR[ 169 ][ 154 ],
   alphaCSR[ 169 ][ 155 ],
   alphaCSR[ 169 ][ 156 ],
   alphaCSR[ 169 ][ 157 ],
   alphaCSR[ 169 ][ 158 ],
   alphaCSR[ 169 ][ 159 ],
   alphaCSR[ 169 ][ 160 ],
   alphaCSR[ 169 ][ 161 ],
   alphaCSR[ 169 ][ 162 ],
   alphaCSR[ 169 ][ 163 ],
   alphaCSR[ 169 ][ 164 ],
   alphaCSR[ 169 ][ 165 ],
   alphaCSR[ 169 ][ 166 ],
   alphaCSR[ 169 ][ 167 ],
   alphaCSR[ 169 ][ 168 ],
   alphaCSR[ 169 ][ 169 ],
   alphaCSR[ 169 ][ 170 ],
   alphaCSR[ 169 ][ 171 ],
   alphaCSR[ 169 ][ 172 ],
   alphaCSR[ 169 ][ 173 ],
   alphaCSR[ 169 ][ 174 ],
   alphaCSR[ 169 ][ 175 ],
   alphaCSR[ 169 ][ 176 ],
   alphaCSR[ 169 ][ 177 ],
   alphaCSR[ 169 ][ 178 ],
   alphaCSR[ 169 ][ 179 ],
   alphaCSR[ 169 ][ 180 ],
   alphaCSR[ 169 ][ 181 ],
   alphaCSR[ 169 ][ 182 ],
   alphaCSR[ 169 ][ 183 ],
   alphaCSR[ 169 ][ 184 ],
   alphaCSR[ 169 ][ 185 ],
   alphaCSR[ 169 ][ 186 ],
   alphaCSR[ 169 ][ 187 ],
   alphaCSR[ 169 ][ 188 ],
   alphaCSR[ 169 ][ 189 ],
   alphaCSR[ 169 ][ 190 ],
   alphaCSR[ 169 ][ 191 ],
   alphaCSR[ 169 ][ 192 ],
   alphaCSR[ 169 ][ 193 ],
   alphaCSR[ 169 ][ 194 ],
   alphaCSR[ 169 ][ 195 ],
   alphaCSR[ 169 ][ 196 ],
   alphaCSR[ 169 ][ 197 ],
   alphaCSR[ 169 ][ 198 ],
   alphaCSR[ 169 ][ 199 ],
   alphaCSR[ 169 ][ 200 ],
   alphaCSR[ 169 ][ 201 ],
   alphaCSR[ 169 ][ 202 ],
   alphaCSR[ 169 ][ 203 ],
   alphaCSR[ 169 ][ 204 ],
   alphaCSR[ 169 ][ 205 ],
   alphaCSR[ 169 ][ 206 ],
   alphaCSR[ 169 ][ 207 ],
   alphaCSR[ 169 ][ 208 ],
   alphaCSR[ 169 ][ 209 ],
   alphaCSR[ 169 ][ 210 ],
   alphaCSR[ 169 ][ 211 ],
   alphaCSR[ 169 ][ 212 ],
   alphaCSR[ 169 ][ 213 ],
   alphaCSR[ 169 ][ 214 ],
   alphaCSR[ 169 ][ 215 ],
   alphaCSR[ 169 ][ 216 ],
   alphaCSR[ 169 ][ 217 ],
   alphaCSR[ 169 ][ 218 ],
   alphaCSR[ 169 ][ 219 ],
   alphaCSR[ 169 ][ 220 ],
   alphaCSR[ 169 ][ 221 ],
   alphaCSR[ 169 ][ 222 ],
   alphaCSR[ 169 ][ 223 ],
   alphaCSR[ 169 ][ 224 ],
   alphaCSR[ 169 ][ 225 ],
   alphaCSR[ 169 ][ 226 ],
   alphaCSR[ 169 ][ 227 ],
   alphaCSR[ 169 ][ 228 ],
   alphaCSR[ 169 ][ 229 ],
   alphaCSR[ 169 ][ 230 ],
   alphaCSR[ 169 ][ 231 ],
   alphaCSR[ 169 ][ 232 ],
   alphaCSR[ 169 ][ 233 ],
   alphaCSR[ 169 ][ 234 ],
   alphaCSR[ 169 ][ 235 ],
   alphaCSR[ 169 ][ 236 ],
   alphaCSR[ 169 ][ 237 ],
   alphaCSR[ 169 ][ 238 ],
   alphaCSR[ 169 ][ 239 ],
   alphaCSR[ 169 ][ 240 ],
   alphaCSR[ 169 ][ 241 ],
   alphaCSR[ 169 ][ 242 ],
   alphaCSR[ 169 ][ 243 ],
   alphaCSR[ 169 ][ 244 ],
   alphaCSR[ 169 ][ 245 ],
   alphaCSR[ 169 ][ 246 ],
   alphaCSR[ 169 ][ 247 ],
   alphaCSR[ 169 ][ 248 ],
   alphaCSR[ 169 ][ 249 ],
   alphaCSR[ 169 ][ 250 ],
   alphaCSR[ 169 ][ 251 ],
   alphaCSR[ 169 ][ 252 ],
   alphaCSR[ 169 ][ 253 ],
   alphaCSR[ 169 ][ 254 ],
   alphaCSR[ 169 ][ 255 ],
   alphaCSR[ 169 ][ 256 ],
   alphaCSR[ 169 ][ 257 ],
   alphaCSR[ 169 ][ 258 ],
   alphaCSR[ 169 ][ 259 ],
   alphaCSR[ 169 ][ 260 ],
   alphaCSR[ 169 ][ 261 ],
   alphaCSR[ 169 ][ 262 ],
   alphaCSR[ 169 ][ 263 ],
   alphaCSR[ 169 ][ 264 ],
   alphaCSR[ 169 ][ 265 ],
   alphaCSR[ 169 ][ 266 ],
   alphaCSR[ 169 ][ 267 ],
   alphaCSR[ 169 ][ 268 ],
   alphaCSR[ 169 ][ 269 ],
   alphaCSR[ 169 ][ 270 ],
   alphaCSR[ 169 ][ 271 ],
   alphaCSR[ 169 ][ 272 ],
   alphaCSR[ 169 ][ 273 ],
   alphaCSR[ 169 ][ 274 ],
   alphaCSR[ 169 ][ 275 ],
   alphaCSR[ 169 ][ 276 ],
   alphaCSR[ 169 ][ 277 ],
   alphaCSR[ 169 ][ 278 ],
   alphaCSR[ 169 ][ 279 ],
   alphaCSR[ 169 ][ 280 ],
   alphaCSR[ 169 ][ 281 ],
   alphaCSR[ 169 ][ 282 ],
   alphaCSR[ 169 ][ 283 ],
   alphaCSR[ 169 ][ 284 ],
   alphaCSR[ 169 ][ 285 ],
   alphaCSR[ 169 ][ 286 ],
   alphaCSR[ 169 ][ 287 ],
   alphaCSR[ 169 ][ 288 ],
   alphaCSR[ 169 ][ 289 ],
   alphaCSR[ 169 ][ 290 ],
   alphaCSR[ 169 ][ 291 ],
   alphaCSR[ 169 ][ 292 ],
   alphaCSR[ 169 ][ 293 ],
   alphaCSR[ 169 ][ 294 ],
   alphaCSR[ 169 ][ 295 ],
   alphaCSR[ 169 ][ 296 ],
   alphaCSR[ 169 ][ 297 ],
   alphaCSR[ 169 ][ 298 ],
   alphaCSR[ 169 ][ 299 ],
   alphaCSR[ 169 ][ 300 ],
   alphaCSR[ 169 ][ 301 ],
   alphaCSR[ 169 ][ 302 ],
   alphaCSR[ 169 ][ 303 ],
   alphaCSR[ 169 ][ 304 ],
   alphaCSR[ 169 ][ 305 ],
   alphaCSR[ 169 ][ 306 ],
   alphaCSR[ 169 ][ 307 ],
   alphaCSR[ 169 ][ 308 ],
   alphaCSR[ 169 ][ 309 ],
   alphaCSR[ 169 ][ 310 ],
   alphaCSR[ 169 ][ 311 ],
   alphaCSR[ 169 ][ 312 ],
   alphaCSR[ 169 ][ 313 ],
   alphaCSR[ 169 ][ 314 ],
   alphaCSR[ 169 ][ 315 ],
   alphaCSR[ 169 ][ 316 ],
   alphaCSR[ 169 ][ 317 ],
   alphaCSR[ 169 ][ 318 ],
   alphaCSR[ 169 ][ 319 ],
   alphaCSR[ 169 ][ 320 ],
   alphaCSR[ 169 ][ 321 ],
   alphaCSR[ 169 ][ 322 ],
   alphaCSR[ 169 ][ 323 ],
   alphaCSR[ 169 ][ 324 ],
   alphaCSR[ 169 ][ 325 ],
   alphaCSR[ 169 ][ 326 ],
   alphaCSR[ 169 ][ 327 ],
   alphaCSR[ 169 ][ 328 ],
   alphaCSR[ 169 ][ 329 ],
   alphaCSR[ 169 ][ 330 ],
   alphaCSR[ 169 ][ 331 ],
   alphaCSR[ 169 ][ 332 ],
   alphaCSR[ 169 ][ 333 ],
   alphaCSR[ 169 ][ 334 ],
   alphaCSR[ 169 ][ 335 ],
   alphaCSR[ 169 ][ 336 ],
   alphaCSR[ 169 ][ 337 ],
   alphaCSR[ 169 ][ 338 ],
   alphaCSR[ 169 ][ 339 ],
   alphaCSR[ 169 ][ 340 ],
   alphaCSR[ 169 ][ 341 ],
   alphaCSR[ 169 ][ 342 ],
   alphaCSR[ 169 ][ 343 ],
   alphaCSR[ 169 ][ 344 ],
   alphaCSR[ 169 ][ 345 ],
   alphaCSR[ 169 ][ 346 ],
   alphaCSR[ 169 ][ 347 ],
   alphaCSR[ 169 ][ 348 ],
   alphaCSR[ 169 ][ 349 ],
   alphaCSR[ 169 ][ 350 ],
   alphaCSR[ 169 ][ 351 ],
   alphaCSR[ 169 ][ 352 ],
   alphaCSR[ 169 ][ 353 ],
   alphaCSR[ 169 ][ 354 ],
   alphaCSR[ 169 ][ 355 ],
   alphaCSR[ 169 ][ 356 ],
   alphaCSR[ 169 ][ 357 ],
   alphaCSR[ 169 ][ 358 ],
   alphaCSR[ 169 ][ 359 ],
   alphaCSR[ 169 ][ 360 ],
   alphaCSR[ 169 ][ 361 ],
   alphaCSR[ 169 ][ 362 ],
   alphaCSR[ 169 ][ 363 ],
   alphaCSR[ 169 ][ 364 ],
   alphaCSR[ 169 ][ 365 ],
   alphaCSR[ 169 ][ 366 ],
   alphaCSR[ 169 ][ 367 ],
   alphaCSR[ 169 ][ 368 ],
   alphaCSR[ 169 ][ 369 ],
   alphaCSR[ 169 ][ 370 ],
   alphaCSR[ 169 ][ 371 ],
   alphaCSR[ 169 ][ 372 ],
   alphaCSR[ 169 ][ 373 ],
   alphaCSR[ 169 ][ 374 ],
   alphaCSR[ 169 ][ 375 ],
   alphaCSR[ 169 ][ 376 ],
   alphaCSR[ 169 ][ 377 ],
   alphaCSR[ 169 ][ 378 ],
   alphaCSR[ 169 ][ 379 ],
   alphaCSR[ 169 ][ 380 ],
   alphaCSR[ 169 ][ 381 ],
   alphaCSR[ 169 ][ 382 ],
   alphaCSR[ 169 ][ 383 ],
   alphaCSR[ 170 ][ 0 ],
   alphaCSR[ 170 ][ 1 ],
   alphaCSR[ 170 ][ 2 ],
   alphaCSR[ 170 ][ 3 ],
   alphaCSR[ 170 ][ 4 ],
   alphaCSR[ 170 ][ 5 ],
   alphaCSR[ 170 ][ 6 ],
   alphaCSR[ 170 ][ 7 ],
   alphaCSR[ 170 ][ 8 ],
   alphaCSR[ 170 ][ 9 ],
   alphaCSR[ 170 ][ 10 ],
   alphaCSR[ 170 ][ 11 ],
   alphaCSR[ 170 ][ 12 ],
   alphaCSR[ 170 ][ 13 ],
   alphaCSR[ 170 ][ 14 ],
   alphaCSR[ 170 ][ 15 ],
   alphaCSR[ 170 ][ 16 ],
   alphaCSR[ 170 ][ 17 ],
   alphaCSR[ 170 ][ 18 ],
   alphaCSR[ 170 ][ 19 ],
   alphaCSR[ 170 ][ 20 ],
   alphaCSR[ 170 ][ 21 ],
   alphaCSR[ 170 ][ 22 ],
   alphaCSR[ 170 ][ 23 ],
   alphaCSR[ 170 ][ 24 ],
   alphaCSR[ 170 ][ 25 ],
   alphaCSR[ 170 ][ 26 ],
   alphaCSR[ 170 ][ 27 ],
   alphaCSR[ 170 ][ 28 ],
   alphaCSR[ 170 ][ 29 ],
   alphaCSR[ 170 ][ 30 ],
   alphaCSR[ 170 ][ 31 ],
   alphaCSR[ 170 ][ 32 ],
   alphaCSR[ 170 ][ 33 ],
   alphaCSR[ 170 ][ 34 ],
   alphaCSR[ 170 ][ 35 ],
   alphaCSR[ 170 ][ 36 ],
   alphaCSR[ 170 ][ 37 ],
   alphaCSR[ 170 ][ 38 ],
   alphaCSR[ 170 ][ 39 ],
   alphaCSR[ 170 ][ 40 ],
   alphaCSR[ 170 ][ 41 ],
   alphaCSR[ 170 ][ 42 ],
   alphaCSR[ 170 ][ 43 ],
   alphaCSR[ 170 ][ 44 ],
   alphaCSR[ 170 ][ 45 ],
   alphaCSR[ 170 ][ 46 ],
   alphaCSR[ 170 ][ 47 ],
   alphaCSR[ 170 ][ 48 ],
   alphaCSR[ 170 ][ 49 ],
   alphaCSR[ 170 ][ 50 ],
   alphaCSR[ 170 ][ 51 ],
   alphaCSR[ 170 ][ 52 ],
   alphaCSR[ 170 ][ 53 ],
   alphaCSR[ 170 ][ 54 ],
   alphaCSR[ 170 ][ 55 ],
   alphaCSR[ 170 ][ 56 ],
   alphaCSR[ 170 ][ 57 ],
   alphaCSR[ 170 ][ 58 ],
   alphaCSR[ 170 ][ 59 ],
   alphaCSR[ 170 ][ 60 ],
   alphaCSR[ 170 ][ 61 ],
   alphaCSR[ 170 ][ 62 ],
   alphaCSR[ 170 ][ 63 ],
   alphaCSR[ 170 ][ 64 ],
   alphaCSR[ 170 ][ 65 ],
   alphaCSR[ 170 ][ 66 ],
   alphaCSR[ 170 ][ 67 ],
   alphaCSR[ 170 ][ 68 ],
   alphaCSR[ 170 ][ 69 ],
   alphaCSR[ 170 ][ 70 ],
   alphaCSR[ 170 ][ 71 ],
   alphaCSR[ 170 ][ 72 ],
   alphaCSR[ 170 ][ 73 ],
   alphaCSR[ 170 ][ 74 ],
   alphaCSR[ 170 ][ 75 ],
   alphaCSR[ 170 ][ 76 ],
   alphaCSR[ 170 ][ 77 ],
   alphaCSR[ 170 ][ 78 ],
   alphaCSR[ 170 ][ 79 ],
   alphaCSR[ 170 ][ 80 ],
   alphaCSR[ 170 ][ 81 ],
   alphaCSR[ 170 ][ 82 ],
   alphaCSR[ 170 ][ 83 ],
   alphaCSR[ 170 ][ 84 ],
   alphaCSR[ 170 ][ 85 ],
   alphaCSR[ 170 ][ 86 ],
   alphaCSR[ 170 ][ 87 ],
   alphaCSR[ 170 ][ 88 ],
   alphaCSR[ 170 ][ 89 ],
   alphaCSR[ 170 ][ 90 ],
   alphaCSR[ 170 ][ 91 ],
   alphaCSR[ 170 ][ 92 ],
   alphaCSR[ 170 ][ 93 ],
   alphaCSR[ 170 ][ 94 ],
   alphaCSR[ 170 ][ 95 ],
   alphaCSR[ 170 ][ 96 ],
   alphaCSR[ 170 ][ 97 ],
   alphaCSR[ 170 ][ 98 ],
   alphaCSR[ 170 ][ 99 ],
   alphaCSR[ 170 ][ 100 ],
   alphaCSR[ 170 ][ 101 ],
   alphaCSR[ 170 ][ 102 ],
   alphaCSR[ 170 ][ 103 ],
   alphaCSR[ 170 ][ 104 ],
   alphaCSR[ 170 ][ 105 ],
   alphaCSR[ 170 ][ 106 ],
   alphaCSR[ 170 ][ 107 ],
   alphaCSR[ 170 ][ 108 ],
   alphaCSR[ 170 ][ 109 ],
   alphaCSR[ 170 ][ 110 ],
   alphaCSR[ 170 ][ 111 ],
   alphaCSR[ 170 ][ 112 ],
   alphaCSR[ 170 ][ 113 ],
   alphaCSR[ 170 ][ 114 ],
   alphaCSR[ 170 ][ 115 ],
   alphaCSR[ 170 ][ 116 ],
   alphaCSR[ 170 ][ 117 ],
   alphaCSR[ 170 ][ 118 ],
   alphaCSR[ 170 ][ 119 ],
   alphaCSR[ 170 ][ 120 ],
   alphaCSR[ 170 ][ 121 ],
   alphaCSR[ 170 ][ 122 ],
   alphaCSR[ 170 ][ 123 ],
   alphaCSR[ 170 ][ 124 ],
   alphaCSR[ 170 ][ 125 ],
   alphaCSR[ 170 ][ 126 ],
   alphaCSR[ 170 ][ 127 ],
   alphaCSR[ 170 ][ 128 ],
   alphaCSR[ 170 ][ 129 ],
   alphaCSR[ 170 ][ 130 ],
   alphaCSR[ 170 ][ 131 ],
   alphaCSR[ 170 ][ 132 ],
   alphaCSR[ 170 ][ 133 ],
   alphaCSR[ 170 ][ 134 ],
   alphaCSR[ 170 ][ 135 ],
   alphaCSR[ 170 ][ 136 ],
   alphaCSR[ 170 ][ 137 ],
   alphaCSR[ 170 ][ 138 ],
   alphaCSR[ 170 ][ 139 ],
   alphaCSR[ 170 ][ 140 ],
   alphaCSR[ 170 ][ 141 ],
   alphaCSR[ 170 ][ 142 ],
   alphaCSR[ 170 ][ 143 ],
   alphaCSR[ 170 ][ 144 ],
   alphaCSR[ 170 ][ 145 ],
   alphaCSR[ 170 ][ 146 ],
   alphaCSR[ 170 ][ 147 ],
   alphaCSR[ 170 ][ 148 ],
   alphaCSR[ 170 ][ 149 ],
   alphaCSR[ 170 ][ 150 ],
   alphaCSR[ 170 ][ 151 ],
   alphaCSR[ 170 ][ 152 ],
   alphaCSR[ 170 ][ 153 ],
   alphaCSR[ 170 ][ 154 ],
   alphaCSR[ 170 ][ 155 ],
   alphaCSR[ 170 ][ 156 ],
   alphaCSR[ 170 ][ 157 ],
   alphaCSR[ 170 ][ 158 ],
   alphaCSR[ 170 ][ 159 ],
   alphaCSR[ 170 ][ 160 ],
   alphaCSR[ 170 ][ 161 ],
   alphaCSR[ 170 ][ 162 ],
   alphaCSR[ 170 ][ 163 ],
   alphaCSR[ 170 ][ 164 ],
   alphaCSR[ 170 ][ 165 ],
   alphaCSR[ 170 ][ 166 ],
   alphaCSR[ 170 ][ 167 ],
   alphaCSR[ 170 ][ 168 ],
   alphaCSR[ 170 ][ 169 ],
   alphaCSR[ 170 ][ 170 ],
   alphaCSR[ 170 ][ 171 ],
   alphaCSR[ 170 ][ 172 ],
   alphaCSR[ 170 ][ 173 ],
   alphaCSR[ 170 ][ 174 ],
   alphaCSR[ 170 ][ 175 ],
   alphaCSR[ 170 ][ 176 ],
   alphaCSR[ 170 ][ 177 ],
   alphaCSR[ 170 ][ 178 ],
   alphaCSR[ 170 ][ 179 ],
   alphaCSR[ 170 ][ 180 ],
   alphaCSR[ 170 ][ 181 ],
   alphaCSR[ 170 ][ 182 ],
   alphaCSR[ 170 ][ 183 ],
   alphaCSR[ 170 ][ 184 ],
   alphaCSR[ 170 ][ 185 ],
   alphaCSR[ 170 ][ 186 ],
   alphaCSR[ 170 ][ 187 ],
   alphaCSR[ 170 ][ 188 ],
   alphaCSR[ 170 ][ 189 ],
   alphaCSR[ 170 ][ 190 ],
   alphaCSR[ 170 ][ 191 ],
   alphaCSR[ 170 ][ 192 ],
   alphaCSR[ 170 ][ 193 ],
   alphaCSR[ 170 ][ 194 ],
   alphaCSR[ 170 ][ 195 ],
   alphaCSR[ 170 ][ 196 ],
   alphaCSR[ 170 ][ 197 ],
   alphaCSR[ 170 ][ 198 ],
   alphaCSR[ 170 ][ 199 ],
   alphaCSR[ 170 ][ 200 ],
   alphaCSR[ 170 ][ 201 ],
   alphaCSR[ 170 ][ 202 ],
   alphaCSR[ 170 ][ 203 ],
   alphaCSR[ 170 ][ 204 ],
   alphaCSR[ 170 ][ 205 ],
   alphaCSR[ 170 ][ 206 ],
   alphaCSR[ 170 ][ 207 ],
   alphaCSR[ 170 ][ 208 ],
   alphaCSR[ 170 ][ 209 ],
   alphaCSR[ 170 ][ 210 ],
   alphaCSR[ 170 ][ 211 ],
   alphaCSR[ 170 ][ 212 ],
   alphaCSR[ 170 ][ 213 ],
   alphaCSR[ 170 ][ 214 ],
   alphaCSR[ 170 ][ 215 ],
   alphaCSR[ 170 ][ 216 ],
   alphaCSR[ 170 ][ 217 ],
   alphaCSR[ 170 ][ 218 ],
   alphaCSR[ 170 ][ 219 ],
   alphaCSR[ 170 ][ 220 ],
   alphaCSR[ 170 ][ 221 ],
   alphaCSR[ 170 ][ 222 ],
   alphaCSR[ 170 ][ 223 ],
   alphaCSR[ 170 ][ 224 ],
   alphaCSR[ 170 ][ 225 ],
   alphaCSR[ 170 ][ 226 ],
   alphaCSR[ 170 ][ 227 ],
   alphaCSR[ 170 ][ 228 ],
   alphaCSR[ 170 ][ 229 ],
   alphaCSR[ 170 ][ 230 ],
   alphaCSR[ 170 ][ 231 ],
   alphaCSR[ 170 ][ 232 ],
   alphaCSR[ 170 ][ 233 ],
   alphaCSR[ 170 ][ 234 ],
   alphaCSR[ 170 ][ 235 ],
   alphaCSR[ 170 ][ 236 ],
   alphaCSR[ 170 ][ 237 ],
   alphaCSR[ 170 ][ 238 ],
   alphaCSR[ 170 ][ 239 ],
   alphaCSR[ 170 ][ 240 ],
   alphaCSR[ 170 ][ 241 ],
   alphaCSR[ 170 ][ 242 ],
   alphaCSR[ 170 ][ 243 ],
   alphaCSR[ 170 ][ 244 ],
   alphaCSR[ 170 ][ 245 ],
   alphaCSR[ 170 ][ 246 ],
   alphaCSR[ 170 ][ 247 ],
   alphaCSR[ 170 ][ 248 ],
   alphaCSR[ 170 ][ 249 ],
   alphaCSR[ 170 ][ 250 ],
   alphaCSR[ 170 ][ 251 ],
   alphaCSR[ 170 ][ 252 ],
   alphaCSR[ 170 ][ 253 ],
   alphaCSR[ 170 ][ 254 ],
   alphaCSR[ 170 ][ 255 ],
   alphaCSR[ 170 ][ 256 ],
   alphaCSR[ 170 ][ 257 ],
   alphaCSR[ 170 ][ 258 ],
   alphaCSR[ 170 ][ 259 ],
   alphaCSR[ 170 ][ 260 ],
   alphaCSR[ 170 ][ 261 ],
   alphaCSR[ 170 ][ 262 ],
   alphaCSR[ 170 ][ 263 ],
   alphaCSR[ 170 ][ 264 ],
   alphaCSR[ 170 ][ 265 ],
   alphaCSR[ 170 ][ 266 ],
   alphaCSR[ 170 ][ 267 ],
   alphaCSR[ 170 ][ 268 ],
   alphaCSR[ 170 ][ 269 ],
   alphaCSR[ 170 ][ 270 ],
   alphaCSR[ 170 ][ 271 ],
   alphaCSR[ 170 ][ 272 ],
   alphaCSR[ 170 ][ 273 ],
   alphaCSR[ 170 ][ 274 ],
   alphaCSR[ 170 ][ 275 ],
   alphaCSR[ 170 ][ 276 ],
   alphaCSR[ 170 ][ 277 ],
   alphaCSR[ 170 ][ 278 ],
   alphaCSR[ 170 ][ 279 ],
   alphaCSR[ 170 ][ 280 ],
   alphaCSR[ 170 ][ 281 ],
   alphaCSR[ 170 ][ 282 ],
   alphaCSR[ 170 ][ 283 ],
   alphaCSR[ 170 ][ 284 ],
   alphaCSR[ 170 ][ 285 ],
   alphaCSR[ 170 ][ 286 ],
   alphaCSR[ 170 ][ 287 ],
   alphaCSR[ 170 ][ 288 ],
   alphaCSR[ 170 ][ 289 ],
   alphaCSR[ 170 ][ 290 ],
   alphaCSR[ 170 ][ 291 ],
   alphaCSR[ 170 ][ 292 ],
   alphaCSR[ 170 ][ 293 ],
   alphaCSR[ 170 ][ 294 ],
   alphaCSR[ 170 ][ 295 ],
   alphaCSR[ 170 ][ 296 ],
   alphaCSR[ 170 ][ 297 ],
   alphaCSR[ 170 ][ 298 ],
   alphaCSR[ 170 ][ 299 ],
   alphaCSR[ 170 ][ 300 ],
   alphaCSR[ 170 ][ 301 ],
   alphaCSR[ 170 ][ 302 ],
   alphaCSR[ 170 ][ 303 ],
   alphaCSR[ 170 ][ 304 ],
   alphaCSR[ 170 ][ 305 ],
   alphaCSR[ 170 ][ 306 ],
   alphaCSR[ 170 ][ 307 ],
   alphaCSR[ 170 ][ 308 ],
   alphaCSR[ 170 ][ 309 ],
   alphaCSR[ 170 ][ 310 ],
   alphaCSR[ 170 ][ 311 ],
   alphaCSR[ 170 ][ 312 ],
   alphaCSR[ 170 ][ 313 ],
   alphaCSR[ 170 ][ 314 ],
   alphaCSR[ 170 ][ 315 ],
   alphaCSR[ 170 ][ 316 ],
   alphaCSR[ 170 ][ 317 ],
   alphaCSR[ 170 ][ 318 ],
   alphaCSR[ 170 ][ 319 ],
   alphaCSR[ 170 ][ 320 ],
   alphaCSR[ 170 ][ 321 ],
   alphaCSR[ 170 ][ 322 ],
   alphaCSR[ 170 ][ 323 ],
   alphaCSR[ 170 ][ 324 ],
   alphaCSR[ 170 ][ 325 ],
   alphaCSR[ 170 ][ 326 ],
   alphaCSR[ 170 ][ 327 ],
   alphaCSR[ 170 ][ 328 ],
   alphaCSR[ 170 ][ 329 ],
   alphaCSR[ 170 ][ 330 ],
   alphaCSR[ 170 ][ 331 ],
   alphaCSR[ 170 ][ 332 ],
   alphaCSR[ 170 ][ 333 ],
   alphaCSR[ 170 ][ 334 ],
   alphaCSR[ 170 ][ 335 ],
   alphaCSR[ 170 ][ 336 ],
   alphaCSR[ 170 ][ 337 ],
   alphaCSR[ 170 ][ 338 ],
   alphaCSR[ 170 ][ 339 ],
   alphaCSR[ 170 ][ 340 ],
   alphaCSR[ 170 ][ 341 ],
   alphaCSR[ 170 ][ 342 ],
   alphaCSR[ 170 ][ 343 ],
   alphaCSR[ 170 ][ 344 ],
   alphaCSR[ 170 ][ 345 ],
   alphaCSR[ 170 ][ 346 ],
   alphaCSR[ 170 ][ 347 ],
   alphaCSR[ 170 ][ 348 ],
   alphaCSR[ 170 ][ 349 ],
   alphaCSR[ 170 ][ 350 ],
   alphaCSR[ 170 ][ 351 ],
   alphaCSR[ 170 ][ 352 ],
   alphaCSR[ 170 ][ 353 ],
   alphaCSR[ 170 ][ 354 ],
   alphaCSR[ 170 ][ 355 ],
   alphaCSR[ 170 ][ 356 ],
   alphaCSR[ 170 ][ 357 ],
   alphaCSR[ 170 ][ 358 ],
   alphaCSR[ 170 ][ 359 ],
   alphaCSR[ 170 ][ 360 ],
   alphaCSR[ 170 ][ 361 ],
   alphaCSR[ 170 ][ 362 ],
   alphaCSR[ 170 ][ 363 ],
   alphaCSR[ 170 ][ 364 ],
   alphaCSR[ 170 ][ 365 ],
   alphaCSR[ 170 ][ 366 ],
   alphaCSR[ 170 ][ 367 ],
   alphaCSR[ 170 ][ 368 ],
   alphaCSR[ 170 ][ 369 ],
   alphaCSR[ 170 ][ 370 ],
   alphaCSR[ 170 ][ 371 ],
   alphaCSR[ 170 ][ 372 ],
   alphaCSR[ 170 ][ 373 ],
   alphaCSR[ 170 ][ 374 ],
   alphaCSR[ 170 ][ 375 ],
   alphaCSR[ 170 ][ 376 ],
   alphaCSR[ 170 ][ 377 ],
   alphaCSR[ 170 ][ 378 ],
   alphaCSR[ 170 ][ 379 ],
   alphaCSR[ 170 ][ 380 ],
   alphaCSR[ 170 ][ 381 ],
   alphaCSR[ 170 ][ 382 ],
   alphaCSR[ 170 ][ 383 ],
   alphaCSR[ 171 ][ 0 ],
   alphaCSR[ 171 ][ 1 ],
   alphaCSR[ 171 ][ 2 ],
   alphaCSR[ 171 ][ 3 ],
   alphaCSR[ 171 ][ 4 ],
   alphaCSR[ 171 ][ 5 ],
   alphaCSR[ 171 ][ 6 ],
   alphaCSR[ 171 ][ 7 ],
   alphaCSR[ 171 ][ 8 ],
   alphaCSR[ 171 ][ 9 ],
   alphaCSR[ 171 ][ 10 ],
   alphaCSR[ 171 ][ 11 ],
   alphaCSR[ 171 ][ 12 ],
   alphaCSR[ 171 ][ 13 ],
   alphaCSR[ 171 ][ 14 ],
   alphaCSR[ 171 ][ 15 ],
   alphaCSR[ 171 ][ 16 ],
   alphaCSR[ 171 ][ 17 ],
   alphaCSR[ 171 ][ 18 ],
   alphaCSR[ 171 ][ 19 ],
   alphaCSR[ 171 ][ 20 ],
   alphaCSR[ 171 ][ 21 ],
   alphaCSR[ 171 ][ 22 ],
   alphaCSR[ 171 ][ 23 ],
   alphaCSR[ 171 ][ 24 ],
   alphaCSR[ 171 ][ 25 ],
   alphaCSR[ 171 ][ 26 ],
   alphaCSR[ 171 ][ 27 ],
   alphaCSR[ 171 ][ 28 ],
   alphaCSR[ 171 ][ 29 ],
   alphaCSR[ 171 ][ 30 ],
   alphaCSR[ 171 ][ 31 ],
   alphaCSR[ 171 ][ 32 ],
   alphaCSR[ 171 ][ 33 ],
   alphaCSR[ 171 ][ 34 ],
   alphaCSR[ 171 ][ 35 ],
   alphaCSR[ 171 ][ 36 ],
   alphaCSR[ 171 ][ 37 ],
   alphaCSR[ 171 ][ 38 ],
   alphaCSR[ 171 ][ 39 ],
   alphaCSR[ 171 ][ 40 ],
   alphaCSR[ 171 ][ 41 ],
   alphaCSR[ 171 ][ 42 ],
   alphaCSR[ 171 ][ 43 ],
   alphaCSR[ 171 ][ 44 ],
   alphaCSR[ 171 ][ 45 ],
   alphaCSR[ 171 ][ 46 ],
   alphaCSR[ 171 ][ 47 ],
   alphaCSR[ 171 ][ 48 ],
   alphaCSR[ 171 ][ 49 ],
   alphaCSR[ 171 ][ 50 ],
   alphaCSR[ 171 ][ 51 ],
   alphaCSR[ 171 ][ 52 ],
   alphaCSR[ 171 ][ 53 ],
   alphaCSR[ 171 ][ 54 ],
   alphaCSR[ 171 ][ 55 ],
   alphaCSR[ 171 ][ 56 ],
   alphaCSR[ 171 ][ 57 ],
   alphaCSR[ 171 ][ 58 ],
   alphaCSR[ 171 ][ 59 ],
   alphaCSR[ 171 ][ 60 ],
   alphaCSR[ 171 ][ 61 ],
   alphaCSR[ 171 ][ 62 ],
   alphaCSR[ 171 ][ 63 ],
   alphaCSR[ 171 ][ 64 ],
   alphaCSR[ 171 ][ 65 ],
   alphaCSR[ 171 ][ 66 ],
   alphaCSR[ 171 ][ 67 ],
   alphaCSR[ 171 ][ 68 ],
   alphaCSR[ 171 ][ 69 ],
   alphaCSR[ 171 ][ 70 ],
   alphaCSR[ 171 ][ 71 ],
   alphaCSR[ 171 ][ 72 ],
   alphaCSR[ 171 ][ 73 ],
   alphaCSR[ 171 ][ 74 ],
   alphaCSR[ 171 ][ 75 ],
   alphaCSR[ 171 ][ 76 ],
   alphaCSR[ 171 ][ 77 ],
   alphaCSR[ 171 ][ 78 ],
   alphaCSR[ 171 ][ 79 ],
   alphaCSR[ 171 ][ 80 ],
   alphaCSR[ 171 ][ 81 ],
   alphaCSR[ 171 ][ 82 ],
   alphaCSR[ 171 ][ 83 ],
   alphaCSR[ 171 ][ 84 ],
   alphaCSR[ 171 ][ 85 ],
   alphaCSR[ 171 ][ 86 ],
   alphaCSR[ 171 ][ 87 ],
   alphaCSR[ 171 ][ 88 ],
   alphaCSR[ 171 ][ 89 ],
   alphaCSR[ 171 ][ 90 ],
   alphaCSR[ 171 ][ 91 ],
   alphaCSR[ 171 ][ 92 ],
   alphaCSR[ 171 ][ 93 ],
   alphaCSR[ 171 ][ 94 ],
   alphaCSR[ 171 ][ 95 ],
   alphaCSR[ 171 ][ 96 ],
   alphaCSR[ 171 ][ 97 ],
   alphaCSR[ 171 ][ 98 ],
   alphaCSR[ 171 ][ 99 ],
   alphaCSR[ 171 ][ 100 ],
   alphaCSR[ 171 ][ 101 ],
   alphaCSR[ 171 ][ 102 ],
   alphaCSR[ 171 ][ 103 ],
   alphaCSR[ 171 ][ 104 ],
   alphaCSR[ 171 ][ 105 ],
   alphaCSR[ 171 ][ 106 ],
   alphaCSR[ 171 ][ 107 ],
   alphaCSR[ 171 ][ 108 ],
   alphaCSR[ 171 ][ 109 ],
   alphaCSR[ 171 ][ 110 ],
   alphaCSR[ 171 ][ 111 ],
   alphaCSR[ 171 ][ 112 ],
   alphaCSR[ 171 ][ 113 ],
   alphaCSR[ 171 ][ 114 ],
   alphaCSR[ 171 ][ 115 ],
   alphaCSR[ 171 ][ 116 ],
   alphaCSR[ 171 ][ 117 ],
   alphaCSR[ 171 ][ 118 ],
   alphaCSR[ 171 ][ 119 ],
   alphaCSR[ 171 ][ 120 ],
   alphaCSR[ 171 ][ 121 ],
   alphaCSR[ 171 ][ 122 ],
   alphaCSR[ 171 ][ 123 ],
   alphaCSR[ 171 ][ 124 ],
   alphaCSR[ 171 ][ 125 ],
   alphaCSR[ 171 ][ 126 ],
   alphaCSR[ 171 ][ 127 ],
   alphaCSR[ 171 ][ 128 ],
   alphaCSR[ 171 ][ 129 ],
   alphaCSR[ 171 ][ 130 ],
   alphaCSR[ 171 ][ 131 ],
   alphaCSR[ 171 ][ 132 ],
   alphaCSR[ 171 ][ 133 ],
   alphaCSR[ 171 ][ 134 ],
   alphaCSR[ 171 ][ 135 ],
   alphaCSR[ 171 ][ 136 ],
   alphaCSR[ 171 ][ 137 ],
   alphaCSR[ 171 ][ 138 ],
   alphaCSR[ 171 ][ 139 ],
   alphaCSR[ 171 ][ 140 ],
   alphaCSR[ 171 ][ 141 ],
   alphaCSR[ 171 ][ 142 ],
   alphaCSR[ 171 ][ 143 ],
   alphaCSR[ 171 ][ 144 ],
   alphaCSR[ 171 ][ 145 ],
   alphaCSR[ 171 ][ 146 ],
   alphaCSR[ 171 ][ 147 ],
   alphaCSR[ 171 ][ 148 ],
   alphaCSR[ 171 ][ 149 ],
   alphaCSR[ 171 ][ 150 ],
   alphaCSR[ 171 ][ 151 ],
   alphaCSR[ 171 ][ 152 ],
   alphaCSR[ 171 ][ 153 ],
   alphaCSR[ 171 ][ 154 ],
   alphaCSR[ 171 ][ 155 ],
   alphaCSR[ 171 ][ 156 ],
   alphaCSR[ 171 ][ 157 ],
   alphaCSR[ 171 ][ 158 ],
   alphaCSR[ 171 ][ 159 ],
   alphaCSR[ 171 ][ 160 ],
   alphaCSR[ 171 ][ 161 ],
   alphaCSR[ 171 ][ 162 ],
   alphaCSR[ 171 ][ 163 ],
   alphaCSR[ 171 ][ 164 ],
   alphaCSR[ 171 ][ 165 ],
   alphaCSR[ 171 ][ 166 ],
   alphaCSR[ 171 ][ 167 ],
   alphaCSR[ 171 ][ 168 ],
   alphaCSR[ 171 ][ 169 ],
   alphaCSR[ 171 ][ 170 ],
   alphaCSR[ 171 ][ 171 ],
   alphaCSR[ 171 ][ 172 ],
   alphaCSR[ 171 ][ 173 ],
   alphaCSR[ 171 ][ 174 ],
   alphaCSR[ 171 ][ 175 ],
   alphaCSR[ 171 ][ 176 ],
   alphaCSR[ 171 ][ 177 ],
   alphaCSR[ 171 ][ 178 ],
   alphaCSR[ 171 ][ 179 ],
   alphaCSR[ 171 ][ 180 ],
   alphaCSR[ 171 ][ 181 ],
   alphaCSR[ 171 ][ 182 ],
   alphaCSR[ 171 ][ 183 ],
   alphaCSR[ 171 ][ 184 ],
   alphaCSR[ 171 ][ 185 ],
   alphaCSR[ 171 ][ 186 ],
   alphaCSR[ 171 ][ 187 ],
   alphaCSR[ 171 ][ 188 ],
   alphaCSR[ 171 ][ 189 ],
   alphaCSR[ 171 ][ 190 ],
   alphaCSR[ 171 ][ 191 ],
   alphaCSR[ 171 ][ 192 ],
   alphaCSR[ 171 ][ 193 ],
   alphaCSR[ 171 ][ 194 ],
   alphaCSR[ 171 ][ 195 ],
   alphaCSR[ 171 ][ 196 ],
   alphaCSR[ 171 ][ 197 ],
   alphaCSR[ 171 ][ 198 ],
   alphaCSR[ 171 ][ 199 ],
   alphaCSR[ 171 ][ 200 ],
   alphaCSR[ 171 ][ 201 ],
   alphaCSR[ 171 ][ 202 ],
   alphaCSR[ 171 ][ 203 ],
   alphaCSR[ 171 ][ 204 ],
   alphaCSR[ 171 ][ 205 ],
   alphaCSR[ 171 ][ 206 ],
   alphaCSR[ 171 ][ 207 ],
   alphaCSR[ 171 ][ 208 ],
   alphaCSR[ 171 ][ 209 ],
   alphaCSR[ 171 ][ 210 ],
   alphaCSR[ 171 ][ 211 ],
   alphaCSR[ 171 ][ 212 ],
   alphaCSR[ 171 ][ 213 ],
   alphaCSR[ 171 ][ 214 ],
   alphaCSR[ 171 ][ 215 ],
   alphaCSR[ 171 ][ 216 ],
   alphaCSR[ 171 ][ 217 ],
   alphaCSR[ 171 ][ 218 ],
   alphaCSR[ 171 ][ 219 ],
   alphaCSR[ 171 ][ 220 ],
   alphaCSR[ 171 ][ 221 ],
   alphaCSR[ 171 ][ 222 ],
   alphaCSR[ 171 ][ 223 ],
   alphaCSR[ 171 ][ 224 ],
   alphaCSR[ 171 ][ 225 ],
   alphaCSR[ 171 ][ 226 ],
   alphaCSR[ 171 ][ 227 ],
   alphaCSR[ 171 ][ 228 ],
   alphaCSR[ 171 ][ 229 ],
   alphaCSR[ 171 ][ 230 ],
   alphaCSR[ 171 ][ 231 ],
   alphaCSR[ 171 ][ 232 ],
   alphaCSR[ 171 ][ 233 ],
   alphaCSR[ 171 ][ 234 ],
   alphaCSR[ 171 ][ 235 ],
   alphaCSR[ 171 ][ 236 ],
   alphaCSR[ 171 ][ 237 ],
   alphaCSR[ 171 ][ 238 ],
   alphaCSR[ 171 ][ 239 ],
   alphaCSR[ 171 ][ 240 ],
   alphaCSR[ 171 ][ 241 ],
   alphaCSR[ 171 ][ 242 ],
   alphaCSR[ 171 ][ 243 ],
   alphaCSR[ 171 ][ 244 ],
   alphaCSR[ 171 ][ 245 ],
   alphaCSR[ 171 ][ 246 ],
   alphaCSR[ 171 ][ 247 ],
   alphaCSR[ 171 ][ 248 ],
   alphaCSR[ 171 ][ 249 ],
   alphaCSR[ 171 ][ 250 ],
   alphaCSR[ 171 ][ 251 ],
   alphaCSR[ 171 ][ 252 ],
   alphaCSR[ 171 ][ 253 ],
   alphaCSR[ 171 ][ 254 ],
   alphaCSR[ 171 ][ 255 ],
   alphaCSR[ 171 ][ 256 ],
   alphaCSR[ 171 ][ 257 ],
   alphaCSR[ 171 ][ 258 ],
   alphaCSR[ 171 ][ 259 ],
   alphaCSR[ 171 ][ 260 ],
   alphaCSR[ 171 ][ 261 ],
   alphaCSR[ 171 ][ 262 ],
   alphaCSR[ 171 ][ 263 ],
   alphaCSR[ 171 ][ 264 ],
   alphaCSR[ 171 ][ 265 ],
   alphaCSR[ 171 ][ 266 ],
   alphaCSR[ 171 ][ 267 ],
   alphaCSR[ 171 ][ 268 ],
   alphaCSR[ 171 ][ 269 ],
   alphaCSR[ 171 ][ 270 ],
   alphaCSR[ 171 ][ 271 ],
   alphaCSR[ 171 ][ 272 ],
   alphaCSR[ 171 ][ 273 ],
   alphaCSR[ 171 ][ 274 ],
   alphaCSR[ 171 ][ 275 ],
   alphaCSR[ 171 ][ 276 ],
   alphaCSR[ 171 ][ 277 ],
   alphaCSR[ 171 ][ 278 ],
   alphaCSR[ 171 ][ 279 ],
   alphaCSR[ 171 ][ 280 ],
   alphaCSR[ 171 ][ 281 ],
   alphaCSR[ 171 ][ 282 ],
   alphaCSR[ 171 ][ 283 ],
   alphaCSR[ 171 ][ 284 ],
   alphaCSR[ 171 ][ 285 ],
   alphaCSR[ 171 ][ 286 ],
   alphaCSR[ 171 ][ 287 ],
   alphaCSR[ 171 ][ 288 ],
   alphaCSR[ 171 ][ 289 ],
   alphaCSR[ 171 ][ 290 ],
   alphaCSR[ 171 ][ 291 ],
   alphaCSR[ 171 ][ 292 ],
   alphaCSR[ 171 ][ 293 ],
   alphaCSR[ 171 ][ 294 ],
   alphaCSR[ 171 ][ 295 ],
   alphaCSR[ 171 ][ 296 ],
   alphaCSR[ 171 ][ 297 ],
   alphaCSR[ 171 ][ 298 ],
   alphaCSR[ 171 ][ 299 ],
   alphaCSR[ 171 ][ 300 ],
   alphaCSR[ 171 ][ 301 ],
   alphaCSR[ 171 ][ 302 ],
   alphaCSR[ 171 ][ 303 ],
   alphaCSR[ 171 ][ 304 ],
   alphaCSR[ 171 ][ 305 ],
   alphaCSR[ 171 ][ 306 ],
   alphaCSR[ 171 ][ 307 ],
   alphaCSR[ 171 ][ 308 ],
   alphaCSR[ 171 ][ 309 ],
   alphaCSR[ 171 ][ 310 ],
   alphaCSR[ 171 ][ 311 ],
   alphaCSR[ 171 ][ 312 ],
   alphaCSR[ 171 ][ 313 ],
   alphaCSR[ 171 ][ 314 ],
   alphaCSR[ 171 ][ 315 ],
   alphaCSR[ 171 ][ 316 ],
   alphaCSR[ 171 ][ 317 ],
   alphaCSR[ 171 ][ 318 ],
   alphaCSR[ 171 ][ 319 ],
   alphaCSR[ 171 ][ 320 ],
   alphaCSR[ 171 ][ 321 ],
   alphaCSR[ 171 ][ 322 ],
   alphaCSR[ 171 ][ 323 ],
   alphaCSR[ 171 ][ 324 ],
   alphaCSR[ 171 ][ 325 ],
   alphaCSR[ 171 ][ 326 ],
   alphaCSR[ 171 ][ 327 ],
   alphaCSR[ 171 ][ 328 ],
   alphaCSR[ 171 ][ 329 ],
   alphaCSR[ 171 ][ 330 ],
   alphaCSR[ 171 ][ 331 ],
   alphaCSR[ 171 ][ 332 ],
   alphaCSR[ 171 ][ 333 ],
   alphaCSR[ 171 ][ 334 ],
   alphaCSR[ 171 ][ 335 ],
   alphaCSR[ 171 ][ 336 ],
   alphaCSR[ 171 ][ 337 ],
   alphaCSR[ 171 ][ 338 ],
   alphaCSR[ 171 ][ 339 ],
   alphaCSR[ 171 ][ 340 ],
   alphaCSR[ 171 ][ 341 ],
   alphaCSR[ 171 ][ 342 ],
   alphaCSR[ 171 ][ 343 ],
   alphaCSR[ 171 ][ 344 ],
   alphaCSR[ 171 ][ 345 ],
   alphaCSR[ 171 ][ 346 ],
   alphaCSR[ 171 ][ 347 ],
   alphaCSR[ 171 ][ 348 ],
   alphaCSR[ 171 ][ 349 ],
   alphaCSR[ 171 ][ 350 ],
   alphaCSR[ 171 ][ 351 ],
   alphaCSR[ 171 ][ 352 ],
   alphaCSR[ 171 ][ 353 ],
   alphaCSR[ 171 ][ 354 ],
   alphaCSR[ 171 ][ 355 ],
   alphaCSR[ 171 ][ 356 ],
   alphaCSR[ 171 ][ 357 ],
   alphaCSR[ 171 ][ 358 ],
   alphaCSR[ 171 ][ 359 ],
   alphaCSR[ 171 ][ 360 ],
   alphaCSR[ 171 ][ 361 ],
   alphaCSR[ 171 ][ 362 ],
   alphaCSR[ 171 ][ 363 ],
   alphaCSR[ 171 ][ 364 ],
   alphaCSR[ 171 ][ 365 ],
   alphaCSR[ 171 ][ 366 ],
   alphaCSR[ 171 ][ 367 ],
   alphaCSR[ 171 ][ 368 ],
   alphaCSR[ 171 ][ 369 ],
   alphaCSR[ 171 ][ 370 ],
   alphaCSR[ 171 ][ 371 ],
   alphaCSR[ 171 ][ 372 ],
   alphaCSR[ 171 ][ 373 ],
   alphaCSR[ 171 ][ 374 ],
   alphaCSR[ 171 ][ 375 ],
   alphaCSR[ 171 ][ 376 ],
   alphaCSR[ 171 ][ 377 ],
   alphaCSR[ 171 ][ 378 ],
   alphaCSR[ 171 ][ 379 ],
   alphaCSR[ 171 ][ 380 ],
   alphaCSR[ 171 ][ 381 ],
   alphaCSR[ 171 ][ 382 ],
   alphaCSR[ 171 ][ 383 ],
   alphaCSR[ 172 ][ 0 ],
   alphaCSR[ 172 ][ 1 ],
   alphaCSR[ 172 ][ 2 ],
   alphaCSR[ 172 ][ 3 ],
   alphaCSR[ 172 ][ 4 ],
   alphaCSR[ 172 ][ 5 ],
   alphaCSR[ 172 ][ 6 ],
   alphaCSR[ 172 ][ 7 ],
   alphaCSR[ 172 ][ 8 ],
   alphaCSR[ 172 ][ 9 ],
   alphaCSR[ 172 ][ 10 ],
   alphaCSR[ 172 ][ 11 ],
   alphaCSR[ 172 ][ 12 ],
   alphaCSR[ 172 ][ 13 ],
   alphaCSR[ 172 ][ 14 ],
   alphaCSR[ 172 ][ 15 ],
   alphaCSR[ 172 ][ 16 ],
   alphaCSR[ 172 ][ 17 ],
   alphaCSR[ 172 ][ 18 ],
   alphaCSR[ 172 ][ 19 ],
   alphaCSR[ 172 ][ 20 ],
   alphaCSR[ 172 ][ 21 ],
   alphaCSR[ 172 ][ 22 ],
   alphaCSR[ 172 ][ 23 ],
   alphaCSR[ 172 ][ 24 ],
   alphaCSR[ 172 ][ 25 ],
   alphaCSR[ 172 ][ 26 ],
   alphaCSR[ 172 ][ 27 ],
   alphaCSR[ 172 ][ 28 ],
   alphaCSR[ 172 ][ 29 ],
   alphaCSR[ 172 ][ 30 ],
   alphaCSR[ 172 ][ 31 ],
   alphaCSR[ 172 ][ 32 ],
   alphaCSR[ 172 ][ 33 ],
   alphaCSR[ 172 ][ 34 ],
   alphaCSR[ 172 ][ 35 ],
   alphaCSR[ 172 ][ 36 ],
   alphaCSR[ 172 ][ 37 ],
   alphaCSR[ 172 ][ 38 ],
   alphaCSR[ 172 ][ 39 ],
   alphaCSR[ 172 ][ 40 ],
   alphaCSR[ 172 ][ 41 ],
   alphaCSR[ 172 ][ 42 ],
   alphaCSR[ 172 ][ 43 ],
   alphaCSR[ 172 ][ 44 ],
   alphaCSR[ 172 ][ 45 ],
   alphaCSR[ 172 ][ 46 ],
   alphaCSR[ 172 ][ 47 ],
   alphaCSR[ 172 ][ 48 ],
   alphaCSR[ 172 ][ 49 ],
   alphaCSR[ 172 ][ 50 ],
   alphaCSR[ 172 ][ 51 ],
   alphaCSR[ 172 ][ 52 ],
   alphaCSR[ 172 ][ 53 ],
   alphaCSR[ 172 ][ 54 ],
   alphaCSR[ 172 ][ 55 ],
   alphaCSR[ 172 ][ 56 ],
   alphaCSR[ 172 ][ 57 ],
   alphaCSR[ 172 ][ 58 ],
   alphaCSR[ 172 ][ 59 ],
   alphaCSR[ 172 ][ 60 ],
   alphaCSR[ 172 ][ 61 ],
   alphaCSR[ 172 ][ 62 ],
   alphaCSR[ 172 ][ 63 ],
   alphaCSR[ 172 ][ 64 ],
   alphaCSR[ 172 ][ 65 ],
   alphaCSR[ 172 ][ 66 ],
   alphaCSR[ 172 ][ 67 ],
   alphaCSR[ 172 ][ 68 ],
   alphaCSR[ 172 ][ 69 ],
   alphaCSR[ 172 ][ 70 ],
   alphaCSR[ 172 ][ 71 ],
   alphaCSR[ 172 ][ 72 ],
   alphaCSR[ 172 ][ 73 ],
   alphaCSR[ 172 ][ 74 ],
   alphaCSR[ 172 ][ 75 ],
   alphaCSR[ 172 ][ 76 ],
   alphaCSR[ 172 ][ 77 ],
   alphaCSR[ 172 ][ 78 ],
   alphaCSR[ 172 ][ 79 ],
   alphaCSR[ 172 ][ 80 ],
   alphaCSR[ 172 ][ 81 ],
   alphaCSR[ 172 ][ 82 ],
   alphaCSR[ 172 ][ 83 ],
   alphaCSR[ 172 ][ 84 ],
   alphaCSR[ 172 ][ 85 ],
   alphaCSR[ 172 ][ 86 ],
   alphaCSR[ 172 ][ 87 ],
   alphaCSR[ 172 ][ 88 ],
   alphaCSR[ 172 ][ 89 ],
   alphaCSR[ 172 ][ 90 ],
   alphaCSR[ 172 ][ 91 ],
   alphaCSR[ 172 ][ 92 ],
   alphaCSR[ 172 ][ 93 ],
   alphaCSR[ 172 ][ 94 ],
   alphaCSR[ 172 ][ 95 ],
   alphaCSR[ 172 ][ 96 ],
   alphaCSR[ 172 ][ 97 ],
   alphaCSR[ 172 ][ 98 ],
   alphaCSR[ 172 ][ 99 ],
   alphaCSR[ 172 ][ 100 ],
   alphaCSR[ 172 ][ 101 ],
   alphaCSR[ 172 ][ 102 ],
   alphaCSR[ 172 ][ 103 ],
   alphaCSR[ 172 ][ 104 ],
   alphaCSR[ 172 ][ 105 ],
   alphaCSR[ 172 ][ 106 ],
   alphaCSR[ 172 ][ 107 ],
   alphaCSR[ 172 ][ 108 ],
   alphaCSR[ 172 ][ 109 ],
   alphaCSR[ 172 ][ 110 ],
   alphaCSR[ 172 ][ 111 ],
   alphaCSR[ 172 ][ 112 ],
   alphaCSR[ 172 ][ 113 ],
   alphaCSR[ 172 ][ 114 ],
   alphaCSR[ 172 ][ 115 ],
   alphaCSR[ 172 ][ 116 ],
   alphaCSR[ 172 ][ 117 ],
   alphaCSR[ 172 ][ 118 ],
   alphaCSR[ 172 ][ 119 ],
   alphaCSR[ 172 ][ 120 ],
   alphaCSR[ 172 ][ 121 ],
   alphaCSR[ 172 ][ 122 ],
   alphaCSR[ 172 ][ 123 ],
   alphaCSR[ 172 ][ 124 ],
   alphaCSR[ 172 ][ 125 ],
   alphaCSR[ 172 ][ 126 ],
   alphaCSR[ 172 ][ 127 ],
   alphaCSR[ 172 ][ 128 ],
   alphaCSR[ 172 ][ 129 ],
   alphaCSR[ 172 ][ 130 ],
   alphaCSR[ 172 ][ 131 ],
   alphaCSR[ 172 ][ 132 ],
   alphaCSR[ 172 ][ 133 ],
   alphaCSR[ 172 ][ 134 ],
   alphaCSR[ 172 ][ 135 ],
   alphaCSR[ 172 ][ 136 ],
   alphaCSR[ 172 ][ 137 ],
   alphaCSR[ 172 ][ 138 ],
   alphaCSR[ 172 ][ 139 ],
   alphaCSR[ 172 ][ 140 ],
   alphaCSR[ 172 ][ 141 ],
   alphaCSR[ 172 ][ 142 ],
   alphaCSR[ 172 ][ 143 ],
   alphaCSR[ 172 ][ 144 ],
   alphaCSR[ 172 ][ 145 ],
   alphaCSR[ 172 ][ 146 ],
   alphaCSR[ 172 ][ 147 ],
   alphaCSR[ 172 ][ 148 ],
   alphaCSR[ 172 ][ 149 ],
   alphaCSR[ 172 ][ 150 ],
   alphaCSR[ 172 ][ 151 ],
   alphaCSR[ 172 ][ 152 ],
   alphaCSR[ 172 ][ 153 ],
   alphaCSR[ 172 ][ 154 ],
   alphaCSR[ 172 ][ 155 ],
   alphaCSR[ 172 ][ 156 ],
   alphaCSR[ 172 ][ 157 ],
   alphaCSR[ 172 ][ 158 ],
   alphaCSR[ 172 ][ 159 ],
   alphaCSR[ 172 ][ 160 ],
   alphaCSR[ 172 ][ 161 ],
   alphaCSR[ 172 ][ 162 ],
   alphaCSR[ 172 ][ 163 ],
   alphaCSR[ 172 ][ 164 ],
   alphaCSR[ 172 ][ 165 ],
   alphaCSR[ 172 ][ 166 ],
   alphaCSR[ 172 ][ 167 ],
   alphaCSR[ 172 ][ 168 ],
   alphaCSR[ 172 ][ 169 ],
   alphaCSR[ 172 ][ 170 ],
   alphaCSR[ 172 ][ 171 ],
   alphaCSR[ 172 ][ 172 ],
   alphaCSR[ 172 ][ 173 ],
   alphaCSR[ 172 ][ 174 ],
   alphaCSR[ 172 ][ 175 ],
   alphaCSR[ 172 ][ 176 ],
   alphaCSR[ 172 ][ 177 ],
   alphaCSR[ 172 ][ 178 ],
   alphaCSR[ 172 ][ 179 ],
   alphaCSR[ 172 ][ 180 ],
   alphaCSR[ 172 ][ 181 ],
   alphaCSR[ 172 ][ 182 ],
   alphaCSR[ 172 ][ 183 ],
   alphaCSR[ 172 ][ 184 ],
   alphaCSR[ 172 ][ 185 ],
   alphaCSR[ 172 ][ 186 ],
   alphaCSR[ 172 ][ 187 ],
   alphaCSR[ 172 ][ 188 ],
   alphaCSR[ 172 ][ 189 ],
   alphaCSR[ 172 ][ 190 ],
   alphaCSR[ 172 ][ 191 ],
   alphaCSR[ 172 ][ 192 ],
   alphaCSR[ 172 ][ 193 ],
   alphaCSR[ 172 ][ 194 ],
   alphaCSR[ 172 ][ 195 ],
   alphaCSR[ 172 ][ 196 ],
   alphaCSR[ 172 ][ 197 ],
   alphaCSR[ 172 ][ 198 ],
   alphaCSR[ 172 ][ 199 ],
   alphaCSR[ 172 ][ 200 ],
   alphaCSR[ 172 ][ 201 ],
   alphaCSR[ 172 ][ 202 ],
   alphaCSR[ 172 ][ 203 ],
   alphaCSR[ 172 ][ 204 ],
   alphaCSR[ 172 ][ 205 ],
   alphaCSR[ 172 ][ 206 ],
   alphaCSR[ 172 ][ 207 ],
   alphaCSR[ 172 ][ 208 ],
   alphaCSR[ 172 ][ 209 ],
   alphaCSR[ 172 ][ 210 ],
   alphaCSR[ 172 ][ 211 ],
   alphaCSR[ 172 ][ 212 ],
   alphaCSR[ 172 ][ 213 ],
   alphaCSR[ 172 ][ 214 ],
   alphaCSR[ 172 ][ 215 ],
   alphaCSR[ 172 ][ 216 ],
   alphaCSR[ 172 ][ 217 ],
   alphaCSR[ 172 ][ 218 ],
   alphaCSR[ 172 ][ 219 ],
   alphaCSR[ 172 ][ 220 ],
   alphaCSR[ 172 ][ 221 ],
   alphaCSR[ 172 ][ 222 ],
   alphaCSR[ 172 ][ 223 ],
   alphaCSR[ 172 ][ 224 ],
   alphaCSR[ 172 ][ 225 ],
   alphaCSR[ 172 ][ 226 ],
   alphaCSR[ 172 ][ 227 ],
   alphaCSR[ 172 ][ 228 ],
   alphaCSR[ 172 ][ 229 ],
   alphaCSR[ 172 ][ 230 ],
   alphaCSR[ 172 ][ 231 ],
   alphaCSR[ 172 ][ 232 ],
   alphaCSR[ 172 ][ 233 ],
   alphaCSR[ 172 ][ 234 ],
   alphaCSR[ 172 ][ 235 ],
   alphaCSR[ 172 ][ 236 ],
   alphaCSR[ 172 ][ 237 ],
   alphaCSR[ 172 ][ 238 ],
   alphaCSR[ 172 ][ 239 ],
   alphaCSR[ 172 ][ 240 ],
   alphaCSR[ 172 ][ 241 ],
   alphaCSR[ 172 ][ 242 ],
   alphaCSR[ 172 ][ 243 ],
   alphaCSR[ 172 ][ 244 ],
   alphaCSR[ 172 ][ 245 ],
   alphaCSR[ 172 ][ 246 ],
   alphaCSR[ 172 ][ 247 ],
   alphaCSR[ 172 ][ 248 ],
   alphaCSR[ 172 ][ 249 ],
   alphaCSR[ 172 ][ 250 ],
   alphaCSR[ 172 ][ 251 ],
   alphaCSR[ 172 ][ 252 ],
   alphaCSR[ 172 ][ 253 ],
   alphaCSR[ 172 ][ 254 ],
   alphaCSR[ 172 ][ 255 ],
   alphaCSR[ 172 ][ 256 ],
   alphaCSR[ 172 ][ 257 ],
   alphaCSR[ 172 ][ 258 ],
   alphaCSR[ 172 ][ 259 ],
   alphaCSR[ 172 ][ 260 ],
   alphaCSR[ 172 ][ 261 ],
   alphaCSR[ 172 ][ 262 ],
   alphaCSR[ 172 ][ 263 ],
   alphaCSR[ 172 ][ 264 ],
   alphaCSR[ 172 ][ 265 ],
   alphaCSR[ 172 ][ 266 ],
   alphaCSR[ 172 ][ 267 ],
   alphaCSR[ 172 ][ 268 ],
   alphaCSR[ 172 ][ 269 ],
   alphaCSR[ 172 ][ 270 ],
   alphaCSR[ 172 ][ 271 ],
   alphaCSR[ 172 ][ 272 ],
   alphaCSR[ 172 ][ 273 ],
   alphaCSR[ 172 ][ 274 ],
   alphaCSR[ 172 ][ 275 ],
   alphaCSR[ 172 ][ 276 ],
   alphaCSR[ 172 ][ 277 ],
   alphaCSR[ 172 ][ 278 ],
   alphaCSR[ 172 ][ 279 ],
   alphaCSR[ 172 ][ 280 ],
   alphaCSR[ 172 ][ 281 ],
   alphaCSR[ 172 ][ 282 ],
   alphaCSR[ 172 ][ 283 ],
   alphaCSR[ 172 ][ 284 ],
   alphaCSR[ 172 ][ 285 ],
   alphaCSR[ 172 ][ 286 ],
   alphaCSR[ 172 ][ 287 ],
   alphaCSR[ 172 ][ 288 ],
   alphaCSR[ 172 ][ 289 ],
   alphaCSR[ 172 ][ 290 ],
   alphaCSR[ 172 ][ 291 ],
   alphaCSR[ 172 ][ 292 ],
   alphaCSR[ 172 ][ 293 ],
   alphaCSR[ 172 ][ 294 ],
   alphaCSR[ 172 ][ 295 ],
   alphaCSR[ 172 ][ 296 ],
   alphaCSR[ 172 ][ 297 ],
   alphaCSR[ 172 ][ 298 ],
   alphaCSR[ 172 ][ 299 ],
   alphaCSR[ 172 ][ 300 ],
   alphaCSR[ 172 ][ 301 ],
   alphaCSR[ 172 ][ 302 ],
   alphaCSR[ 172 ][ 303 ],
   alphaCSR[ 172 ][ 304 ],
   alphaCSR[ 172 ][ 305 ],
   alphaCSR[ 172 ][ 306 ],
   alphaCSR[ 172 ][ 307 ],
   alphaCSR[ 172 ][ 308 ],
   alphaCSR[ 172 ][ 309 ],
   alphaCSR[ 172 ][ 310 ],
   alphaCSR[ 172 ][ 311 ],
   alphaCSR[ 172 ][ 312 ],
   alphaCSR[ 172 ][ 313 ],
   alphaCSR[ 172 ][ 314 ],
   alphaCSR[ 172 ][ 315 ],
   alphaCSR[ 172 ][ 316 ],
   alphaCSR[ 172 ][ 317 ],
   alphaCSR[ 172 ][ 318 ],
   alphaCSR[ 172 ][ 319 ],
   alphaCSR[ 172 ][ 320 ],
   alphaCSR[ 172 ][ 321 ],
   alphaCSR[ 172 ][ 322 ],
   alphaCSR[ 172 ][ 323 ],
   alphaCSR[ 172 ][ 324 ],
   alphaCSR[ 172 ][ 325 ],
   alphaCSR[ 172 ][ 326 ],
   alphaCSR[ 172 ][ 327 ],
   alphaCSR[ 172 ][ 328 ],
   alphaCSR[ 172 ][ 329 ],
   alphaCSR[ 172 ][ 330 ],
   alphaCSR[ 172 ][ 331 ],
   alphaCSR[ 172 ][ 332 ],
   alphaCSR[ 172 ][ 333 ],
   alphaCSR[ 172 ][ 334 ],
   alphaCSR[ 172 ][ 335 ],
   alphaCSR[ 172 ][ 336 ],
   alphaCSR[ 172 ][ 337 ],
   alphaCSR[ 172 ][ 338 ],
   alphaCSR[ 172 ][ 339 ],
   alphaCSR[ 172 ][ 340 ],
   alphaCSR[ 172 ][ 341 ],
   alphaCSR[ 172 ][ 342 ],
   alphaCSR[ 172 ][ 343 ],
   alphaCSR[ 172 ][ 344 ],
   alphaCSR[ 172 ][ 345 ],
   alphaCSR[ 172 ][ 346 ],
   alphaCSR[ 172 ][ 347 ],
   alphaCSR[ 172 ][ 348 ],
   alphaCSR[ 172 ][ 349 ],
   alphaCSR[ 172 ][ 350 ],
   alphaCSR[ 172 ][ 351 ],
   alphaCSR[ 172 ][ 352 ],
   alphaCSR[ 172 ][ 353 ],
   alphaCSR[ 172 ][ 354 ],
   alphaCSR[ 172 ][ 355 ],
   alphaCSR[ 172 ][ 356 ],
   alphaCSR[ 172 ][ 357 ],
   alphaCSR[ 172 ][ 358 ],
   alphaCSR[ 172 ][ 359 ],
   alphaCSR[ 172 ][ 360 ],
   alphaCSR[ 172 ][ 361 ],
   alphaCSR[ 172 ][ 362 ],
   alphaCSR[ 172 ][ 363 ],
   alphaCSR[ 172 ][ 364 ],
   alphaCSR[ 172 ][ 365 ],
   alphaCSR[ 172 ][ 366 ],
   alphaCSR[ 172 ][ 367 ],
   alphaCSR[ 172 ][ 368 ],
   alphaCSR[ 172 ][ 369 ],
   alphaCSR[ 172 ][ 370 ],
   alphaCSR[ 172 ][ 371 ],
   alphaCSR[ 172 ][ 372 ],
   alphaCSR[ 172 ][ 373 ],
   alphaCSR[ 172 ][ 374 ],
   alphaCSR[ 172 ][ 375 ],
   alphaCSR[ 172 ][ 376 ],
   alphaCSR[ 172 ][ 377 ],
   alphaCSR[ 172 ][ 378 ],
   alphaCSR[ 172 ][ 379 ],
   alphaCSR[ 172 ][ 380 ],
   alphaCSR[ 172 ][ 381 ],
   alphaCSR[ 172 ][ 382 ],
   alphaCSR[ 172 ][ 383 ],
   alphaCSR[ 173 ][ 0 ],
   alphaCSR[ 173 ][ 1 ],
   alphaCSR[ 173 ][ 2 ],
   alphaCSR[ 173 ][ 3 ],
   alphaCSR[ 173 ][ 4 ],
   alphaCSR[ 173 ][ 5 ],
   alphaCSR[ 173 ][ 6 ],
   alphaCSR[ 173 ][ 7 ],
   alphaCSR[ 173 ][ 8 ],
   alphaCSR[ 173 ][ 9 ],
   alphaCSR[ 173 ][ 10 ],
   alphaCSR[ 173 ][ 11 ],
   alphaCSR[ 173 ][ 12 ],
   alphaCSR[ 173 ][ 13 ],
   alphaCSR[ 173 ][ 14 ],
   alphaCSR[ 173 ][ 15 ],
   alphaCSR[ 173 ][ 16 ],
   alphaCSR[ 173 ][ 17 ],
   alphaCSR[ 173 ][ 18 ],
   alphaCSR[ 173 ][ 19 ],
   alphaCSR[ 173 ][ 20 ],
   alphaCSR[ 173 ][ 21 ],
   alphaCSR[ 173 ][ 22 ],
   alphaCSR[ 173 ][ 23 ],
   alphaCSR[ 173 ][ 24 ],
   alphaCSR[ 173 ][ 25 ],
   alphaCSR[ 173 ][ 26 ],
   alphaCSR[ 173 ][ 27 ],
   alphaCSR[ 173 ][ 28 ],
   alphaCSR[ 173 ][ 29 ],
   alphaCSR[ 173 ][ 30 ],
   alphaCSR[ 173 ][ 31 ],
   alphaCSR[ 173 ][ 32 ],
   alphaCSR[ 173 ][ 33 ],
   alphaCSR[ 173 ][ 34 ],
   alphaCSR[ 173 ][ 35 ],
   alphaCSR[ 173 ][ 36 ],
   alphaCSR[ 173 ][ 37 ],
   alphaCSR[ 173 ][ 38 ],
   alphaCSR[ 173 ][ 39 ],
   alphaCSR[ 173 ][ 40 ],
   alphaCSR[ 173 ][ 41 ],
   alphaCSR[ 173 ][ 42 ],
   alphaCSR[ 173 ][ 43 ],
   alphaCSR[ 173 ][ 44 ],
   alphaCSR[ 173 ][ 45 ],
   alphaCSR[ 173 ][ 46 ],
   alphaCSR[ 173 ][ 47 ],
   alphaCSR[ 173 ][ 48 ],
   alphaCSR[ 173 ][ 49 ],
   alphaCSR[ 173 ][ 50 ],
   alphaCSR[ 173 ][ 51 ],
   alphaCSR[ 173 ][ 52 ],
   alphaCSR[ 173 ][ 53 ],
   alphaCSR[ 173 ][ 54 ],
   alphaCSR[ 173 ][ 55 ],
   alphaCSR[ 173 ][ 56 ],
   alphaCSR[ 173 ][ 57 ],
   alphaCSR[ 173 ][ 58 ],
   alphaCSR[ 173 ][ 59 ],
   alphaCSR[ 173 ][ 60 ],
   alphaCSR[ 173 ][ 61 ],
   alphaCSR[ 173 ][ 62 ],
   alphaCSR[ 173 ][ 63 ],
   alphaCSR[ 173 ][ 64 ],
   alphaCSR[ 173 ][ 65 ],
   alphaCSR[ 173 ][ 66 ],
   alphaCSR[ 173 ][ 67 ],
   alphaCSR[ 173 ][ 68 ],
   alphaCSR[ 173 ][ 69 ],
   alphaCSR[ 173 ][ 70 ],
   alphaCSR[ 173 ][ 71 ],
   alphaCSR[ 173 ][ 72 ],
   alphaCSR[ 173 ][ 73 ],
   alphaCSR[ 173 ][ 74 ],
   alphaCSR[ 173 ][ 75 ],
   alphaCSR[ 173 ][ 76 ],
   alphaCSR[ 173 ][ 77 ],
   alphaCSR[ 173 ][ 78 ],
   alphaCSR[ 173 ][ 79 ],
   alphaCSR[ 173 ][ 80 ],
   alphaCSR[ 173 ][ 81 ],
   alphaCSR[ 173 ][ 82 ],
   alphaCSR[ 173 ][ 83 ],
   alphaCSR[ 173 ][ 84 ],
   alphaCSR[ 173 ][ 85 ],
   alphaCSR[ 173 ][ 86 ],
   alphaCSR[ 173 ][ 87 ],
   alphaCSR[ 173 ][ 88 ],
   alphaCSR[ 173 ][ 89 ],
   alphaCSR[ 173 ][ 90 ],
   alphaCSR[ 173 ][ 91 ],
   alphaCSR[ 173 ][ 92 ],
   alphaCSR[ 173 ][ 93 ],
   alphaCSR[ 173 ][ 94 ],
   alphaCSR[ 173 ][ 95 ],
   alphaCSR[ 173 ][ 96 ],
   alphaCSR[ 173 ][ 97 ],
   alphaCSR[ 173 ][ 98 ],
   alphaCSR[ 173 ][ 99 ],
   alphaCSR[ 173 ][ 100 ],
   alphaCSR[ 173 ][ 101 ],
   alphaCSR[ 173 ][ 102 ],
   alphaCSR[ 173 ][ 103 ],
   alphaCSR[ 173 ][ 104 ],
   alphaCSR[ 173 ][ 105 ],
   alphaCSR[ 173 ][ 106 ],
   alphaCSR[ 173 ][ 107 ],
   alphaCSR[ 173 ][ 108 ],
   alphaCSR[ 173 ][ 109 ],
   alphaCSR[ 173 ][ 110 ],
   alphaCSR[ 173 ][ 111 ],
   alphaCSR[ 173 ][ 112 ],
   alphaCSR[ 173 ][ 113 ],
   alphaCSR[ 173 ][ 114 ],
   alphaCSR[ 173 ][ 115 ],
   alphaCSR[ 173 ][ 116 ],
   alphaCSR[ 173 ][ 117 ],
   alphaCSR[ 173 ][ 118 ],
   alphaCSR[ 173 ][ 119 ],
   alphaCSR[ 173 ][ 120 ],
   alphaCSR[ 173 ][ 121 ],
   alphaCSR[ 173 ][ 122 ],
   alphaCSR[ 173 ][ 123 ],
   alphaCSR[ 173 ][ 124 ],
   alphaCSR[ 173 ][ 125 ],
   alphaCSR[ 173 ][ 126 ],
   alphaCSR[ 173 ][ 127 ],
   alphaCSR[ 173 ][ 128 ],
   alphaCSR[ 173 ][ 129 ],
   alphaCSR[ 173 ][ 130 ],
   alphaCSR[ 173 ][ 131 ],
   alphaCSR[ 173 ][ 132 ],
   alphaCSR[ 173 ][ 133 ],
   alphaCSR[ 173 ][ 134 ],
   alphaCSR[ 173 ][ 135 ],
   alphaCSR[ 173 ][ 136 ],
   alphaCSR[ 173 ][ 137 ],
   alphaCSR[ 173 ][ 138 ],
   alphaCSR[ 173 ][ 139 ],
   alphaCSR[ 173 ][ 140 ],
   alphaCSR[ 173 ][ 141 ],
   alphaCSR[ 173 ][ 142 ],
   alphaCSR[ 173 ][ 143 ],
   alphaCSR[ 173 ][ 144 ],
   alphaCSR[ 173 ][ 145 ],
   alphaCSR[ 173 ][ 146 ],
   alphaCSR[ 173 ][ 147 ],
   alphaCSR[ 173 ][ 148 ],
   alphaCSR[ 173 ][ 149 ],
   alphaCSR[ 173 ][ 150 ],
   alphaCSR[ 173 ][ 151 ],
   alphaCSR[ 173 ][ 152 ],
   alphaCSR[ 173 ][ 153 ],
   alphaCSR[ 173 ][ 154 ],
   alphaCSR[ 173 ][ 155 ],
   alphaCSR[ 173 ][ 156 ],
   alphaCSR[ 173 ][ 157 ],
   alphaCSR[ 173 ][ 158 ],
   alphaCSR[ 173 ][ 159 ],
   alphaCSR[ 173 ][ 160 ],
   alphaCSR[ 173 ][ 161 ],
   alphaCSR[ 173 ][ 162 ],
   alphaCSR[ 173 ][ 163 ],
   alphaCSR[ 173 ][ 164 ],
   alphaCSR[ 173 ][ 165 ],
   alphaCSR[ 173 ][ 166 ],
   alphaCSR[ 173 ][ 167 ],
   alphaCSR[ 173 ][ 168 ],
   alphaCSR[ 173 ][ 169 ],
   alphaCSR[ 173 ][ 170 ],
   alphaCSR[ 173 ][ 171 ],
   alphaCSR[ 173 ][ 172 ],
   alphaCSR[ 173 ][ 173 ],
   alphaCSR[ 173 ][ 174 ],
   alphaCSR[ 173 ][ 175 ],
   alphaCSR[ 173 ][ 176 ],
   alphaCSR[ 173 ][ 177 ],
   alphaCSR[ 173 ][ 178 ],
   alphaCSR[ 173 ][ 179 ],
   alphaCSR[ 173 ][ 180 ],
   alphaCSR[ 173 ][ 181 ],
   alphaCSR[ 173 ][ 182 ],
   alphaCSR[ 173 ][ 183 ],
   alphaCSR[ 173 ][ 184 ],
   alphaCSR[ 173 ][ 185 ],
   alphaCSR[ 173 ][ 186 ],
   alphaCSR[ 173 ][ 187 ],
   alphaCSR[ 173 ][ 188 ],
   alphaCSR[ 173 ][ 189 ],
   alphaCSR[ 173 ][ 190 ],
   alphaCSR[ 173 ][ 191 ],
   alphaCSR[ 173 ][ 192 ],
   alphaCSR[ 173 ][ 193 ],
   alphaCSR[ 173 ][ 194 ],
   alphaCSR[ 173 ][ 195 ],
   alphaCSR[ 173 ][ 196 ],
   alphaCSR[ 173 ][ 197 ],
   alphaCSR[ 173 ][ 198 ],
   alphaCSR[ 173 ][ 199 ],
   alphaCSR[ 173 ][ 200 ],
   alphaCSR[ 173 ][ 201 ],
   alphaCSR[ 173 ][ 202 ],
   alphaCSR[ 173 ][ 203 ],
   alphaCSR[ 173 ][ 204 ],
   alphaCSR[ 173 ][ 205 ],
   alphaCSR[ 173 ][ 206 ],
   alphaCSR[ 173 ][ 207 ],
   alphaCSR[ 173 ][ 208 ],
   alphaCSR[ 173 ][ 209 ],
   alphaCSR[ 173 ][ 210 ],
   alphaCSR[ 173 ][ 211 ],
   alphaCSR[ 173 ][ 212 ],
   alphaCSR[ 173 ][ 213 ],
   alphaCSR[ 173 ][ 214 ],
   alphaCSR[ 173 ][ 215 ],
   alphaCSR[ 173 ][ 216 ],
   alphaCSR[ 173 ][ 217 ],
   alphaCSR[ 173 ][ 218 ],
   alphaCSR[ 173 ][ 219 ],
   alphaCSR[ 173 ][ 220 ],
   alphaCSR[ 173 ][ 221 ],
   alphaCSR[ 173 ][ 222 ],
   alphaCSR[ 173 ][ 223 ],
   alphaCSR[ 173 ][ 224 ],
   alphaCSR[ 173 ][ 225 ],
   alphaCSR[ 173 ][ 226 ],
   alphaCSR[ 173 ][ 227 ],
   alphaCSR[ 173 ][ 228 ],
   alphaCSR[ 173 ][ 229 ],
   alphaCSR[ 173 ][ 230 ],
   alphaCSR[ 173 ][ 231 ],
   alphaCSR[ 173 ][ 232 ],
   alphaCSR[ 173 ][ 233 ],
   alphaCSR[ 173 ][ 234 ],
   alphaCSR[ 173 ][ 235 ],
   alphaCSR[ 173 ][ 236 ],
   alphaCSR[ 173 ][ 237 ],
   alphaCSR[ 173 ][ 238 ],
   alphaCSR[ 173 ][ 239 ],
   alphaCSR[ 173 ][ 240 ],
   alphaCSR[ 173 ][ 241 ],
   alphaCSR[ 173 ][ 242 ],
   alphaCSR[ 173 ][ 243 ],
   alphaCSR[ 173 ][ 244 ],
   alphaCSR[ 173 ][ 245 ],
   alphaCSR[ 173 ][ 246 ],
   alphaCSR[ 173 ][ 247 ],
   alphaCSR[ 173 ][ 248 ],
   alphaCSR[ 173 ][ 249 ],
   alphaCSR[ 173 ][ 250 ],
   alphaCSR[ 173 ][ 251 ],
   alphaCSR[ 173 ][ 252 ],
   alphaCSR[ 173 ][ 253 ],
   alphaCSR[ 173 ][ 254 ],
   alphaCSR[ 173 ][ 255 ],
   alphaCSR[ 173 ][ 256 ],
   alphaCSR[ 173 ][ 257 ],
   alphaCSR[ 173 ][ 258 ],
   alphaCSR[ 173 ][ 259 ],
   alphaCSR[ 173 ][ 260 ],
   alphaCSR[ 173 ][ 261 ],
   alphaCSR[ 173 ][ 262 ],
   alphaCSR[ 173 ][ 263 ],
   alphaCSR[ 173 ][ 264 ],
   alphaCSR[ 173 ][ 265 ],
   alphaCSR[ 173 ][ 266 ],
   alphaCSR[ 173 ][ 267 ],
   alphaCSR[ 173 ][ 268 ],
   alphaCSR[ 173 ][ 269 ],
   alphaCSR[ 173 ][ 270 ],
   alphaCSR[ 173 ][ 271 ],
   alphaCSR[ 173 ][ 272 ],
   alphaCSR[ 173 ][ 273 ],
   alphaCSR[ 173 ][ 274 ],
   alphaCSR[ 173 ][ 275 ],
   alphaCSR[ 173 ][ 276 ],
   alphaCSR[ 173 ][ 277 ],
   alphaCSR[ 173 ][ 278 ],
   alphaCSR[ 173 ][ 279 ],
   alphaCSR[ 173 ][ 280 ],
   alphaCSR[ 173 ][ 281 ],
   alphaCSR[ 173 ][ 282 ],
   alphaCSR[ 173 ][ 283 ],
   alphaCSR[ 173 ][ 284 ],
   alphaCSR[ 173 ][ 285 ],
   alphaCSR[ 173 ][ 286 ],
   alphaCSR[ 173 ][ 287 ],
   alphaCSR[ 173 ][ 288 ],
   alphaCSR[ 173 ][ 289 ],
   alphaCSR[ 173 ][ 290 ],
   alphaCSR[ 173 ][ 291 ],
   alphaCSR[ 173 ][ 292 ],
   alphaCSR[ 173 ][ 293 ],
   alphaCSR[ 173 ][ 294 ],
   alphaCSR[ 173 ][ 295 ],
   alphaCSR[ 173 ][ 296 ],
   alphaCSR[ 173 ][ 297 ],
   alphaCSR[ 173 ][ 298 ],
   alphaCSR[ 173 ][ 299 ],
   alphaCSR[ 173 ][ 300 ],
   alphaCSR[ 173 ][ 301 ],
   alphaCSR[ 173 ][ 302 ],
   alphaCSR[ 173 ][ 303 ],
   alphaCSR[ 173 ][ 304 ],
   alphaCSR[ 173 ][ 305 ],
   alphaCSR[ 173 ][ 306 ],
   alphaCSR[ 173 ][ 307 ],
   alphaCSR[ 173 ][ 308 ],
   alphaCSR[ 173 ][ 309 ],
   alphaCSR[ 173 ][ 310 ],
   alphaCSR[ 173 ][ 311 ],
   alphaCSR[ 173 ][ 312 ],
   alphaCSR[ 173 ][ 313 ],
   alphaCSR[ 173 ][ 314 ],
   alphaCSR[ 173 ][ 315 ],
   alphaCSR[ 173 ][ 316 ],
   alphaCSR[ 173 ][ 317 ],
   alphaCSR[ 173 ][ 318 ],
   alphaCSR[ 173 ][ 319 ],
   alphaCSR[ 173 ][ 320 ],
   alphaCSR[ 173 ][ 321 ],
   alphaCSR[ 173 ][ 322 ],
   alphaCSR[ 173 ][ 323 ],
   alphaCSR[ 173 ][ 324 ],
   alphaCSR[ 173 ][ 325 ],
   alphaCSR[ 173 ][ 326 ],
   alphaCSR[ 173 ][ 327 ],
   alphaCSR[ 173 ][ 328 ],
   alphaCSR[ 173 ][ 329 ],
   alphaCSR[ 173 ][ 330 ],
   alphaCSR[ 173 ][ 331 ],
   alphaCSR[ 173 ][ 332 ],
   alphaCSR[ 173 ][ 333 ],
   alphaCSR[ 173 ][ 334 ],
   alphaCSR[ 173 ][ 335 ],
   alphaCSR[ 173 ][ 336 ],
   alphaCSR[ 173 ][ 337 ],
   alphaCSR[ 173 ][ 338 ],
   alphaCSR[ 173 ][ 339 ],
   alphaCSR[ 173 ][ 340 ],
   alphaCSR[ 173 ][ 341 ],
   alphaCSR[ 173 ][ 342 ],
   alphaCSR[ 173 ][ 343 ],
   alphaCSR[ 173 ][ 344 ],
   alphaCSR[ 173 ][ 345 ],
   alphaCSR[ 173 ][ 346 ],
   alphaCSR[ 173 ][ 347 ],
   alphaCSR[ 173 ][ 348 ],
   alphaCSR[ 173 ][ 349 ],
   alphaCSR[ 173 ][ 350 ],
   alphaCSR[ 173 ][ 351 ],
   alphaCSR[ 173 ][ 352 ],
   alphaCSR[ 173 ][ 353 ],
   alphaCSR[ 173 ][ 354 ],
   alphaCSR[ 173 ][ 355 ],
   alphaCSR[ 173 ][ 356 ],
   alphaCSR[ 173 ][ 357 ],
   alphaCSR[ 173 ][ 358 ],
   alphaCSR[ 173 ][ 359 ],
   alphaCSR[ 173 ][ 360 ],
   alphaCSR[ 173 ][ 361 ],
   alphaCSR[ 173 ][ 362 ],
   alphaCSR[ 173 ][ 363 ],
   alphaCSR[ 173 ][ 364 ],
   alphaCSR[ 173 ][ 365 ],
   alphaCSR[ 173 ][ 366 ],
   alphaCSR[ 173 ][ 367 ],
   alphaCSR[ 173 ][ 368 ],
   alphaCSR[ 173 ][ 369 ],
   alphaCSR[ 173 ][ 370 ],
   alphaCSR[ 173 ][ 371 ],
   alphaCSR[ 173 ][ 372 ],
   alphaCSR[ 173 ][ 373 ],
   alphaCSR[ 173 ][ 374 ],
   alphaCSR[ 173 ][ 375 ],
   alphaCSR[ 173 ][ 376 ],
   alphaCSR[ 173 ][ 377 ],
   alphaCSR[ 173 ][ 378 ],
   alphaCSR[ 173 ][ 379 ],
   alphaCSR[ 173 ][ 380 ],
   alphaCSR[ 173 ][ 381 ],
   alphaCSR[ 173 ][ 382 ],
   alphaCSR[ 173 ][ 383 ],
   alphaCSR[ 174 ][ 0 ],
   alphaCSR[ 174 ][ 1 ],
   alphaCSR[ 174 ][ 2 ],
   alphaCSR[ 174 ][ 3 ],
   alphaCSR[ 174 ][ 4 ],
   alphaCSR[ 174 ][ 5 ],
   alphaCSR[ 174 ][ 6 ],
   alphaCSR[ 174 ][ 7 ],
   alphaCSR[ 174 ][ 8 ],
   alphaCSR[ 174 ][ 9 ],
   alphaCSR[ 174 ][ 10 ],
   alphaCSR[ 174 ][ 11 ],
   alphaCSR[ 174 ][ 12 ],
   alphaCSR[ 174 ][ 13 ],
   alphaCSR[ 174 ][ 14 ],
   alphaCSR[ 174 ][ 15 ],
   alphaCSR[ 174 ][ 16 ],
   alphaCSR[ 174 ][ 17 ],
   alphaCSR[ 174 ][ 18 ],
   alphaCSR[ 174 ][ 19 ],
   alphaCSR[ 174 ][ 20 ],
   alphaCSR[ 174 ][ 21 ],
   alphaCSR[ 174 ][ 22 ],
   alphaCSR[ 174 ][ 23 ],
   alphaCSR[ 174 ][ 24 ],
   alphaCSR[ 174 ][ 25 ],
   alphaCSR[ 174 ][ 26 ],
   alphaCSR[ 174 ][ 27 ],
   alphaCSR[ 174 ][ 28 ],
   alphaCSR[ 174 ][ 29 ],
   alphaCSR[ 174 ][ 30 ],
   alphaCSR[ 174 ][ 31 ],
   alphaCSR[ 174 ][ 32 ],
   alphaCSR[ 174 ][ 33 ],
   alphaCSR[ 174 ][ 34 ],
   alphaCSR[ 174 ][ 35 ],
   alphaCSR[ 174 ][ 36 ],
   alphaCSR[ 174 ][ 37 ],
   alphaCSR[ 174 ][ 38 ],
   alphaCSR[ 174 ][ 39 ],
   alphaCSR[ 174 ][ 40 ],
   alphaCSR[ 174 ][ 41 ],
   alphaCSR[ 174 ][ 42 ],
   alphaCSR[ 174 ][ 43 ],
   alphaCSR[ 174 ][ 44 ],
   alphaCSR[ 174 ][ 45 ],
   alphaCSR[ 174 ][ 46 ],
   alphaCSR[ 174 ][ 47 ],
   alphaCSR[ 174 ][ 48 ],
   alphaCSR[ 174 ][ 49 ],
   alphaCSR[ 174 ][ 50 ],
   alphaCSR[ 174 ][ 51 ],
   alphaCSR[ 174 ][ 52 ],
   alphaCSR[ 174 ][ 53 ],
   alphaCSR[ 174 ][ 54 ],
   alphaCSR[ 174 ][ 55 ],
   alphaCSR[ 174 ][ 56 ],
   alphaCSR[ 174 ][ 57 ],
   alphaCSR[ 174 ][ 58 ],
   alphaCSR[ 174 ][ 59 ],
   alphaCSR[ 174 ][ 60 ],
   alphaCSR[ 174 ][ 61 ],
   alphaCSR[ 174 ][ 62 ],
   alphaCSR[ 174 ][ 63 ],
   alphaCSR[ 174 ][ 64 ],
   alphaCSR[ 174 ][ 65 ],
   alphaCSR[ 174 ][ 66 ],
   alphaCSR[ 174 ][ 67 ],
   alphaCSR[ 174 ][ 68 ],
   alphaCSR[ 174 ][ 69 ],
   alphaCSR[ 174 ][ 70 ],
   alphaCSR[ 174 ][ 71 ],
   alphaCSR[ 174 ][ 72 ],
   alphaCSR[ 174 ][ 73 ],
   alphaCSR[ 174 ][ 74 ],
   alphaCSR[ 174 ][ 75 ],
   alphaCSR[ 174 ][ 76 ],
   alphaCSR[ 174 ][ 77 ],
   alphaCSR[ 174 ][ 78 ],
   alphaCSR[ 174 ][ 79 ],
   alphaCSR[ 174 ][ 80 ],
   alphaCSR[ 174 ][ 81 ],
   alphaCSR[ 174 ][ 82 ],
   alphaCSR[ 174 ][ 83 ],
   alphaCSR[ 174 ][ 84 ],
   alphaCSR[ 174 ][ 85 ],
   alphaCSR[ 174 ][ 86 ],
   alphaCSR[ 174 ][ 87 ],
   alphaCSR[ 174 ][ 88 ],
   alphaCSR[ 174 ][ 89 ],
   alphaCSR[ 174 ][ 90 ],
   alphaCSR[ 174 ][ 91 ],
   alphaCSR[ 174 ][ 92 ],
   alphaCSR[ 174 ][ 93 ],
   alphaCSR[ 174 ][ 94 ],
   alphaCSR[ 174 ][ 95 ],
   alphaCSR[ 174 ][ 96 ],
   alphaCSR[ 174 ][ 97 ],
   alphaCSR[ 174 ][ 98 ],
   alphaCSR[ 174 ][ 99 ],
   alphaCSR[ 174 ][ 100 ],
   alphaCSR[ 174 ][ 101 ],
   alphaCSR[ 174 ][ 102 ],
   alphaCSR[ 174 ][ 103 ],
   alphaCSR[ 174 ][ 104 ],
   alphaCSR[ 174 ][ 105 ],
   alphaCSR[ 174 ][ 106 ],
   alphaCSR[ 174 ][ 107 ],
   alphaCSR[ 174 ][ 108 ],
   alphaCSR[ 174 ][ 109 ],
   alphaCSR[ 174 ][ 110 ],
   alphaCSR[ 174 ][ 111 ],
   alphaCSR[ 174 ][ 112 ],
   alphaCSR[ 174 ][ 113 ],
   alphaCSR[ 174 ][ 114 ],
   alphaCSR[ 174 ][ 115 ],
   alphaCSR[ 174 ][ 116 ],
   alphaCSR[ 174 ][ 117 ],
   alphaCSR[ 174 ][ 118 ],
   alphaCSR[ 174 ][ 119 ],
   alphaCSR[ 174 ][ 120 ],
   alphaCSR[ 174 ][ 121 ],
   alphaCSR[ 174 ][ 122 ],
   alphaCSR[ 174 ][ 123 ],
   alphaCSR[ 174 ][ 124 ],
   alphaCSR[ 174 ][ 125 ],
   alphaCSR[ 174 ][ 126 ],
   alphaCSR[ 174 ][ 127 ],
   alphaCSR[ 174 ][ 128 ],
   alphaCSR[ 174 ][ 129 ],
   alphaCSR[ 174 ][ 130 ],
   alphaCSR[ 174 ][ 131 ],
   alphaCSR[ 174 ][ 132 ],
   alphaCSR[ 174 ][ 133 ],
   alphaCSR[ 174 ][ 134 ],
   alphaCSR[ 174 ][ 135 ],
   alphaCSR[ 174 ][ 136 ],
   alphaCSR[ 174 ][ 137 ],
   alphaCSR[ 174 ][ 138 ],
   alphaCSR[ 174 ][ 139 ],
   alphaCSR[ 174 ][ 140 ],
   alphaCSR[ 174 ][ 141 ],
   alphaCSR[ 174 ][ 142 ],
   alphaCSR[ 174 ][ 143 ],
   alphaCSR[ 174 ][ 144 ],
   alphaCSR[ 174 ][ 145 ],
   alphaCSR[ 174 ][ 146 ],
   alphaCSR[ 174 ][ 147 ],
   alphaCSR[ 174 ][ 148 ],
   alphaCSR[ 174 ][ 149 ],
   alphaCSR[ 174 ][ 150 ],
   alphaCSR[ 174 ][ 151 ],
   alphaCSR[ 174 ][ 152 ],
   alphaCSR[ 174 ][ 153 ],
   alphaCSR[ 174 ][ 154 ],
   alphaCSR[ 174 ][ 155 ],
   alphaCSR[ 174 ][ 156 ],
   alphaCSR[ 174 ][ 157 ],
   alphaCSR[ 174 ][ 158 ],
   alphaCSR[ 174 ][ 159 ],
   alphaCSR[ 174 ][ 160 ],
   alphaCSR[ 174 ][ 161 ],
   alphaCSR[ 174 ][ 162 ],
   alphaCSR[ 174 ][ 163 ],
   alphaCSR[ 174 ][ 164 ],
   alphaCSR[ 174 ][ 165 ],
   alphaCSR[ 174 ][ 166 ],
   alphaCSR[ 174 ][ 167 ],
   alphaCSR[ 174 ][ 168 ],
   alphaCSR[ 174 ][ 169 ],
   alphaCSR[ 174 ][ 170 ],
   alphaCSR[ 174 ][ 171 ],
   alphaCSR[ 174 ][ 172 ],
   alphaCSR[ 174 ][ 173 ],
   alphaCSR[ 174 ][ 174 ],
   alphaCSR[ 174 ][ 175 ],
   alphaCSR[ 174 ][ 176 ],
   alphaCSR[ 174 ][ 177 ],
   alphaCSR[ 174 ][ 178 ],
   alphaCSR[ 174 ][ 179 ],
   alphaCSR[ 174 ][ 180 ],
   alphaCSR[ 174 ][ 181 ],
   alphaCSR[ 174 ][ 182 ],
   alphaCSR[ 174 ][ 183 ],
   alphaCSR[ 174 ][ 184 ],
   alphaCSR[ 174 ][ 185 ],
   alphaCSR[ 174 ][ 186 ],
   alphaCSR[ 174 ][ 187 ],
   alphaCSR[ 174 ][ 188 ],
   alphaCSR[ 174 ][ 189 ],
   alphaCSR[ 174 ][ 190 ],
   alphaCSR[ 174 ][ 191 ],
   alphaCSR[ 174 ][ 192 ],
   alphaCSR[ 174 ][ 193 ],
   alphaCSR[ 174 ][ 194 ],
   alphaCSR[ 174 ][ 195 ],
   alphaCSR[ 174 ][ 196 ],
   alphaCSR[ 174 ][ 197 ],
   alphaCSR[ 174 ][ 198 ],
   alphaCSR[ 174 ][ 199 ],
   alphaCSR[ 174 ][ 200 ],
   alphaCSR[ 174 ][ 201 ],
   alphaCSR[ 174 ][ 202 ],
   alphaCSR[ 174 ][ 203 ],
   alphaCSR[ 174 ][ 204 ],
   alphaCSR[ 174 ][ 205 ],
   alphaCSR[ 174 ][ 206 ],
   alphaCSR[ 174 ][ 207 ],
   alphaCSR[ 174 ][ 208 ],
   alphaCSR[ 174 ][ 209 ],
   alphaCSR[ 174 ][ 210 ],
   alphaCSR[ 174 ][ 211 ],
   alphaCSR[ 174 ][ 212 ],
   alphaCSR[ 174 ][ 213 ],
   alphaCSR[ 174 ][ 214 ],
   alphaCSR[ 174 ][ 215 ],
   alphaCSR[ 174 ][ 216 ],
   alphaCSR[ 174 ][ 217 ],
   alphaCSR[ 174 ][ 218 ],
   alphaCSR[ 174 ][ 219 ],
   alphaCSR[ 174 ][ 220 ],
   alphaCSR[ 174 ][ 221 ],
   alphaCSR[ 174 ][ 222 ],
   alphaCSR[ 174 ][ 223 ],
   alphaCSR[ 174 ][ 224 ],
   alphaCSR[ 174 ][ 225 ],
   alphaCSR[ 174 ][ 226 ],
   alphaCSR[ 174 ][ 227 ],
   alphaCSR[ 174 ][ 228 ],
   alphaCSR[ 174 ][ 229 ],
   alphaCSR[ 174 ][ 230 ],
   alphaCSR[ 174 ][ 231 ],
   alphaCSR[ 174 ][ 232 ],
   alphaCSR[ 174 ][ 233 ],
   alphaCSR[ 174 ][ 234 ],
   alphaCSR[ 174 ][ 235 ],
   alphaCSR[ 174 ][ 236 ],
   alphaCSR[ 174 ][ 237 ],
   alphaCSR[ 174 ][ 238 ],
   alphaCSR[ 174 ][ 239 ],
   alphaCSR[ 174 ][ 240 ],
   alphaCSR[ 174 ][ 241 ],
   alphaCSR[ 174 ][ 242 ],
   alphaCSR[ 174 ][ 243 ],
   alphaCSR[ 174 ][ 244 ],
   alphaCSR[ 174 ][ 245 ],
   alphaCSR[ 174 ][ 246 ],
   alphaCSR[ 174 ][ 247 ],
   alphaCSR[ 174 ][ 248 ],
   alphaCSR[ 174 ][ 249 ],
   alphaCSR[ 174 ][ 250 ],
   alphaCSR[ 174 ][ 251 ],
   alphaCSR[ 174 ][ 252 ],
   alphaCSR[ 174 ][ 253 ],
   alphaCSR[ 174 ][ 254 ],
   alphaCSR[ 174 ][ 255 ],
   alphaCSR[ 174 ][ 256 ],
   alphaCSR[ 174 ][ 257 ],
   alphaCSR[ 174 ][ 258 ],
   alphaCSR[ 174 ][ 259 ],
   alphaCSR[ 174 ][ 260 ],
   alphaCSR[ 174 ][ 261 ],
   alphaCSR[ 174 ][ 262 ],
   alphaCSR[ 174 ][ 263 ],
   alphaCSR[ 174 ][ 264 ],
   alphaCSR[ 174 ][ 265 ],
   alphaCSR[ 174 ][ 266 ],
   alphaCSR[ 174 ][ 267 ],
   alphaCSR[ 174 ][ 268 ],
   alphaCSR[ 174 ][ 269 ],
   alphaCSR[ 174 ][ 270 ],
   alphaCSR[ 174 ][ 271 ],
   alphaCSR[ 174 ][ 272 ],
   alphaCSR[ 174 ][ 273 ],
   alphaCSR[ 174 ][ 274 ],
   alphaCSR[ 174 ][ 275 ],
   alphaCSR[ 174 ][ 276 ],
   alphaCSR[ 174 ][ 277 ],
   alphaCSR[ 174 ][ 278 ],
   alphaCSR[ 174 ][ 279 ],
   alphaCSR[ 174 ][ 280 ],
   alphaCSR[ 174 ][ 281 ],
   alphaCSR[ 174 ][ 282 ],
   alphaCSR[ 174 ][ 283 ],
   alphaCSR[ 174 ][ 284 ],
   alphaCSR[ 174 ][ 285 ],
   alphaCSR[ 174 ][ 286 ],
   alphaCSR[ 174 ][ 287 ],
   alphaCSR[ 174 ][ 288 ],
   alphaCSR[ 174 ][ 289 ],
   alphaCSR[ 174 ][ 290 ],
   alphaCSR[ 174 ][ 291 ],
   alphaCSR[ 174 ][ 292 ],
   alphaCSR[ 174 ][ 293 ],
   alphaCSR[ 174 ][ 294 ],
   alphaCSR[ 174 ][ 295 ],
   alphaCSR[ 174 ][ 296 ],
   alphaCSR[ 174 ][ 297 ],
   alphaCSR[ 174 ][ 298 ],
   alphaCSR[ 174 ][ 299 ],
   alphaCSR[ 174 ][ 300 ],
   alphaCSR[ 174 ][ 301 ],
   alphaCSR[ 174 ][ 302 ],
   alphaCSR[ 174 ][ 303 ],
   alphaCSR[ 174 ][ 304 ],
   alphaCSR[ 174 ][ 305 ],
   alphaCSR[ 174 ][ 306 ],
   alphaCSR[ 174 ][ 307 ],
   alphaCSR[ 174 ][ 308 ],
   alphaCSR[ 174 ][ 309 ],
   alphaCSR[ 174 ][ 310 ],
   alphaCSR[ 174 ][ 311 ],
   alphaCSR[ 174 ][ 312 ],
   alphaCSR[ 174 ][ 313 ],
   alphaCSR[ 174 ][ 314 ],
   alphaCSR[ 174 ][ 315 ],
   alphaCSR[ 174 ][ 316 ],
   alphaCSR[ 174 ][ 317 ],
   alphaCSR[ 174 ][ 318 ],
   alphaCSR[ 174 ][ 319 ],
   alphaCSR[ 174 ][ 320 ],
   alphaCSR[ 174 ][ 321 ],
   alphaCSR[ 174 ][ 322 ],
   alphaCSR[ 174 ][ 323 ],
   alphaCSR[ 174 ][ 324 ],
   alphaCSR[ 174 ][ 325 ],
   alphaCSR[ 174 ][ 326 ],
   alphaCSR[ 174 ][ 327 ],
   alphaCSR[ 174 ][ 328 ],
   alphaCSR[ 174 ][ 329 ],
   alphaCSR[ 174 ][ 330 ],
   alphaCSR[ 174 ][ 331 ],
   alphaCSR[ 174 ][ 332 ],
   alphaCSR[ 174 ][ 333 ],
   alphaCSR[ 174 ][ 334 ],
   alphaCSR[ 174 ][ 335 ],
   alphaCSR[ 174 ][ 336 ],
   alphaCSR[ 174 ][ 337 ],
   alphaCSR[ 174 ][ 338 ],
   alphaCSR[ 174 ][ 339 ],
   alphaCSR[ 174 ][ 340 ],
   alphaCSR[ 174 ][ 341 ],
   alphaCSR[ 174 ][ 342 ],
   alphaCSR[ 174 ][ 343 ],
   alphaCSR[ 174 ][ 344 ],
   alphaCSR[ 174 ][ 345 ],
   alphaCSR[ 174 ][ 346 ],
   alphaCSR[ 174 ][ 347 ],
   alphaCSR[ 174 ][ 348 ],
   alphaCSR[ 174 ][ 349 ],
   alphaCSR[ 174 ][ 350 ],
   alphaCSR[ 174 ][ 351 ],
   alphaCSR[ 174 ][ 352 ],
   alphaCSR[ 174 ][ 353 ],
   alphaCSR[ 174 ][ 354 ],
   alphaCSR[ 174 ][ 355 ],
   alphaCSR[ 174 ][ 356 ],
   alphaCSR[ 174 ][ 357 ],
   alphaCSR[ 174 ][ 358 ],
   alphaCSR[ 174 ][ 359 ],
   alphaCSR[ 174 ][ 360 ],
   alphaCSR[ 174 ][ 361 ],
   alphaCSR[ 174 ][ 362 ],
   alphaCSR[ 174 ][ 363 ],
   alphaCSR[ 174 ][ 364 ],
   alphaCSR[ 174 ][ 365 ],
   alphaCSR[ 174 ][ 366 ],
   alphaCSR[ 174 ][ 367 ],
   alphaCSR[ 174 ][ 368 ],
   alphaCSR[ 174 ][ 369 ],
   alphaCSR[ 174 ][ 370 ],
   alphaCSR[ 174 ][ 371 ],
   alphaCSR[ 174 ][ 372 ],
   alphaCSR[ 174 ][ 373 ],
   alphaCSR[ 174 ][ 374 ],
   alphaCSR[ 174 ][ 375 ],
   alphaCSR[ 174 ][ 376 ],
   alphaCSR[ 174 ][ 377 ],
   alphaCSR[ 174 ][ 378 ],
   alphaCSR[ 174 ][ 379 ],
   alphaCSR[ 174 ][ 380 ],
   alphaCSR[ 174 ][ 381 ],
   alphaCSR[ 174 ][ 382 ],
   alphaCSR[ 174 ][ 383 ],
   alphaCSR[ 175 ][ 0 ],
   alphaCSR[ 175 ][ 1 ],
   alphaCSR[ 175 ][ 2 ],
   alphaCSR[ 175 ][ 3 ],
   alphaCSR[ 175 ][ 4 ],
   alphaCSR[ 175 ][ 5 ],
   alphaCSR[ 175 ][ 6 ],
   alphaCSR[ 175 ][ 7 ],
   alphaCSR[ 175 ][ 8 ],
   alphaCSR[ 175 ][ 9 ],
   alphaCSR[ 175 ][ 10 ],
   alphaCSR[ 175 ][ 11 ],
   alphaCSR[ 175 ][ 12 ],
   alphaCSR[ 175 ][ 13 ],
   alphaCSR[ 175 ][ 14 ],
   alphaCSR[ 175 ][ 15 ],
   alphaCSR[ 175 ][ 16 ],
   alphaCSR[ 175 ][ 17 ],
   alphaCSR[ 175 ][ 18 ],
   alphaCSR[ 175 ][ 19 ],
   alphaCSR[ 175 ][ 20 ],
   alphaCSR[ 175 ][ 21 ],
   alphaCSR[ 175 ][ 22 ],
   alphaCSR[ 175 ][ 23 ],
   alphaCSR[ 175 ][ 24 ],
   alphaCSR[ 175 ][ 25 ],
   alphaCSR[ 175 ][ 26 ],
   alphaCSR[ 175 ][ 27 ],
   alphaCSR[ 175 ][ 28 ],
   alphaCSR[ 175 ][ 29 ],
   alphaCSR[ 175 ][ 30 ],
   alphaCSR[ 175 ][ 31 ],
   alphaCSR[ 175 ][ 32 ],
   alphaCSR[ 175 ][ 33 ],
   alphaCSR[ 175 ][ 34 ],
   alphaCSR[ 175 ][ 35 ],
   alphaCSR[ 175 ][ 36 ],
   alphaCSR[ 175 ][ 37 ],
   alphaCSR[ 175 ][ 38 ],
   alphaCSR[ 175 ][ 39 ],
   alphaCSR[ 175 ][ 40 ],
   alphaCSR[ 175 ][ 41 ],
   alphaCSR[ 175 ][ 42 ],
   alphaCSR[ 175 ][ 43 ],
   alphaCSR[ 175 ][ 44 ],
   alphaCSR[ 175 ][ 45 ],
   alphaCSR[ 175 ][ 46 ],
   alphaCSR[ 175 ][ 47 ],
   alphaCSR[ 175 ][ 48 ],
   alphaCSR[ 175 ][ 49 ],
   alphaCSR[ 175 ][ 50 ],
   alphaCSR[ 175 ][ 51 ],
   alphaCSR[ 175 ][ 52 ],
   alphaCSR[ 175 ][ 53 ],
   alphaCSR[ 175 ][ 54 ],
   alphaCSR[ 175 ][ 55 ],
   alphaCSR[ 175 ][ 56 ],
   alphaCSR[ 175 ][ 57 ],
   alphaCSR[ 175 ][ 58 ],
   alphaCSR[ 175 ][ 59 ],
   alphaCSR[ 175 ][ 60 ],
   alphaCSR[ 175 ][ 61 ],
   alphaCSR[ 175 ][ 62 ],
   alphaCSR[ 175 ][ 63 ],
   alphaCSR[ 175 ][ 64 ],
   alphaCSR[ 175 ][ 65 ],
   alphaCSR[ 175 ][ 66 ],
   alphaCSR[ 175 ][ 67 ],
   alphaCSR[ 175 ][ 68 ],
   alphaCSR[ 175 ][ 69 ],
   alphaCSR[ 175 ][ 70 ],
   alphaCSR[ 175 ][ 71 ],
   alphaCSR[ 175 ][ 72 ],
   alphaCSR[ 175 ][ 73 ],
   alphaCSR[ 175 ][ 74 ],
   alphaCSR[ 175 ][ 75 ],
   alphaCSR[ 175 ][ 76 ],
   alphaCSR[ 175 ][ 77 ],
   alphaCSR[ 175 ][ 78 ],
   alphaCSR[ 175 ][ 79 ],
   alphaCSR[ 175 ][ 80 ],
   alphaCSR[ 175 ][ 81 ],
   alphaCSR[ 175 ][ 82 ],
   alphaCSR[ 175 ][ 83 ],
   alphaCSR[ 175 ][ 84 ],
   alphaCSR[ 175 ][ 85 ],
   alphaCSR[ 175 ][ 86 ],
   alphaCSR[ 175 ][ 87 ],
   alphaCSR[ 175 ][ 88 ],
   alphaCSR[ 175 ][ 89 ],
   alphaCSR[ 175 ][ 90 ],
   alphaCSR[ 175 ][ 91 ],
   alphaCSR[ 175 ][ 92 ],
   alphaCSR[ 175 ][ 93 ],
   alphaCSR[ 175 ][ 94 ],
   alphaCSR[ 175 ][ 95 ],
   alphaCSR[ 175 ][ 96 ],
   alphaCSR[ 175 ][ 97 ],
   alphaCSR[ 175 ][ 98 ],
   alphaCSR[ 175 ][ 99 ],
   alphaCSR[ 175 ][ 100 ],
   alphaCSR[ 175 ][ 101 ],
   alphaCSR[ 175 ][ 102 ],
   alphaCSR[ 175 ][ 103 ],
   alphaCSR[ 175 ][ 104 ],
   alphaCSR[ 175 ][ 105 ],
   alphaCSR[ 175 ][ 106 ],
   alphaCSR[ 175 ][ 107 ],
   alphaCSR[ 175 ][ 108 ],
   alphaCSR[ 175 ][ 109 ],
   alphaCSR[ 175 ][ 110 ],
   alphaCSR[ 175 ][ 111 ],
   alphaCSR[ 175 ][ 112 ],
   alphaCSR[ 175 ][ 113 ],
   alphaCSR[ 175 ][ 114 ],
   alphaCSR[ 175 ][ 115 ],
   alphaCSR[ 175 ][ 116 ],
   alphaCSR[ 175 ][ 117 ],
   alphaCSR[ 175 ][ 118 ],
   alphaCSR[ 175 ][ 119 ],
   alphaCSR[ 175 ][ 120 ],
   alphaCSR[ 175 ][ 121 ],
   alphaCSR[ 175 ][ 122 ],
   alphaCSR[ 175 ][ 123 ],
   alphaCSR[ 175 ][ 124 ],
   alphaCSR[ 175 ][ 125 ],
   alphaCSR[ 175 ][ 126 ],
   alphaCSR[ 175 ][ 127 ],
   alphaCSR[ 175 ][ 128 ],
   alphaCSR[ 175 ][ 129 ],
   alphaCSR[ 175 ][ 130 ],
   alphaCSR[ 175 ][ 131 ],
   alphaCSR[ 175 ][ 132 ],
   alphaCSR[ 175 ][ 133 ],
   alphaCSR[ 175 ][ 134 ],
   alphaCSR[ 175 ][ 135 ],
   alphaCSR[ 175 ][ 136 ],
   alphaCSR[ 175 ][ 137 ],
   alphaCSR[ 175 ][ 138 ],
   alphaCSR[ 175 ][ 139 ],
   alphaCSR[ 175 ][ 140 ],
   alphaCSR[ 175 ][ 141 ],
   alphaCSR[ 175 ][ 142 ],
   alphaCSR[ 175 ][ 143 ],
   alphaCSR[ 175 ][ 144 ],
   alphaCSR[ 175 ][ 145 ],
   alphaCSR[ 175 ][ 146 ],
   alphaCSR[ 175 ][ 147 ],
   alphaCSR[ 175 ][ 148 ],
   alphaCSR[ 175 ][ 149 ],
   alphaCSR[ 175 ][ 150 ],
   alphaCSR[ 175 ][ 151 ],
   alphaCSR[ 175 ][ 152 ],
   alphaCSR[ 175 ][ 153 ],
   alphaCSR[ 175 ][ 154 ],
   alphaCSR[ 175 ][ 155 ],
   alphaCSR[ 175 ][ 156 ],
   alphaCSR[ 175 ][ 157 ],
   alphaCSR[ 175 ][ 158 ],
   alphaCSR[ 175 ][ 159 ],
   alphaCSR[ 175 ][ 160 ],
   alphaCSR[ 175 ][ 161 ],
   alphaCSR[ 175 ][ 162 ],
   alphaCSR[ 175 ][ 163 ],
   alphaCSR[ 175 ][ 164 ],
   alphaCSR[ 175 ][ 165 ],
   alphaCSR[ 175 ][ 166 ],
   alphaCSR[ 175 ][ 167 ],
   alphaCSR[ 175 ][ 168 ],
   alphaCSR[ 175 ][ 169 ],
   alphaCSR[ 175 ][ 170 ],
   alphaCSR[ 175 ][ 171 ],
   alphaCSR[ 175 ][ 172 ],
   alphaCSR[ 175 ][ 173 ],
   alphaCSR[ 175 ][ 174 ],
   alphaCSR[ 175 ][ 175 ],
   alphaCSR[ 175 ][ 176 ],
   alphaCSR[ 175 ][ 177 ],
   alphaCSR[ 175 ][ 178 ],
   alphaCSR[ 175 ][ 179 ],
   alphaCSR[ 175 ][ 180 ],
   alphaCSR[ 175 ][ 181 ],
   alphaCSR[ 175 ][ 182 ],
   alphaCSR[ 175 ][ 183 ],
   alphaCSR[ 175 ][ 184 ],
   alphaCSR[ 175 ][ 185 ],
   alphaCSR[ 175 ][ 186 ],
   alphaCSR[ 175 ][ 187 ],
   alphaCSR[ 175 ][ 188 ],
   alphaCSR[ 175 ][ 189 ],
   alphaCSR[ 175 ][ 190 ],
   alphaCSR[ 175 ][ 191 ],
   alphaCSR[ 175 ][ 192 ],
   alphaCSR[ 175 ][ 193 ],
   alphaCSR[ 175 ][ 194 ],
   alphaCSR[ 175 ][ 195 ],
   alphaCSR[ 175 ][ 196 ],
   alphaCSR[ 175 ][ 197 ],
   alphaCSR[ 175 ][ 198 ],
   alphaCSR[ 175 ][ 199 ],
   alphaCSR[ 175 ][ 200 ],
   alphaCSR[ 175 ][ 201 ],
   alphaCSR[ 175 ][ 202 ],
   alphaCSR[ 175 ][ 203 ],
   alphaCSR[ 175 ][ 204 ],
   alphaCSR[ 175 ][ 205 ],
   alphaCSR[ 175 ][ 206 ],
   alphaCSR[ 175 ][ 207 ],
   alphaCSR[ 175 ][ 208 ],
   alphaCSR[ 175 ][ 209 ],
   alphaCSR[ 175 ][ 210 ],
   alphaCSR[ 175 ][ 211 ],
   alphaCSR[ 175 ][ 212 ],
   alphaCSR[ 175 ][ 213 ],
   alphaCSR[ 175 ][ 214 ],
   alphaCSR[ 175 ][ 215 ],
   alphaCSR[ 175 ][ 216 ],
   alphaCSR[ 175 ][ 217 ],
   alphaCSR[ 175 ][ 218 ],
   alphaCSR[ 175 ][ 219 ],
   alphaCSR[ 175 ][ 220 ],
   alphaCSR[ 175 ][ 221 ],
   alphaCSR[ 175 ][ 222 ],
   alphaCSR[ 175 ][ 223 ],
   alphaCSR[ 175 ][ 224 ],
   alphaCSR[ 175 ][ 225 ],
   alphaCSR[ 175 ][ 226 ],
   alphaCSR[ 175 ][ 227 ],
   alphaCSR[ 175 ][ 228 ],
   alphaCSR[ 175 ][ 229 ],
   alphaCSR[ 175 ][ 230 ],
   alphaCSR[ 175 ][ 231 ],
   alphaCSR[ 175 ][ 232 ],
   alphaCSR[ 175 ][ 233 ],
   alphaCSR[ 175 ][ 234 ],
   alphaCSR[ 175 ][ 235 ],
   alphaCSR[ 175 ][ 236 ],
   alphaCSR[ 175 ][ 237 ],
   alphaCSR[ 175 ][ 238 ],
   alphaCSR[ 175 ][ 239 ],
   alphaCSR[ 175 ][ 240 ],
   alphaCSR[ 175 ][ 241 ],
   alphaCSR[ 175 ][ 242 ],
   alphaCSR[ 175 ][ 243 ],
   alphaCSR[ 175 ][ 244 ],
   alphaCSR[ 175 ][ 245 ],
   alphaCSR[ 175 ][ 246 ],
   alphaCSR[ 175 ][ 247 ],
   alphaCSR[ 175 ][ 248 ],
   alphaCSR[ 175 ][ 249 ],
   alphaCSR[ 175 ][ 250 ],
   alphaCSR[ 175 ][ 251 ],
   alphaCSR[ 175 ][ 252 ],
   alphaCSR[ 175 ][ 253 ],
   alphaCSR[ 175 ][ 254 ],
   alphaCSR[ 175 ][ 255 ],
   alphaCSR[ 175 ][ 256 ],
   alphaCSR[ 175 ][ 257 ],
   alphaCSR[ 175 ][ 258 ],
   alphaCSR[ 175 ][ 259 ],
   alphaCSR[ 175 ][ 260 ],
   alphaCSR[ 175 ][ 261 ],
   alphaCSR[ 175 ][ 262 ],
   alphaCSR[ 175 ][ 263 ],
   alphaCSR[ 175 ][ 264 ],
   alphaCSR[ 175 ][ 265 ],
   alphaCSR[ 175 ][ 266 ],
   alphaCSR[ 175 ][ 267 ],
   alphaCSR[ 175 ][ 268 ],
   alphaCSR[ 175 ][ 269 ],
   alphaCSR[ 175 ][ 270 ],
   alphaCSR[ 175 ][ 271 ],
   alphaCSR[ 175 ][ 272 ],
   alphaCSR[ 175 ][ 273 ],
   alphaCSR[ 175 ][ 274 ],
   alphaCSR[ 175 ][ 275 ],
   alphaCSR[ 175 ][ 276 ],
   alphaCSR[ 175 ][ 277 ],
   alphaCSR[ 175 ][ 278 ],
   alphaCSR[ 175 ][ 279 ],
   alphaCSR[ 175 ][ 280 ],
   alphaCSR[ 175 ][ 281 ],
   alphaCSR[ 175 ][ 282 ],
   alphaCSR[ 175 ][ 283 ],
   alphaCSR[ 175 ][ 284 ],
   alphaCSR[ 175 ][ 285 ],
   alphaCSR[ 175 ][ 286 ],
   alphaCSR[ 175 ][ 287 ],
   alphaCSR[ 175 ][ 288 ],
   alphaCSR[ 175 ][ 289 ],
   alphaCSR[ 175 ][ 290 ],
   alphaCSR[ 175 ][ 291 ],
   alphaCSR[ 175 ][ 292 ],
   alphaCSR[ 175 ][ 293 ],
   alphaCSR[ 175 ][ 294 ],
   alphaCSR[ 175 ][ 295 ],
   alphaCSR[ 175 ][ 296 ],
   alphaCSR[ 175 ][ 297 ],
   alphaCSR[ 175 ][ 298 ],
   alphaCSR[ 175 ][ 299 ],
   alphaCSR[ 175 ][ 300 ],
   alphaCSR[ 175 ][ 301 ],
   alphaCSR[ 175 ][ 302 ],
   alphaCSR[ 175 ][ 303 ],
   alphaCSR[ 175 ][ 304 ],
   alphaCSR[ 175 ][ 305 ],
   alphaCSR[ 175 ][ 306 ],
   alphaCSR[ 175 ][ 307 ],
   alphaCSR[ 175 ][ 308 ],
   alphaCSR[ 175 ][ 309 ],
   alphaCSR[ 175 ][ 310 ],
   alphaCSR[ 175 ][ 311 ],
   alphaCSR[ 175 ][ 312 ],
   alphaCSR[ 175 ][ 313 ],
   alphaCSR[ 175 ][ 314 ],
   alphaCSR[ 175 ][ 315 ],
   alphaCSR[ 175 ][ 316 ],
   alphaCSR[ 175 ][ 317 ],
   alphaCSR[ 175 ][ 318 ],
   alphaCSR[ 175 ][ 319 ],
   alphaCSR[ 175 ][ 320 ],
   alphaCSR[ 175 ][ 321 ],
   alphaCSR[ 175 ][ 322 ],
   alphaCSR[ 175 ][ 323 ],
   alphaCSR[ 175 ][ 324 ],
   alphaCSR[ 175 ][ 325 ],
   alphaCSR[ 175 ][ 326 ],
   alphaCSR[ 175 ][ 327 ],
   alphaCSR[ 175 ][ 328 ],
   alphaCSR[ 175 ][ 329 ],
   alphaCSR[ 175 ][ 330 ],
   alphaCSR[ 175 ][ 331 ],
   alphaCSR[ 175 ][ 332 ],
   alphaCSR[ 175 ][ 333 ],
   alphaCSR[ 175 ][ 334 ],
   alphaCSR[ 175 ][ 335 ],
   alphaCSR[ 175 ][ 336 ],
   alphaCSR[ 175 ][ 337 ],
   alphaCSR[ 175 ][ 338 ],
   alphaCSR[ 175 ][ 339 ],
   alphaCSR[ 175 ][ 340 ],
   alphaCSR[ 175 ][ 341 ],
   alphaCSR[ 175 ][ 342 ],
   alphaCSR[ 175 ][ 343 ],
   alphaCSR[ 175 ][ 344 ],
   alphaCSR[ 175 ][ 345 ],
   alphaCSR[ 175 ][ 346 ],
   alphaCSR[ 175 ][ 347 ],
   alphaCSR[ 175 ][ 348 ],
   alphaCSR[ 175 ][ 349 ],
   alphaCSR[ 175 ][ 350 ],
   alphaCSR[ 175 ][ 351 ],
   alphaCSR[ 175 ][ 352 ],
   alphaCSR[ 175 ][ 353 ],
   alphaCSR[ 175 ][ 354 ],
   alphaCSR[ 175 ][ 355 ],
   alphaCSR[ 175 ][ 356 ],
   alphaCSR[ 175 ][ 357 ],
   alphaCSR[ 175 ][ 358 ],
   alphaCSR[ 175 ][ 359 ],
   alphaCSR[ 175 ][ 360 ],
   alphaCSR[ 175 ][ 361 ],
   alphaCSR[ 175 ][ 362 ],
   alphaCSR[ 175 ][ 363 ],
   alphaCSR[ 175 ][ 364 ],
   alphaCSR[ 175 ][ 365 ],
   alphaCSR[ 175 ][ 366 ],
   alphaCSR[ 175 ][ 367 ],
   alphaCSR[ 175 ][ 368 ],
   alphaCSR[ 175 ][ 369 ],
   alphaCSR[ 175 ][ 370 ],
   alphaCSR[ 175 ][ 371 ],
   alphaCSR[ 175 ][ 372 ],
   alphaCSR[ 175 ][ 373 ],
   alphaCSR[ 175 ][ 374 ],
   alphaCSR[ 175 ][ 375 ],
   alphaCSR[ 175 ][ 376 ],
   alphaCSR[ 175 ][ 377 ],
   alphaCSR[ 175 ][ 378 ],
   alphaCSR[ 175 ][ 379 ],
   alphaCSR[ 175 ][ 380 ],
   alphaCSR[ 175 ][ 381 ],
   alphaCSR[ 175 ][ 382 ],
   alphaCSR[ 175 ][ 383 ],
   alphaCSR[ 176 ][ 0 ],
   alphaCSR[ 176 ][ 1 ],
   alphaCSR[ 176 ][ 2 ],
   alphaCSR[ 176 ][ 3 ],
   alphaCSR[ 176 ][ 4 ],
   alphaCSR[ 176 ][ 5 ],
   alphaCSR[ 176 ][ 6 ],
   alphaCSR[ 176 ][ 7 ],
   alphaCSR[ 176 ][ 8 ],
   alphaCSR[ 176 ][ 9 ],
   alphaCSR[ 176 ][ 10 ],
   alphaCSR[ 176 ][ 11 ],
   alphaCSR[ 176 ][ 12 ],
   alphaCSR[ 176 ][ 13 ],
   alphaCSR[ 176 ][ 14 ],
   alphaCSR[ 176 ][ 15 ],
   alphaCSR[ 176 ][ 16 ],
   alphaCSR[ 176 ][ 17 ],
   alphaCSR[ 176 ][ 18 ],
   alphaCSR[ 176 ][ 19 ],
   alphaCSR[ 176 ][ 20 ],
   alphaCSR[ 176 ][ 21 ],
   alphaCSR[ 176 ][ 22 ],
   alphaCSR[ 176 ][ 23 ],
   alphaCSR[ 176 ][ 24 ],
   alphaCSR[ 176 ][ 25 ],
   alphaCSR[ 176 ][ 26 ],
   alphaCSR[ 176 ][ 27 ],
   alphaCSR[ 176 ][ 28 ],
   alphaCSR[ 176 ][ 29 ],
   alphaCSR[ 176 ][ 30 ],
   alphaCSR[ 176 ][ 31 ],
   alphaCSR[ 176 ][ 32 ],
   alphaCSR[ 176 ][ 33 ],
   alphaCSR[ 176 ][ 34 ],
   alphaCSR[ 176 ][ 35 ],
   alphaCSR[ 176 ][ 36 ],
   alphaCSR[ 176 ][ 37 ],
   alphaCSR[ 176 ][ 38 ],
   alphaCSR[ 176 ][ 39 ],
   alphaCSR[ 176 ][ 40 ],
   alphaCSR[ 176 ][ 41 ],
   alphaCSR[ 176 ][ 42 ],
   alphaCSR[ 176 ][ 43 ],
   alphaCSR[ 176 ][ 44 ],
   alphaCSR[ 176 ][ 45 ],
   alphaCSR[ 176 ][ 46 ],
   alphaCSR[ 176 ][ 47 ],
   alphaCSR[ 176 ][ 48 ],
   alphaCSR[ 176 ][ 49 ],
   alphaCSR[ 176 ][ 50 ],
   alphaCSR[ 176 ][ 51 ],
   alphaCSR[ 176 ][ 52 ],
   alphaCSR[ 176 ][ 53 ],
   alphaCSR[ 176 ][ 54 ],
   alphaCSR[ 176 ][ 55 ],
   alphaCSR[ 176 ][ 56 ],
   alphaCSR[ 176 ][ 57 ],
   alphaCSR[ 176 ][ 58 ],
   alphaCSR[ 176 ][ 59 ],
   alphaCSR[ 176 ][ 60 ],
   alphaCSR[ 176 ][ 61 ],
   alphaCSR[ 176 ][ 62 ],
   alphaCSR[ 176 ][ 63 ],
   alphaCSR[ 176 ][ 64 ],
   alphaCSR[ 176 ][ 65 ],
   alphaCSR[ 176 ][ 66 ],
   alphaCSR[ 176 ][ 67 ],
   alphaCSR[ 176 ][ 68 ],
   alphaCSR[ 176 ][ 69 ],
   alphaCSR[ 176 ][ 70 ],
   alphaCSR[ 176 ][ 71 ],
   alphaCSR[ 176 ][ 72 ],
   alphaCSR[ 176 ][ 73 ],
   alphaCSR[ 176 ][ 74 ],
   alphaCSR[ 176 ][ 75 ],
   alphaCSR[ 176 ][ 76 ],
   alphaCSR[ 176 ][ 77 ],
   alphaCSR[ 176 ][ 78 ],
   alphaCSR[ 176 ][ 79 ],
   alphaCSR[ 176 ][ 80 ],
   alphaCSR[ 176 ][ 81 ],
   alphaCSR[ 176 ][ 82 ],
   alphaCSR[ 176 ][ 83 ],
   alphaCSR[ 176 ][ 84 ],
   alphaCSR[ 176 ][ 85 ],
   alphaCSR[ 176 ][ 86 ],
   alphaCSR[ 176 ][ 87 ],
   alphaCSR[ 176 ][ 88 ],
   alphaCSR[ 176 ][ 89 ],
   alphaCSR[ 176 ][ 90 ],
   alphaCSR[ 176 ][ 91 ],
   alphaCSR[ 176 ][ 92 ],
   alphaCSR[ 176 ][ 93 ],
   alphaCSR[ 176 ][ 94 ],
   alphaCSR[ 176 ][ 95 ],
   alphaCSR[ 176 ][ 96 ],
   alphaCSR[ 176 ][ 97 ],
   alphaCSR[ 176 ][ 98 ],
   alphaCSR[ 176 ][ 99 ],
   alphaCSR[ 176 ][ 100 ],
   alphaCSR[ 176 ][ 101 ],
   alphaCSR[ 176 ][ 102 ],
   alphaCSR[ 176 ][ 103 ],
   alphaCSR[ 176 ][ 104 ],
   alphaCSR[ 176 ][ 105 ],
   alphaCSR[ 176 ][ 106 ],
   alphaCSR[ 176 ][ 107 ],
   alphaCSR[ 176 ][ 108 ],
   alphaCSR[ 176 ][ 109 ],
   alphaCSR[ 176 ][ 110 ],
   alphaCSR[ 176 ][ 111 ],
   alphaCSR[ 176 ][ 112 ],
   alphaCSR[ 176 ][ 113 ],
   alphaCSR[ 176 ][ 114 ],
   alphaCSR[ 176 ][ 115 ],
   alphaCSR[ 176 ][ 116 ],
   alphaCSR[ 176 ][ 117 ],
   alphaCSR[ 176 ][ 118 ],
   alphaCSR[ 176 ][ 119 ],
   alphaCSR[ 176 ][ 120 ],
   alphaCSR[ 176 ][ 121 ],
   alphaCSR[ 176 ][ 122 ],
   alphaCSR[ 176 ][ 123 ],
   alphaCSR[ 176 ][ 124 ],
   alphaCSR[ 176 ][ 125 ],
   alphaCSR[ 176 ][ 126 ],
   alphaCSR[ 176 ][ 127 ],
   alphaCSR[ 176 ][ 128 ],
   alphaCSR[ 176 ][ 129 ],
   alphaCSR[ 176 ][ 130 ],
   alphaCSR[ 176 ][ 131 ],
   alphaCSR[ 176 ][ 132 ],
   alphaCSR[ 176 ][ 133 ],
   alphaCSR[ 176 ][ 134 ],
   alphaCSR[ 176 ][ 135 ],
   alphaCSR[ 176 ][ 136 ],
   alphaCSR[ 176 ][ 137 ],
   alphaCSR[ 176 ][ 138 ],
   alphaCSR[ 176 ][ 139 ],
   alphaCSR[ 176 ][ 140 ],
   alphaCSR[ 176 ][ 141 ],
   alphaCSR[ 176 ][ 142 ],
   alphaCSR[ 176 ][ 143 ],
   alphaCSR[ 176 ][ 144 ],
   alphaCSR[ 176 ][ 145 ],
   alphaCSR[ 176 ][ 146 ],
   alphaCSR[ 176 ][ 147 ],
   alphaCSR[ 176 ][ 148 ],
   alphaCSR[ 176 ][ 149 ],
   alphaCSR[ 176 ][ 150 ],
   alphaCSR[ 176 ][ 151 ],
   alphaCSR[ 176 ][ 152 ],
   alphaCSR[ 176 ][ 153 ],
   alphaCSR[ 176 ][ 154 ],
   alphaCSR[ 176 ][ 155 ],
   alphaCSR[ 176 ][ 156 ],
   alphaCSR[ 176 ][ 157 ],
   alphaCSR[ 176 ][ 158 ],
   alphaCSR[ 176 ][ 159 ],
   alphaCSR[ 176 ][ 160 ],
   alphaCSR[ 176 ][ 161 ],
   alphaCSR[ 176 ][ 162 ],
   alphaCSR[ 176 ][ 163 ],
   alphaCSR[ 176 ][ 164 ],
   alphaCSR[ 176 ][ 165 ],
   alphaCSR[ 176 ][ 166 ],
   alphaCSR[ 176 ][ 167 ],
   alphaCSR[ 176 ][ 168 ],
   alphaCSR[ 176 ][ 169 ],
   alphaCSR[ 176 ][ 170 ],
   alphaCSR[ 176 ][ 171 ],
   alphaCSR[ 176 ][ 172 ],
   alphaCSR[ 176 ][ 173 ],
   alphaCSR[ 176 ][ 174 ],
   alphaCSR[ 176 ][ 175 ],
   alphaCSR[ 176 ][ 176 ],
   alphaCSR[ 176 ][ 177 ],
   alphaCSR[ 176 ][ 178 ],
   alphaCSR[ 176 ][ 179 ],
   alphaCSR[ 176 ][ 180 ],
   alphaCSR[ 176 ][ 181 ],
   alphaCSR[ 176 ][ 182 ],
   alphaCSR[ 176 ][ 183 ],
   alphaCSR[ 176 ][ 184 ],
   alphaCSR[ 176 ][ 185 ],
   alphaCSR[ 176 ][ 186 ],
   alphaCSR[ 176 ][ 187 ],
   alphaCSR[ 176 ][ 188 ],
   alphaCSR[ 176 ][ 189 ],
   alphaCSR[ 176 ][ 190 ],
   alphaCSR[ 176 ][ 191 ],
   alphaCSR[ 176 ][ 192 ],
   alphaCSR[ 176 ][ 193 ],
   alphaCSR[ 176 ][ 194 ],
   alphaCSR[ 176 ][ 195 ],
   alphaCSR[ 176 ][ 196 ],
   alphaCSR[ 176 ][ 197 ],
   alphaCSR[ 176 ][ 198 ],
   alphaCSR[ 176 ][ 199 ],
   alphaCSR[ 176 ][ 200 ],
   alphaCSR[ 176 ][ 201 ],
   alphaCSR[ 176 ][ 202 ],
   alphaCSR[ 176 ][ 203 ],
   alphaCSR[ 176 ][ 204 ],
   alphaCSR[ 176 ][ 205 ],
   alphaCSR[ 176 ][ 206 ],
   alphaCSR[ 176 ][ 207 ],
   alphaCSR[ 176 ][ 208 ],
   alphaCSR[ 176 ][ 209 ],
   alphaCSR[ 176 ][ 210 ],
   alphaCSR[ 176 ][ 211 ],
   alphaCSR[ 176 ][ 212 ],
   alphaCSR[ 176 ][ 213 ],
   alphaCSR[ 176 ][ 214 ],
   alphaCSR[ 176 ][ 215 ],
   alphaCSR[ 176 ][ 216 ],
   alphaCSR[ 176 ][ 217 ],
   alphaCSR[ 176 ][ 218 ],
   alphaCSR[ 176 ][ 219 ],
   alphaCSR[ 176 ][ 220 ],
   alphaCSR[ 176 ][ 221 ],
   alphaCSR[ 176 ][ 222 ],
   alphaCSR[ 176 ][ 223 ],
   alphaCSR[ 176 ][ 224 ],
   alphaCSR[ 176 ][ 225 ],
   alphaCSR[ 176 ][ 226 ],
   alphaCSR[ 176 ][ 227 ],
   alphaCSR[ 176 ][ 228 ],
   alphaCSR[ 176 ][ 229 ],
   alphaCSR[ 176 ][ 230 ],
   alphaCSR[ 176 ][ 231 ],
   alphaCSR[ 176 ][ 232 ],
   alphaCSR[ 176 ][ 233 ],
   alphaCSR[ 176 ][ 234 ],
   alphaCSR[ 176 ][ 235 ],
   alphaCSR[ 176 ][ 236 ],
   alphaCSR[ 176 ][ 237 ],
   alphaCSR[ 176 ][ 238 ],
   alphaCSR[ 176 ][ 239 ],
   alphaCSR[ 176 ][ 240 ],
   alphaCSR[ 176 ][ 241 ],
   alphaCSR[ 176 ][ 242 ],
   alphaCSR[ 176 ][ 243 ],
   alphaCSR[ 176 ][ 244 ],
   alphaCSR[ 176 ][ 245 ],
   alphaCSR[ 176 ][ 246 ],
   alphaCSR[ 176 ][ 247 ],
   alphaCSR[ 176 ][ 248 ],
   alphaCSR[ 176 ][ 249 ],
   alphaCSR[ 176 ][ 250 ],
   alphaCSR[ 176 ][ 251 ],
   alphaCSR[ 176 ][ 252 ],
   alphaCSR[ 176 ][ 253 ],
   alphaCSR[ 176 ][ 254 ],
   alphaCSR[ 176 ][ 255 ],
   alphaCSR[ 176 ][ 256 ],
   alphaCSR[ 176 ][ 257 ],
   alphaCSR[ 176 ][ 258 ],
   alphaCSR[ 176 ][ 259 ],
   alphaCSR[ 176 ][ 260 ],
   alphaCSR[ 176 ][ 261 ],
   alphaCSR[ 176 ][ 262 ],
   alphaCSR[ 176 ][ 263 ],
   alphaCSR[ 176 ][ 264 ],
   alphaCSR[ 176 ][ 265 ],
   alphaCSR[ 176 ][ 266 ],
   alphaCSR[ 176 ][ 267 ],
   alphaCSR[ 176 ][ 268 ],
   alphaCSR[ 176 ][ 269 ],
   alphaCSR[ 176 ][ 270 ],
   alphaCSR[ 176 ][ 271 ],
   alphaCSR[ 176 ][ 272 ],
   alphaCSR[ 176 ][ 273 ],
   alphaCSR[ 176 ][ 274 ],
   alphaCSR[ 176 ][ 275 ],
   alphaCSR[ 176 ][ 276 ],
   alphaCSR[ 176 ][ 277 ],
   alphaCSR[ 176 ][ 278 ],
   alphaCSR[ 176 ][ 279 ],
   alphaCSR[ 176 ][ 280 ],
   alphaCSR[ 176 ][ 281 ],
   alphaCSR[ 176 ][ 282 ],
   alphaCSR[ 176 ][ 283 ],
   alphaCSR[ 176 ][ 284 ],
   alphaCSR[ 176 ][ 285 ],
   alphaCSR[ 176 ][ 286 ],
   alphaCSR[ 176 ][ 287 ],
   alphaCSR[ 176 ][ 288 ],
   alphaCSR[ 176 ][ 289 ],
   alphaCSR[ 176 ][ 290 ],
   alphaCSR[ 176 ][ 291 ],
   alphaCSR[ 176 ][ 292 ],
   alphaCSR[ 176 ][ 293 ],
   alphaCSR[ 176 ][ 294 ],
   alphaCSR[ 176 ][ 295 ],
   alphaCSR[ 176 ][ 296 ],
   alphaCSR[ 176 ][ 297 ],
   alphaCSR[ 176 ][ 298 ],
   alphaCSR[ 176 ][ 299 ],
   alphaCSR[ 176 ][ 300 ],
   alphaCSR[ 176 ][ 301 ],
   alphaCSR[ 176 ][ 302 ],
   alphaCSR[ 176 ][ 303 ],
   alphaCSR[ 176 ][ 304 ],
   alphaCSR[ 176 ][ 305 ],
   alphaCSR[ 176 ][ 306 ],
   alphaCSR[ 176 ][ 307 ],
   alphaCSR[ 176 ][ 308 ],
   alphaCSR[ 176 ][ 309 ],
   alphaCSR[ 176 ][ 310 ],
   alphaCSR[ 176 ][ 311 ],
   alphaCSR[ 176 ][ 312 ],
   alphaCSR[ 176 ][ 313 ],
   alphaCSR[ 176 ][ 314 ],
   alphaCSR[ 176 ][ 315 ],
   alphaCSR[ 176 ][ 316 ],
   alphaCSR[ 176 ][ 317 ],
   alphaCSR[ 176 ][ 318 ],
   alphaCSR[ 176 ][ 319 ],
   alphaCSR[ 176 ][ 320 ],
   alphaCSR[ 176 ][ 321 ],
   alphaCSR[ 176 ][ 322 ],
   alphaCSR[ 176 ][ 323 ],
   alphaCSR[ 176 ][ 324 ],
   alphaCSR[ 176 ][ 325 ],
   alphaCSR[ 176 ][ 326 ],
   alphaCSR[ 176 ][ 327 ],
   alphaCSR[ 176 ][ 328 ],
   alphaCSR[ 176 ][ 329 ],
   alphaCSR[ 176 ][ 330 ],
   alphaCSR[ 176 ][ 331 ],
   alphaCSR[ 176 ][ 332 ],
   alphaCSR[ 176 ][ 333 ],
   alphaCSR[ 176 ][ 334 ],
   alphaCSR[ 176 ][ 335 ],
   alphaCSR[ 176 ][ 336 ],
   alphaCSR[ 176 ][ 337 ],
   alphaCSR[ 176 ][ 338 ],
   alphaCSR[ 176 ][ 339 ],
   alphaCSR[ 176 ][ 340 ],
   alphaCSR[ 176 ][ 341 ],
   alphaCSR[ 176 ][ 342 ],
   alphaCSR[ 176 ][ 343 ],
   alphaCSR[ 176 ][ 344 ],
   alphaCSR[ 176 ][ 345 ],
   alphaCSR[ 176 ][ 346 ],
   alphaCSR[ 176 ][ 347 ],
   alphaCSR[ 176 ][ 348 ],
   alphaCSR[ 176 ][ 349 ],
   alphaCSR[ 176 ][ 350 ],
   alphaCSR[ 176 ][ 351 ],
   alphaCSR[ 176 ][ 352 ],
   alphaCSR[ 176 ][ 353 ],
   alphaCSR[ 176 ][ 354 ],
   alphaCSR[ 176 ][ 355 ],
   alphaCSR[ 176 ][ 356 ],
   alphaCSR[ 176 ][ 357 ],
   alphaCSR[ 176 ][ 358 ],
   alphaCSR[ 176 ][ 359 ],
   alphaCSR[ 176 ][ 360 ],
   alphaCSR[ 176 ][ 361 ],
   alphaCSR[ 176 ][ 362 ],
   alphaCSR[ 176 ][ 363 ],
   alphaCSR[ 176 ][ 364 ],
   alphaCSR[ 176 ][ 365 ],
   alphaCSR[ 176 ][ 366 ],
   alphaCSR[ 176 ][ 367 ],
   alphaCSR[ 176 ][ 368 ],
   alphaCSR[ 176 ][ 369 ],
   alphaCSR[ 176 ][ 370 ],
   alphaCSR[ 176 ][ 371 ],
   alphaCSR[ 176 ][ 372 ],
   alphaCSR[ 176 ][ 373 ],
   alphaCSR[ 176 ][ 374 ],
   alphaCSR[ 176 ][ 375 ],
   alphaCSR[ 176 ][ 376 ],
   alphaCSR[ 176 ][ 377 ],
   alphaCSR[ 176 ][ 378 ],
   alphaCSR[ 176 ][ 379 ],
   alphaCSR[ 176 ][ 380 ],
   alphaCSR[ 176 ][ 381 ],
   alphaCSR[ 176 ][ 382 ],
   alphaCSR[ 176 ][ 383 ],
   alphaCSR[ 177 ][ 0 ],
   alphaCSR[ 177 ][ 1 ],
   alphaCSR[ 177 ][ 2 ],
   alphaCSR[ 177 ][ 3 ],
   alphaCSR[ 177 ][ 4 ],
   alphaCSR[ 177 ][ 5 ],
   alphaCSR[ 177 ][ 6 ],
   alphaCSR[ 177 ][ 7 ],
   alphaCSR[ 177 ][ 8 ],
   alphaCSR[ 177 ][ 9 ],
   alphaCSR[ 177 ][ 10 ],
   alphaCSR[ 177 ][ 11 ],
   alphaCSR[ 177 ][ 12 ],
   alphaCSR[ 177 ][ 13 ],
   alphaCSR[ 177 ][ 14 ],
   alphaCSR[ 177 ][ 15 ],
   alphaCSR[ 177 ][ 16 ],
   alphaCSR[ 177 ][ 17 ],
   alphaCSR[ 177 ][ 18 ],
   alphaCSR[ 177 ][ 19 ],
   alphaCSR[ 177 ][ 20 ],
   alphaCSR[ 177 ][ 21 ],
   alphaCSR[ 177 ][ 22 ],
   alphaCSR[ 177 ][ 23 ],
   alphaCSR[ 177 ][ 24 ],
   alphaCSR[ 177 ][ 25 ],
   alphaCSR[ 177 ][ 26 ],
   alphaCSR[ 177 ][ 27 ],
   alphaCSR[ 177 ][ 28 ],
   alphaCSR[ 177 ][ 29 ],
   alphaCSR[ 177 ][ 30 ],
   alphaCSR[ 177 ][ 31 ],
   alphaCSR[ 177 ][ 32 ],
   alphaCSR[ 177 ][ 33 ],
   alphaCSR[ 177 ][ 34 ],
   alphaCSR[ 177 ][ 35 ],
   alphaCSR[ 177 ][ 36 ],
   alphaCSR[ 177 ][ 37 ],
   alphaCSR[ 177 ][ 38 ],
   alphaCSR[ 177 ][ 39 ],
   alphaCSR[ 177 ][ 40 ],
   alphaCSR[ 177 ][ 41 ],
   alphaCSR[ 177 ][ 42 ],
   alphaCSR[ 177 ][ 43 ],
   alphaCSR[ 177 ][ 44 ],
   alphaCSR[ 177 ][ 45 ],
   alphaCSR[ 177 ][ 46 ],
   alphaCSR[ 177 ][ 47 ],
   alphaCSR[ 177 ][ 48 ],
   alphaCSR[ 177 ][ 49 ],
   alphaCSR[ 177 ][ 50 ],
   alphaCSR[ 177 ][ 51 ],
   alphaCSR[ 177 ][ 52 ],
   alphaCSR[ 177 ][ 53 ],
   alphaCSR[ 177 ][ 54 ],
   alphaCSR[ 177 ][ 55 ],
   alphaCSR[ 177 ][ 56 ],
   alphaCSR[ 177 ][ 57 ],
   alphaCSR[ 177 ][ 58 ],
   alphaCSR[ 177 ][ 59 ],
   alphaCSR[ 177 ][ 60 ],
   alphaCSR[ 177 ][ 61 ],
   alphaCSR[ 177 ][ 62 ],
   alphaCSR[ 177 ][ 63 ],
   alphaCSR[ 177 ][ 64 ],
   alphaCSR[ 177 ][ 65 ],
   alphaCSR[ 177 ][ 66 ],
   alphaCSR[ 177 ][ 67 ],
   alphaCSR[ 177 ][ 68 ],
   alphaCSR[ 177 ][ 69 ],
   alphaCSR[ 177 ][ 70 ],
   alphaCSR[ 177 ][ 71 ],
   alphaCSR[ 177 ][ 72 ],
   alphaCSR[ 177 ][ 73 ],
   alphaCSR[ 177 ][ 74 ],
   alphaCSR[ 177 ][ 75 ],
   alphaCSR[ 177 ][ 76 ],
   alphaCSR[ 177 ][ 77 ],
   alphaCSR[ 177 ][ 78 ],
   alphaCSR[ 177 ][ 79 ],
   alphaCSR[ 177 ][ 80 ],
   alphaCSR[ 177 ][ 81 ],
   alphaCSR[ 177 ][ 82 ],
   alphaCSR[ 177 ][ 83 ],
   alphaCSR[ 177 ][ 84 ],
   alphaCSR[ 177 ][ 85 ],
   alphaCSR[ 177 ][ 86 ],
   alphaCSR[ 177 ][ 87 ],
   alphaCSR[ 177 ][ 88 ],
   alphaCSR[ 177 ][ 89 ],
   alphaCSR[ 177 ][ 90 ],
   alphaCSR[ 177 ][ 91 ],
   alphaCSR[ 177 ][ 92 ],
   alphaCSR[ 177 ][ 93 ],
   alphaCSR[ 177 ][ 94 ],
   alphaCSR[ 177 ][ 95 ],
   alphaCSR[ 177 ][ 96 ],
   alphaCSR[ 177 ][ 97 ],
   alphaCSR[ 177 ][ 98 ],
   alphaCSR[ 177 ][ 99 ],
   alphaCSR[ 177 ][ 100 ],
   alphaCSR[ 177 ][ 101 ],
   alphaCSR[ 177 ][ 102 ],
   alphaCSR[ 177 ][ 103 ],
   alphaCSR[ 177 ][ 104 ],
   alphaCSR[ 177 ][ 105 ],
   alphaCSR[ 177 ][ 106 ],
   alphaCSR[ 177 ][ 107 ],
   alphaCSR[ 177 ][ 108 ],
   alphaCSR[ 177 ][ 109 ],
   alphaCSR[ 177 ][ 110 ],
   alphaCSR[ 177 ][ 111 ],
   alphaCSR[ 177 ][ 112 ],
   alphaCSR[ 177 ][ 113 ],
   alphaCSR[ 177 ][ 114 ],
   alphaCSR[ 177 ][ 115 ],
   alphaCSR[ 177 ][ 116 ],
   alphaCSR[ 177 ][ 117 ],
   alphaCSR[ 177 ][ 118 ],
   alphaCSR[ 177 ][ 119 ],
   alphaCSR[ 177 ][ 120 ],
   alphaCSR[ 177 ][ 121 ],
   alphaCSR[ 177 ][ 122 ],
   alphaCSR[ 177 ][ 123 ],
   alphaCSR[ 177 ][ 124 ],
   alphaCSR[ 177 ][ 125 ],
   alphaCSR[ 177 ][ 126 ],
   alphaCSR[ 177 ][ 127 ],
   alphaCSR[ 177 ][ 128 ],
   alphaCSR[ 177 ][ 129 ],
   alphaCSR[ 177 ][ 130 ],
   alphaCSR[ 177 ][ 131 ],
   alphaCSR[ 177 ][ 132 ],
   alphaCSR[ 177 ][ 133 ],
   alphaCSR[ 177 ][ 134 ],
   alphaCSR[ 177 ][ 135 ],
   alphaCSR[ 177 ][ 136 ],
   alphaCSR[ 177 ][ 137 ],
   alphaCSR[ 177 ][ 138 ],
   alphaCSR[ 177 ][ 139 ],
   alphaCSR[ 177 ][ 140 ],
   alphaCSR[ 177 ][ 141 ],
   alphaCSR[ 177 ][ 142 ],
   alphaCSR[ 177 ][ 143 ],
   alphaCSR[ 177 ][ 144 ],
   alphaCSR[ 177 ][ 145 ],
   alphaCSR[ 177 ][ 146 ],
   alphaCSR[ 177 ][ 147 ],
   alphaCSR[ 177 ][ 148 ],
   alphaCSR[ 177 ][ 149 ],
   alphaCSR[ 177 ][ 150 ],
   alphaCSR[ 177 ][ 151 ],
   alphaCSR[ 177 ][ 152 ],
   alphaCSR[ 177 ][ 153 ],
   alphaCSR[ 177 ][ 154 ],
   alphaCSR[ 177 ][ 155 ],
   alphaCSR[ 177 ][ 156 ],
   alphaCSR[ 177 ][ 157 ],
   alphaCSR[ 177 ][ 158 ],
   alphaCSR[ 177 ][ 159 ],
   alphaCSR[ 177 ][ 160 ],
   alphaCSR[ 177 ][ 161 ],
   alphaCSR[ 177 ][ 162 ],
   alphaCSR[ 177 ][ 163 ],
   alphaCSR[ 177 ][ 164 ],
   alphaCSR[ 177 ][ 165 ],
   alphaCSR[ 177 ][ 166 ],
   alphaCSR[ 177 ][ 167 ],
   alphaCSR[ 177 ][ 168 ],
   alphaCSR[ 177 ][ 169 ],
   alphaCSR[ 177 ][ 170 ],
   alphaCSR[ 177 ][ 171 ],
   alphaCSR[ 177 ][ 172 ],
   alphaCSR[ 177 ][ 173 ],
   alphaCSR[ 177 ][ 174 ],
   alphaCSR[ 177 ][ 175 ],
   alphaCSR[ 177 ][ 176 ],
   alphaCSR[ 177 ][ 177 ],
   alphaCSR[ 177 ][ 178 ],
   alphaCSR[ 177 ][ 179 ],
   alphaCSR[ 177 ][ 180 ],
   alphaCSR[ 177 ][ 181 ],
   alphaCSR[ 177 ][ 182 ],
   alphaCSR[ 177 ][ 183 ],
   alphaCSR[ 177 ][ 184 ],
   alphaCSR[ 177 ][ 185 ],
   alphaCSR[ 177 ][ 186 ],
   alphaCSR[ 177 ][ 187 ],
   alphaCSR[ 177 ][ 188 ],
   alphaCSR[ 177 ][ 189 ],
   alphaCSR[ 177 ][ 190 ],
   alphaCSR[ 177 ][ 191 ],
   alphaCSR[ 177 ][ 192 ],
   alphaCSR[ 177 ][ 193 ],
   alphaCSR[ 177 ][ 194 ],
   alphaCSR[ 177 ][ 195 ],
   alphaCSR[ 177 ][ 196 ],
   alphaCSR[ 177 ][ 197 ],
   alphaCSR[ 177 ][ 198 ],
   alphaCSR[ 177 ][ 199 ],
   alphaCSR[ 177 ][ 200 ],
   alphaCSR[ 177 ][ 201 ],
   alphaCSR[ 177 ][ 202 ],
   alphaCSR[ 177 ][ 203 ],
   alphaCSR[ 177 ][ 204 ],
   alphaCSR[ 177 ][ 205 ],
   alphaCSR[ 177 ][ 206 ],
   alphaCSR[ 177 ][ 207 ],
   alphaCSR[ 177 ][ 208 ],
   alphaCSR[ 177 ][ 209 ],
   alphaCSR[ 177 ][ 210 ],
   alphaCSR[ 177 ][ 211 ],
   alphaCSR[ 177 ][ 212 ],
   alphaCSR[ 177 ][ 213 ],
   alphaCSR[ 177 ][ 214 ],
   alphaCSR[ 177 ][ 215 ],
   alphaCSR[ 177 ][ 216 ],
   alphaCSR[ 177 ][ 217 ],
   alphaCSR[ 177 ][ 218 ],
   alphaCSR[ 177 ][ 219 ],
   alphaCSR[ 177 ][ 220 ],
   alphaCSR[ 177 ][ 221 ],
   alphaCSR[ 177 ][ 222 ],
   alphaCSR[ 177 ][ 223 ],
   alphaCSR[ 177 ][ 224 ],
   alphaCSR[ 177 ][ 225 ],
   alphaCSR[ 177 ][ 226 ],
   alphaCSR[ 177 ][ 227 ],
   alphaCSR[ 177 ][ 228 ],
   alphaCSR[ 177 ][ 229 ],
   alphaCSR[ 177 ][ 230 ],
   alphaCSR[ 177 ][ 231 ],
   alphaCSR[ 177 ][ 232 ],
   alphaCSR[ 177 ][ 233 ],
   alphaCSR[ 177 ][ 234 ],
   alphaCSR[ 177 ][ 235 ],
   alphaCSR[ 177 ][ 236 ],
   alphaCSR[ 177 ][ 237 ],
   alphaCSR[ 177 ][ 238 ],
   alphaCSR[ 177 ][ 239 ],
   alphaCSR[ 177 ][ 240 ],
   alphaCSR[ 177 ][ 241 ],
   alphaCSR[ 177 ][ 242 ],
   alphaCSR[ 177 ][ 243 ],
   alphaCSR[ 177 ][ 244 ],
   alphaCSR[ 177 ][ 245 ],
   alphaCSR[ 177 ][ 246 ],
   alphaCSR[ 177 ][ 247 ],
   alphaCSR[ 177 ][ 248 ],
   alphaCSR[ 177 ][ 249 ],
   alphaCSR[ 177 ][ 250 ],
   alphaCSR[ 177 ][ 251 ],
   alphaCSR[ 177 ][ 252 ],
   alphaCSR[ 177 ][ 253 ],
   alphaCSR[ 177 ][ 254 ],
   alphaCSR[ 177 ][ 255 ],
   alphaCSR[ 177 ][ 256 ],
   alphaCSR[ 177 ][ 257 ],
   alphaCSR[ 177 ][ 258 ],
   alphaCSR[ 177 ][ 259 ],
   alphaCSR[ 177 ][ 260 ],
   alphaCSR[ 177 ][ 261 ],
   alphaCSR[ 177 ][ 262 ],
   alphaCSR[ 177 ][ 263 ],
   alphaCSR[ 177 ][ 264 ],
   alphaCSR[ 177 ][ 265 ],
   alphaCSR[ 177 ][ 266 ],
   alphaCSR[ 177 ][ 267 ],
   alphaCSR[ 177 ][ 268 ],
   alphaCSR[ 177 ][ 269 ],
   alphaCSR[ 177 ][ 270 ],
   alphaCSR[ 177 ][ 271 ],
   alphaCSR[ 177 ][ 272 ],
   alphaCSR[ 177 ][ 273 ],
   alphaCSR[ 177 ][ 274 ],
   alphaCSR[ 177 ][ 275 ],
   alphaCSR[ 177 ][ 276 ],
   alphaCSR[ 177 ][ 277 ],
   alphaCSR[ 177 ][ 278 ],
   alphaCSR[ 177 ][ 279 ],
   alphaCSR[ 177 ][ 280 ],
   alphaCSR[ 177 ][ 281 ],
   alphaCSR[ 177 ][ 282 ],
   alphaCSR[ 177 ][ 283 ],
   alphaCSR[ 177 ][ 284 ],
   alphaCSR[ 177 ][ 285 ],
   alphaCSR[ 177 ][ 286 ],
   alphaCSR[ 177 ][ 287 ],
   alphaCSR[ 177 ][ 288 ],
   alphaCSR[ 177 ][ 289 ],
   alphaCSR[ 177 ][ 290 ],
   alphaCSR[ 177 ][ 291 ],
   alphaCSR[ 177 ][ 292 ],
   alphaCSR[ 177 ][ 293 ],
   alphaCSR[ 177 ][ 294 ],
   alphaCSR[ 177 ][ 295 ],
   alphaCSR[ 177 ][ 296 ],
   alphaCSR[ 177 ][ 297 ],
   alphaCSR[ 177 ][ 298 ],
   alphaCSR[ 177 ][ 299 ],
   alphaCSR[ 177 ][ 300 ],
   alphaCSR[ 177 ][ 301 ],
   alphaCSR[ 177 ][ 302 ],
   alphaCSR[ 177 ][ 303 ],
   alphaCSR[ 177 ][ 304 ],
   alphaCSR[ 177 ][ 305 ],
   alphaCSR[ 177 ][ 306 ],
   alphaCSR[ 177 ][ 307 ],
   alphaCSR[ 177 ][ 308 ],
   alphaCSR[ 177 ][ 309 ],
   alphaCSR[ 177 ][ 310 ],
   alphaCSR[ 177 ][ 311 ],
   alphaCSR[ 177 ][ 312 ],
   alphaCSR[ 177 ][ 313 ],
   alphaCSR[ 177 ][ 314 ],
   alphaCSR[ 177 ][ 315 ],
   alphaCSR[ 177 ][ 316 ],
   alphaCSR[ 177 ][ 317 ],
   alphaCSR[ 177 ][ 318 ],
   alphaCSR[ 177 ][ 319 ],
   alphaCSR[ 177 ][ 320 ],
   alphaCSR[ 177 ][ 321 ],
   alphaCSR[ 177 ][ 322 ],
   alphaCSR[ 177 ][ 323 ],
   alphaCSR[ 177 ][ 324 ],
   alphaCSR[ 177 ][ 325 ],
   alphaCSR[ 177 ][ 326 ],
   alphaCSR[ 177 ][ 327 ],
   alphaCSR[ 177 ][ 328 ],
   alphaCSR[ 177 ][ 329 ],
   alphaCSR[ 177 ][ 330 ],
   alphaCSR[ 177 ][ 331 ],
   alphaCSR[ 177 ][ 332 ],
   alphaCSR[ 177 ][ 333 ],
   alphaCSR[ 177 ][ 334 ],
   alphaCSR[ 177 ][ 335 ],
   alphaCSR[ 177 ][ 336 ],
   alphaCSR[ 177 ][ 337 ],
   alphaCSR[ 177 ][ 338 ],
   alphaCSR[ 177 ][ 339 ],
   alphaCSR[ 177 ][ 340 ],
   alphaCSR[ 177 ][ 341 ],
   alphaCSR[ 177 ][ 342 ],
   alphaCSR[ 177 ][ 343 ],
   alphaCSR[ 177 ][ 344 ],
   alphaCSR[ 177 ][ 345 ],
   alphaCSR[ 177 ][ 346 ],
   alphaCSR[ 177 ][ 347 ],
   alphaCSR[ 177 ][ 348 ],
   alphaCSR[ 177 ][ 349 ],
   alphaCSR[ 177 ][ 350 ],
   alphaCSR[ 177 ][ 351 ],
   alphaCSR[ 177 ][ 352 ],
   alphaCSR[ 177 ][ 353 ],
   alphaCSR[ 177 ][ 354 ],
   alphaCSR[ 177 ][ 355 ],
   alphaCSR[ 177 ][ 356 ],
   alphaCSR[ 177 ][ 357 ],
   alphaCSR[ 177 ][ 358 ],
   alphaCSR[ 177 ][ 359 ],
   alphaCSR[ 177 ][ 360 ],
   alphaCSR[ 177 ][ 361 ],
   alphaCSR[ 177 ][ 362 ],
   alphaCSR[ 177 ][ 363 ],
   alphaCSR[ 177 ][ 364 ],
   alphaCSR[ 177 ][ 365 ],
   alphaCSR[ 177 ][ 366 ],
   alphaCSR[ 177 ][ 367 ],
   alphaCSR[ 177 ][ 368 ],
   alphaCSR[ 177 ][ 369 ],
   alphaCSR[ 177 ][ 370 ],
   alphaCSR[ 177 ][ 371 ],
   alphaCSR[ 177 ][ 372 ],
   alphaCSR[ 177 ][ 373 ],
   alphaCSR[ 177 ][ 374 ],
   alphaCSR[ 177 ][ 375 ],
   alphaCSR[ 177 ][ 376 ],
   alphaCSR[ 177 ][ 377 ],
   alphaCSR[ 177 ][ 378 ],
   alphaCSR[ 177 ][ 379 ],
   alphaCSR[ 177 ][ 380 ],
   alphaCSR[ 177 ][ 381 ],
   alphaCSR[ 177 ][ 382 ],
   alphaCSR[ 177 ][ 383 ],
   alphaCSR[ 178 ][ 0 ],
   alphaCSR[ 178 ][ 1 ],
   alphaCSR[ 178 ][ 2 ],
   alphaCSR[ 178 ][ 3 ],
   alphaCSR[ 178 ][ 4 ],
   alphaCSR[ 178 ][ 5 ],
   alphaCSR[ 178 ][ 6 ],
   alphaCSR[ 178 ][ 7 ],
   alphaCSR[ 178 ][ 8 ],
   alphaCSR[ 178 ][ 9 ],
   alphaCSR[ 178 ][ 10 ],
   alphaCSR[ 178 ][ 11 ],
   alphaCSR[ 178 ][ 12 ],
   alphaCSR[ 178 ][ 13 ],
   alphaCSR[ 178 ][ 14 ],
   alphaCSR[ 178 ][ 15 ],
   alphaCSR[ 178 ][ 16 ],
   alphaCSR[ 178 ][ 17 ],
   alphaCSR[ 178 ][ 18 ],
   alphaCSR[ 178 ][ 19 ],
   alphaCSR[ 178 ][ 20 ],
   alphaCSR[ 178 ][ 21 ],
   alphaCSR[ 178 ][ 22 ],
   alphaCSR[ 178 ][ 23 ],
   alphaCSR[ 178 ][ 24 ],
   alphaCSR[ 178 ][ 25 ],
   alphaCSR[ 178 ][ 26 ],
   alphaCSR[ 178 ][ 27 ],
   alphaCSR[ 178 ][ 28 ],
   alphaCSR[ 178 ][ 29 ],
   alphaCSR[ 178 ][ 30 ],
   alphaCSR[ 178 ][ 31 ],
   alphaCSR[ 178 ][ 32 ],
   alphaCSR[ 178 ][ 33 ],
   alphaCSR[ 178 ][ 34 ],
   alphaCSR[ 178 ][ 35 ],
   alphaCSR[ 178 ][ 36 ],
   alphaCSR[ 178 ][ 37 ],
   alphaCSR[ 178 ][ 38 ],
   alphaCSR[ 178 ][ 39 ],
   alphaCSR[ 178 ][ 40 ],
   alphaCSR[ 178 ][ 41 ],
   alphaCSR[ 178 ][ 42 ],
   alphaCSR[ 178 ][ 43 ],
   alphaCSR[ 178 ][ 44 ],
   alphaCSR[ 178 ][ 45 ],
   alphaCSR[ 178 ][ 46 ],
   alphaCSR[ 178 ][ 47 ],
   alphaCSR[ 178 ][ 48 ],
   alphaCSR[ 178 ][ 49 ],
   alphaCSR[ 178 ][ 50 ],
   alphaCSR[ 178 ][ 51 ],
   alphaCSR[ 178 ][ 52 ],
   alphaCSR[ 178 ][ 53 ],
   alphaCSR[ 178 ][ 54 ],
   alphaCSR[ 178 ][ 55 ],
   alphaCSR[ 178 ][ 56 ],
   alphaCSR[ 178 ][ 57 ],
   alphaCSR[ 178 ][ 58 ],
   alphaCSR[ 178 ][ 59 ],
   alphaCSR[ 178 ][ 60 ],
   alphaCSR[ 178 ][ 61 ],
   alphaCSR[ 178 ][ 62 ],
   alphaCSR[ 178 ][ 63 ],
   alphaCSR[ 178 ][ 64 ],
   alphaCSR[ 178 ][ 65 ],
   alphaCSR[ 178 ][ 66 ],
   alphaCSR[ 178 ][ 67 ],
   alphaCSR[ 178 ][ 68 ],
   alphaCSR[ 178 ][ 69 ],
   alphaCSR[ 178 ][ 70 ],
   alphaCSR[ 178 ][ 71 ],
   alphaCSR[ 178 ][ 72 ],
   alphaCSR[ 178 ][ 73 ],
   alphaCSR[ 178 ][ 74 ],
   alphaCSR[ 178 ][ 75 ],
   alphaCSR[ 178 ][ 76 ],
   alphaCSR[ 178 ][ 77 ],
   alphaCSR[ 178 ][ 78 ],
   alphaCSR[ 178 ][ 79 ],
   alphaCSR[ 178 ][ 80 ],
   alphaCSR[ 178 ][ 81 ],
   alphaCSR[ 178 ][ 82 ],
   alphaCSR[ 178 ][ 83 ],
   alphaCSR[ 178 ][ 84 ],
   alphaCSR[ 178 ][ 85 ],
   alphaCSR[ 178 ][ 86 ],
   alphaCSR[ 178 ][ 87 ],
   alphaCSR[ 178 ][ 88 ],
   alphaCSR[ 178 ][ 89 ],
   alphaCSR[ 178 ][ 90 ],
   alphaCSR[ 178 ][ 91 ],
   alphaCSR[ 178 ][ 92 ],
   alphaCSR[ 178 ][ 93 ],
   alphaCSR[ 178 ][ 94 ],
   alphaCSR[ 178 ][ 95 ],
   alphaCSR[ 178 ][ 96 ],
   alphaCSR[ 178 ][ 97 ],
   alphaCSR[ 178 ][ 98 ],
   alphaCSR[ 178 ][ 99 ],
   alphaCSR[ 178 ][ 100 ],
   alphaCSR[ 178 ][ 101 ],
   alphaCSR[ 178 ][ 102 ],
   alphaCSR[ 178 ][ 103 ],
   alphaCSR[ 178 ][ 104 ],
   alphaCSR[ 178 ][ 105 ],
   alphaCSR[ 178 ][ 106 ],
   alphaCSR[ 178 ][ 107 ],
   alphaCSR[ 178 ][ 108 ],
   alphaCSR[ 178 ][ 109 ],
   alphaCSR[ 178 ][ 110 ],
   alphaCSR[ 178 ][ 111 ],
   alphaCSR[ 178 ][ 112 ],
   alphaCSR[ 178 ][ 113 ],
   alphaCSR[ 178 ][ 114 ],
   alphaCSR[ 178 ][ 115 ],
   alphaCSR[ 178 ][ 116 ],
   alphaCSR[ 178 ][ 117 ],
   alphaCSR[ 178 ][ 118 ],
   alphaCSR[ 178 ][ 119 ],
   alphaCSR[ 178 ][ 120 ],
   alphaCSR[ 178 ][ 121 ],
   alphaCSR[ 178 ][ 122 ],
   alphaCSR[ 178 ][ 123 ],
   alphaCSR[ 178 ][ 124 ],
   alphaCSR[ 178 ][ 125 ],
   alphaCSR[ 178 ][ 126 ],
   alphaCSR[ 178 ][ 127 ],
   alphaCSR[ 178 ][ 128 ],
   alphaCSR[ 178 ][ 129 ],
   alphaCSR[ 178 ][ 130 ],
   alphaCSR[ 178 ][ 131 ],
   alphaCSR[ 178 ][ 132 ],
   alphaCSR[ 178 ][ 133 ],
   alphaCSR[ 178 ][ 134 ],
   alphaCSR[ 178 ][ 135 ],
   alphaCSR[ 178 ][ 136 ],
   alphaCSR[ 178 ][ 137 ],
   alphaCSR[ 178 ][ 138 ],
   alphaCSR[ 178 ][ 139 ],
   alphaCSR[ 178 ][ 140 ],
   alphaCSR[ 178 ][ 141 ],
   alphaCSR[ 178 ][ 142 ],
   alphaCSR[ 178 ][ 143 ],
   alphaCSR[ 178 ][ 144 ],
   alphaCSR[ 178 ][ 145 ],
   alphaCSR[ 178 ][ 146 ],
   alphaCSR[ 178 ][ 147 ],
   alphaCSR[ 178 ][ 148 ],
   alphaCSR[ 178 ][ 149 ],
   alphaCSR[ 178 ][ 150 ],
   alphaCSR[ 178 ][ 151 ],
   alphaCSR[ 178 ][ 152 ],
   alphaCSR[ 178 ][ 153 ],
   alphaCSR[ 178 ][ 154 ],
   alphaCSR[ 178 ][ 155 ],
   alphaCSR[ 178 ][ 156 ],
   alphaCSR[ 178 ][ 157 ],
   alphaCSR[ 178 ][ 158 ],
   alphaCSR[ 178 ][ 159 ],
   alphaCSR[ 178 ][ 160 ],
   alphaCSR[ 178 ][ 161 ],
   alphaCSR[ 178 ][ 162 ],
   alphaCSR[ 178 ][ 163 ],
   alphaCSR[ 178 ][ 164 ],
   alphaCSR[ 178 ][ 165 ],
   alphaCSR[ 178 ][ 166 ],
   alphaCSR[ 178 ][ 167 ],
   alphaCSR[ 178 ][ 168 ],
   alphaCSR[ 178 ][ 169 ],
   alphaCSR[ 178 ][ 170 ],
   alphaCSR[ 178 ][ 171 ],
   alphaCSR[ 178 ][ 172 ],
   alphaCSR[ 178 ][ 173 ],
   alphaCSR[ 178 ][ 174 ],
   alphaCSR[ 178 ][ 175 ],
   alphaCSR[ 178 ][ 176 ],
   alphaCSR[ 178 ][ 177 ],
   alphaCSR[ 178 ][ 178 ],
   alphaCSR[ 178 ][ 179 ],
   alphaCSR[ 178 ][ 180 ],
   alphaCSR[ 178 ][ 181 ],
   alphaCSR[ 178 ][ 182 ],
   alphaCSR[ 178 ][ 183 ],
   alphaCSR[ 178 ][ 184 ],
   alphaCSR[ 178 ][ 185 ],
   alphaCSR[ 178 ][ 186 ],
   alphaCSR[ 178 ][ 187 ],
   alphaCSR[ 178 ][ 188 ],
   alphaCSR[ 178 ][ 189 ],
   alphaCSR[ 178 ][ 190 ],
   alphaCSR[ 178 ][ 191 ],
   alphaCSR[ 178 ][ 192 ],
   alphaCSR[ 178 ][ 193 ],
   alphaCSR[ 178 ][ 194 ],
   alphaCSR[ 178 ][ 195 ],
   alphaCSR[ 178 ][ 196 ],
   alphaCSR[ 178 ][ 197 ],
   alphaCSR[ 178 ][ 198 ],
   alphaCSR[ 178 ][ 199 ],
   alphaCSR[ 178 ][ 200 ],
   alphaCSR[ 178 ][ 201 ],
   alphaCSR[ 178 ][ 202 ],
   alphaCSR[ 178 ][ 203 ],
   alphaCSR[ 178 ][ 204 ],
   alphaCSR[ 178 ][ 205 ],
   alphaCSR[ 178 ][ 206 ],
   alphaCSR[ 178 ][ 207 ],
   alphaCSR[ 178 ][ 208 ],
   alphaCSR[ 178 ][ 209 ],
   alphaCSR[ 178 ][ 210 ],
   alphaCSR[ 178 ][ 211 ],
   alphaCSR[ 178 ][ 212 ],
   alphaCSR[ 178 ][ 213 ],
   alphaCSR[ 178 ][ 214 ],
   alphaCSR[ 178 ][ 215 ],
   alphaCSR[ 178 ][ 216 ],
   alphaCSR[ 178 ][ 217 ],
   alphaCSR[ 178 ][ 218 ],
   alphaCSR[ 178 ][ 219 ],
   alphaCSR[ 178 ][ 220 ],
   alphaCSR[ 178 ][ 221 ],
   alphaCSR[ 178 ][ 222 ],
   alphaCSR[ 178 ][ 223 ],
   alphaCSR[ 178 ][ 224 ],
   alphaCSR[ 178 ][ 225 ],
   alphaCSR[ 178 ][ 226 ],
   alphaCSR[ 178 ][ 227 ],
   alphaCSR[ 178 ][ 228 ],
   alphaCSR[ 178 ][ 229 ],
   alphaCSR[ 178 ][ 230 ],
   alphaCSR[ 178 ][ 231 ],
   alphaCSR[ 178 ][ 232 ],
   alphaCSR[ 178 ][ 233 ],
   alphaCSR[ 178 ][ 234 ],
   alphaCSR[ 178 ][ 235 ],
   alphaCSR[ 178 ][ 236 ],
   alphaCSR[ 178 ][ 237 ],
   alphaCSR[ 178 ][ 238 ],
   alphaCSR[ 178 ][ 239 ],
   alphaCSR[ 178 ][ 240 ],
   alphaCSR[ 178 ][ 241 ],
   alphaCSR[ 178 ][ 242 ],
   alphaCSR[ 178 ][ 243 ],
   alphaCSR[ 178 ][ 244 ],
   alphaCSR[ 178 ][ 245 ],
   alphaCSR[ 178 ][ 246 ],
   alphaCSR[ 178 ][ 247 ],
   alphaCSR[ 178 ][ 248 ],
   alphaCSR[ 178 ][ 249 ],
   alphaCSR[ 178 ][ 250 ],
   alphaCSR[ 178 ][ 251 ],
   alphaCSR[ 178 ][ 252 ],
   alphaCSR[ 178 ][ 253 ],
   alphaCSR[ 178 ][ 254 ],
   alphaCSR[ 178 ][ 255 ],
   alphaCSR[ 178 ][ 256 ],
   alphaCSR[ 178 ][ 257 ],
   alphaCSR[ 178 ][ 258 ],
   alphaCSR[ 178 ][ 259 ],
   alphaCSR[ 178 ][ 260 ],
   alphaCSR[ 178 ][ 261 ],
   alphaCSR[ 178 ][ 262 ],
   alphaCSR[ 178 ][ 263 ],
   alphaCSR[ 178 ][ 264 ],
   alphaCSR[ 178 ][ 265 ],
   alphaCSR[ 178 ][ 266 ],
   alphaCSR[ 178 ][ 267 ],
   alphaCSR[ 178 ][ 268 ],
   alphaCSR[ 178 ][ 269 ],
   alphaCSR[ 178 ][ 270 ],
   alphaCSR[ 178 ][ 271 ],
   alphaCSR[ 178 ][ 272 ],
   alphaCSR[ 178 ][ 273 ],
   alphaCSR[ 178 ][ 274 ],
   alphaCSR[ 178 ][ 275 ],
   alphaCSR[ 178 ][ 276 ],
   alphaCSR[ 178 ][ 277 ],
   alphaCSR[ 178 ][ 278 ],
   alphaCSR[ 178 ][ 279 ],
   alphaCSR[ 178 ][ 280 ],
   alphaCSR[ 178 ][ 281 ],
   alphaCSR[ 178 ][ 282 ],
   alphaCSR[ 178 ][ 283 ],
   alphaCSR[ 178 ][ 284 ],
   alphaCSR[ 178 ][ 285 ],
   alphaCSR[ 178 ][ 286 ],
   alphaCSR[ 178 ][ 287 ],
   alphaCSR[ 178 ][ 288 ],
   alphaCSR[ 178 ][ 289 ],
   alphaCSR[ 178 ][ 290 ],
   alphaCSR[ 178 ][ 291 ],
   alphaCSR[ 178 ][ 292 ],
   alphaCSR[ 178 ][ 293 ],
   alphaCSR[ 178 ][ 294 ],
   alphaCSR[ 178 ][ 295 ],
   alphaCSR[ 178 ][ 296 ],
   alphaCSR[ 178 ][ 297 ],
   alphaCSR[ 178 ][ 298 ],
   alphaCSR[ 178 ][ 299 ],
   alphaCSR[ 178 ][ 300 ],
   alphaCSR[ 178 ][ 301 ],
   alphaCSR[ 178 ][ 302 ],
   alphaCSR[ 178 ][ 303 ],
   alphaCSR[ 178 ][ 304 ],
   alphaCSR[ 178 ][ 305 ],
   alphaCSR[ 178 ][ 306 ],
   alphaCSR[ 178 ][ 307 ],
   alphaCSR[ 178 ][ 308 ],
   alphaCSR[ 178 ][ 309 ],
   alphaCSR[ 178 ][ 310 ],
   alphaCSR[ 178 ][ 311 ],
   alphaCSR[ 178 ][ 312 ],
   alphaCSR[ 178 ][ 313 ],
   alphaCSR[ 178 ][ 314 ],
   alphaCSR[ 178 ][ 315 ],
   alphaCSR[ 178 ][ 316 ],
   alphaCSR[ 178 ][ 317 ],
   alphaCSR[ 178 ][ 318 ],
   alphaCSR[ 178 ][ 319 ],
   alphaCSR[ 178 ][ 320 ],
   alphaCSR[ 178 ][ 321 ],
   alphaCSR[ 178 ][ 322 ],
   alphaCSR[ 178 ][ 323 ],
   alphaCSR[ 178 ][ 324 ],
   alphaCSR[ 178 ][ 325 ],
   alphaCSR[ 178 ][ 326 ],
   alphaCSR[ 178 ][ 327 ],
   alphaCSR[ 178 ][ 328 ],
   alphaCSR[ 178 ][ 329 ],
   alphaCSR[ 178 ][ 330 ],
   alphaCSR[ 178 ][ 331 ],
   alphaCSR[ 178 ][ 332 ],
   alphaCSR[ 178 ][ 333 ],
   alphaCSR[ 178 ][ 334 ],
   alphaCSR[ 178 ][ 335 ],
   alphaCSR[ 178 ][ 336 ],
   alphaCSR[ 178 ][ 337 ],
   alphaCSR[ 178 ][ 338 ],
   alphaCSR[ 178 ][ 339 ],
   alphaCSR[ 178 ][ 340 ],
   alphaCSR[ 178 ][ 341 ],
   alphaCSR[ 178 ][ 342 ],
   alphaCSR[ 178 ][ 343 ],
   alphaCSR[ 178 ][ 344 ],
   alphaCSR[ 178 ][ 345 ],
   alphaCSR[ 178 ][ 346 ],
   alphaCSR[ 178 ][ 347 ],
   alphaCSR[ 178 ][ 348 ],
   alphaCSR[ 178 ][ 349 ],
   alphaCSR[ 178 ][ 350 ],
   alphaCSR[ 178 ][ 351 ],
   alphaCSR[ 178 ][ 352 ],
   alphaCSR[ 178 ][ 353 ],
   alphaCSR[ 178 ][ 354 ],
   alphaCSR[ 178 ][ 355 ],
   alphaCSR[ 178 ][ 356 ],
   alphaCSR[ 178 ][ 357 ],
   alphaCSR[ 178 ][ 358 ],
   alphaCSR[ 178 ][ 359 ],
   alphaCSR[ 178 ][ 360 ],
   alphaCSR[ 178 ][ 361 ],
   alphaCSR[ 178 ][ 362 ],
   alphaCSR[ 178 ][ 363 ],
   alphaCSR[ 178 ][ 364 ],
   alphaCSR[ 178 ][ 365 ],
   alphaCSR[ 178 ][ 366 ],
   alphaCSR[ 178 ][ 367 ],
   alphaCSR[ 178 ][ 368 ],
   alphaCSR[ 178 ][ 369 ],
   alphaCSR[ 178 ][ 370 ],
   alphaCSR[ 178 ][ 371 ],
   alphaCSR[ 178 ][ 372 ],
   alphaCSR[ 178 ][ 373 ],
   alphaCSR[ 178 ][ 374 ],
   alphaCSR[ 178 ][ 375 ],
   alphaCSR[ 178 ][ 376 ],
   alphaCSR[ 178 ][ 377 ],
   alphaCSR[ 178 ][ 378 ],
   alphaCSR[ 178 ][ 379 ],
   alphaCSR[ 178 ][ 380 ],
   alphaCSR[ 178 ][ 381 ],
   alphaCSR[ 178 ][ 382 ],
   alphaCSR[ 178 ][ 383 ],
   alphaCSR[ 179 ][ 0 ],
   alphaCSR[ 179 ][ 1 ],
   alphaCSR[ 179 ][ 2 ],
   alphaCSR[ 179 ][ 3 ],
   alphaCSR[ 179 ][ 4 ],
   alphaCSR[ 179 ][ 5 ],
   alphaCSR[ 179 ][ 6 ],
   alphaCSR[ 179 ][ 7 ],
   alphaCSR[ 179 ][ 8 ],
   alphaCSR[ 179 ][ 9 ],
   alphaCSR[ 179 ][ 10 ],
   alphaCSR[ 179 ][ 11 ],
   alphaCSR[ 179 ][ 12 ],
   alphaCSR[ 179 ][ 13 ],
   alphaCSR[ 179 ][ 14 ],
   alphaCSR[ 179 ][ 15 ],
   alphaCSR[ 179 ][ 16 ],
   alphaCSR[ 179 ][ 17 ],
   alphaCSR[ 179 ][ 18 ],
   alphaCSR[ 179 ][ 19 ],
   alphaCSR[ 179 ][ 20 ],
   alphaCSR[ 179 ][ 21 ],
   alphaCSR[ 179 ][ 22 ],
   alphaCSR[ 179 ][ 23 ],
   alphaCSR[ 179 ][ 24 ],
   alphaCSR[ 179 ][ 25 ],
   alphaCSR[ 179 ][ 26 ],
   alphaCSR[ 179 ][ 27 ],
   alphaCSR[ 179 ][ 28 ],
   alphaCSR[ 179 ][ 29 ],
   alphaCSR[ 179 ][ 30 ],
   alphaCSR[ 179 ][ 31 ],
   alphaCSR[ 179 ][ 32 ],
   alphaCSR[ 179 ][ 33 ],
   alphaCSR[ 179 ][ 34 ],
   alphaCSR[ 179 ][ 35 ],
   alphaCSR[ 179 ][ 36 ],
   alphaCSR[ 179 ][ 37 ],
   alphaCSR[ 179 ][ 38 ],
   alphaCSR[ 179 ][ 39 ],
   alphaCSR[ 179 ][ 40 ],
   alphaCSR[ 179 ][ 41 ],
   alphaCSR[ 179 ][ 42 ],
   alphaCSR[ 179 ][ 43 ],
   alphaCSR[ 179 ][ 44 ],
   alphaCSR[ 179 ][ 45 ],
   alphaCSR[ 179 ][ 46 ],
   alphaCSR[ 179 ][ 47 ],
   alphaCSR[ 179 ][ 48 ],
   alphaCSR[ 179 ][ 49 ],
   alphaCSR[ 179 ][ 50 ],
   alphaCSR[ 179 ][ 51 ],
   alphaCSR[ 179 ][ 52 ],
   alphaCSR[ 179 ][ 53 ],
   alphaCSR[ 179 ][ 54 ],
   alphaCSR[ 179 ][ 55 ],
   alphaCSR[ 179 ][ 56 ],
   alphaCSR[ 179 ][ 57 ],
   alphaCSR[ 179 ][ 58 ],
   alphaCSR[ 179 ][ 59 ],
   alphaCSR[ 179 ][ 60 ],
   alphaCSR[ 179 ][ 61 ],
   alphaCSR[ 179 ][ 62 ],
   alphaCSR[ 179 ][ 63 ],
   alphaCSR[ 179 ][ 64 ],
   alphaCSR[ 179 ][ 65 ],
   alphaCSR[ 179 ][ 66 ],
   alphaCSR[ 179 ][ 67 ],
   alphaCSR[ 179 ][ 68 ],
   alphaCSR[ 179 ][ 69 ],
   alphaCSR[ 179 ][ 70 ],
   alphaCSR[ 179 ][ 71 ],
   alphaCSR[ 179 ][ 72 ],
   alphaCSR[ 179 ][ 73 ],
   alphaCSR[ 179 ][ 74 ],
   alphaCSR[ 179 ][ 75 ],
   alphaCSR[ 179 ][ 76 ],
   alphaCSR[ 179 ][ 77 ],
   alphaCSR[ 179 ][ 78 ],
   alphaCSR[ 179 ][ 79 ],
   alphaCSR[ 179 ][ 80 ],
   alphaCSR[ 179 ][ 81 ],
   alphaCSR[ 179 ][ 82 ],
   alphaCSR[ 179 ][ 83 ],
   alphaCSR[ 179 ][ 84 ],
   alphaCSR[ 179 ][ 85 ],
   alphaCSR[ 179 ][ 86 ],
   alphaCSR[ 179 ][ 87 ],
   alphaCSR[ 179 ][ 88 ],
   alphaCSR[ 179 ][ 89 ],
   alphaCSR[ 179 ][ 90 ],
   alphaCSR[ 179 ][ 91 ],
   alphaCSR[ 179 ][ 92 ],
   alphaCSR[ 179 ][ 93 ],
   alphaCSR[ 179 ][ 94 ],
   alphaCSR[ 179 ][ 95 ],
   alphaCSR[ 179 ][ 96 ],
   alphaCSR[ 179 ][ 97 ],
   alphaCSR[ 179 ][ 98 ],
   alphaCSR[ 179 ][ 99 ],
   alphaCSR[ 179 ][ 100 ],
   alphaCSR[ 179 ][ 101 ],
   alphaCSR[ 179 ][ 102 ],
   alphaCSR[ 179 ][ 103 ],
   alphaCSR[ 179 ][ 104 ],
   alphaCSR[ 179 ][ 105 ],
   alphaCSR[ 179 ][ 106 ],
   alphaCSR[ 179 ][ 107 ],
   alphaCSR[ 179 ][ 108 ],
   alphaCSR[ 179 ][ 109 ],
   alphaCSR[ 179 ][ 110 ],
   alphaCSR[ 179 ][ 111 ],
   alphaCSR[ 179 ][ 112 ],
   alphaCSR[ 179 ][ 113 ],
   alphaCSR[ 179 ][ 114 ],
   alphaCSR[ 179 ][ 115 ],
   alphaCSR[ 179 ][ 116 ],
   alphaCSR[ 179 ][ 117 ],
   alphaCSR[ 179 ][ 118 ],
   alphaCSR[ 179 ][ 119 ],
   alphaCSR[ 179 ][ 120 ],
   alphaCSR[ 179 ][ 121 ],
   alphaCSR[ 179 ][ 122 ],
   alphaCSR[ 179 ][ 123 ],
   alphaCSR[ 179 ][ 124 ],
   alphaCSR[ 179 ][ 125 ],
   alphaCSR[ 179 ][ 126 ],
   alphaCSR[ 179 ][ 127 ],
   alphaCSR[ 179 ][ 128 ],
   alphaCSR[ 179 ][ 129 ],
   alphaCSR[ 179 ][ 130 ],
   alphaCSR[ 179 ][ 131 ],
   alphaCSR[ 179 ][ 132 ],
   alphaCSR[ 179 ][ 133 ],
   alphaCSR[ 179 ][ 134 ],
   alphaCSR[ 179 ][ 135 ],
   alphaCSR[ 179 ][ 136 ],
   alphaCSR[ 179 ][ 137 ],
   alphaCSR[ 179 ][ 138 ],
   alphaCSR[ 179 ][ 139 ],
   alphaCSR[ 179 ][ 140 ],
   alphaCSR[ 179 ][ 141 ],
   alphaCSR[ 179 ][ 142 ],
   alphaCSR[ 179 ][ 143 ],
   alphaCSR[ 179 ][ 144 ],
   alphaCSR[ 179 ][ 145 ],
   alphaCSR[ 179 ][ 146 ],
   alphaCSR[ 179 ][ 147 ],
   alphaCSR[ 179 ][ 148 ],
   alphaCSR[ 179 ][ 149 ],
   alphaCSR[ 179 ][ 150 ],
   alphaCSR[ 179 ][ 151 ],
   alphaCSR[ 179 ][ 152 ],
   alphaCSR[ 179 ][ 153 ],
   alphaCSR[ 179 ][ 154 ],
   alphaCSR[ 179 ][ 155 ],
   alphaCSR[ 179 ][ 156 ],
   alphaCSR[ 179 ][ 157 ],
   alphaCSR[ 179 ][ 158 ],
   alphaCSR[ 179 ][ 159 ],
   alphaCSR[ 179 ][ 160 ],
   alphaCSR[ 179 ][ 161 ],
   alphaCSR[ 179 ][ 162 ],
   alphaCSR[ 179 ][ 163 ],
   alphaCSR[ 179 ][ 164 ],
   alphaCSR[ 179 ][ 165 ],
   alphaCSR[ 179 ][ 166 ],
   alphaCSR[ 179 ][ 167 ],
   alphaCSR[ 179 ][ 168 ],
   alphaCSR[ 179 ][ 169 ],
   alphaCSR[ 179 ][ 170 ],
   alphaCSR[ 179 ][ 171 ],
   alphaCSR[ 179 ][ 172 ],
   alphaCSR[ 179 ][ 173 ],
   alphaCSR[ 179 ][ 174 ],
   alphaCSR[ 179 ][ 175 ],
   alphaCSR[ 179 ][ 176 ],
   alphaCSR[ 179 ][ 177 ],
   alphaCSR[ 179 ][ 178 ],
   alphaCSR[ 179 ][ 179 ],
   alphaCSR[ 179 ][ 180 ],
   alphaCSR[ 179 ][ 181 ],
   alphaCSR[ 179 ][ 182 ],
   alphaCSR[ 179 ][ 183 ],
   alphaCSR[ 179 ][ 184 ],
   alphaCSR[ 179 ][ 185 ],
   alphaCSR[ 179 ][ 186 ],
   alphaCSR[ 179 ][ 187 ],
   alphaCSR[ 179 ][ 188 ],
   alphaCSR[ 179 ][ 189 ],
   alphaCSR[ 179 ][ 190 ],
   alphaCSR[ 179 ][ 191 ],
   alphaCSR[ 179 ][ 192 ],
   alphaCSR[ 179 ][ 193 ],
   alphaCSR[ 179 ][ 194 ],
   alphaCSR[ 179 ][ 195 ],
   alphaCSR[ 179 ][ 196 ],
   alphaCSR[ 179 ][ 197 ],
   alphaCSR[ 179 ][ 198 ],
   alphaCSR[ 179 ][ 199 ],
   alphaCSR[ 179 ][ 200 ],
   alphaCSR[ 179 ][ 201 ],
   alphaCSR[ 179 ][ 202 ],
   alphaCSR[ 179 ][ 203 ],
   alphaCSR[ 179 ][ 204 ],
   alphaCSR[ 179 ][ 205 ],
   alphaCSR[ 179 ][ 206 ],
   alphaCSR[ 179 ][ 207 ],
   alphaCSR[ 179 ][ 208 ],
   alphaCSR[ 179 ][ 209 ],
   alphaCSR[ 179 ][ 210 ],
   alphaCSR[ 179 ][ 211 ],
   alphaCSR[ 179 ][ 212 ],
   alphaCSR[ 179 ][ 213 ],
   alphaCSR[ 179 ][ 214 ],
   alphaCSR[ 179 ][ 215 ],
   alphaCSR[ 179 ][ 216 ],
   alphaCSR[ 179 ][ 217 ],
   alphaCSR[ 179 ][ 218 ],
   alphaCSR[ 179 ][ 219 ],
   alphaCSR[ 179 ][ 220 ],
   alphaCSR[ 179 ][ 221 ],
   alphaCSR[ 179 ][ 222 ],
   alphaCSR[ 179 ][ 223 ],
   alphaCSR[ 179 ][ 224 ],
   alphaCSR[ 179 ][ 225 ],
   alphaCSR[ 179 ][ 226 ],
   alphaCSR[ 179 ][ 227 ],
   alphaCSR[ 179 ][ 228 ],
   alphaCSR[ 179 ][ 229 ],
   alphaCSR[ 179 ][ 230 ],
   alphaCSR[ 179 ][ 231 ],
   alphaCSR[ 179 ][ 232 ],
   alphaCSR[ 179 ][ 233 ],
   alphaCSR[ 179 ][ 234 ],
   alphaCSR[ 179 ][ 235 ],
   alphaCSR[ 179 ][ 236 ],
   alphaCSR[ 179 ][ 237 ],
   alphaCSR[ 179 ][ 238 ],
   alphaCSR[ 179 ][ 239 ],
   alphaCSR[ 179 ][ 240 ],
   alphaCSR[ 179 ][ 241 ],
   alphaCSR[ 179 ][ 242 ],
   alphaCSR[ 179 ][ 243 ],
   alphaCSR[ 179 ][ 244 ],
   alphaCSR[ 179 ][ 245 ],
   alphaCSR[ 179 ][ 246 ],
   alphaCSR[ 179 ][ 247 ],
   alphaCSR[ 179 ][ 248 ],
   alphaCSR[ 179 ][ 249 ],
   alphaCSR[ 179 ][ 250 ],
   alphaCSR[ 179 ][ 251 ],
   alphaCSR[ 179 ][ 252 ],
   alphaCSR[ 179 ][ 253 ],
   alphaCSR[ 179 ][ 254 ],
   alphaCSR[ 179 ][ 255 ],
   alphaCSR[ 179 ][ 256 ],
   alphaCSR[ 179 ][ 257 ],
   alphaCSR[ 179 ][ 258 ],
   alphaCSR[ 179 ][ 259 ],
   alphaCSR[ 179 ][ 260 ],
   alphaCSR[ 179 ][ 261 ],
   alphaCSR[ 179 ][ 262 ],
   alphaCSR[ 179 ][ 263 ],
   alphaCSR[ 179 ][ 264 ],
   alphaCSR[ 179 ][ 265 ],
   alphaCSR[ 179 ][ 266 ],
   alphaCSR[ 179 ][ 267 ],
   alphaCSR[ 179 ][ 268 ],
   alphaCSR[ 179 ][ 269 ],
   alphaCSR[ 179 ][ 270 ],
   alphaCSR[ 179 ][ 271 ],
   alphaCSR[ 179 ][ 272 ],
   alphaCSR[ 179 ][ 273 ],
   alphaCSR[ 179 ][ 274 ],
   alphaCSR[ 179 ][ 275 ],
   alphaCSR[ 179 ][ 276 ],
   alphaCSR[ 179 ][ 277 ],
   alphaCSR[ 179 ][ 278 ],
   alphaCSR[ 179 ][ 279 ],
   alphaCSR[ 179 ][ 280 ],
   alphaCSR[ 179 ][ 281 ],
   alphaCSR[ 179 ][ 282 ],
   alphaCSR[ 179 ][ 283 ],
   alphaCSR[ 179 ][ 284 ],
   alphaCSR[ 179 ][ 285 ],
   alphaCSR[ 179 ][ 286 ],
   alphaCSR[ 179 ][ 287 ],
   alphaCSR[ 179 ][ 288 ],
   alphaCSR[ 179 ][ 289 ],
   alphaCSR[ 179 ][ 290 ],
   alphaCSR[ 179 ][ 291 ],
   alphaCSR[ 179 ][ 292 ],
   alphaCSR[ 179 ][ 293 ],
   alphaCSR[ 179 ][ 294 ],
   alphaCSR[ 179 ][ 295 ],
   alphaCSR[ 179 ][ 296 ],
   alphaCSR[ 179 ][ 297 ],
   alphaCSR[ 179 ][ 298 ],
   alphaCSR[ 179 ][ 299 ],
   alphaCSR[ 179 ][ 300 ],
   alphaCSR[ 179 ][ 301 ],
   alphaCSR[ 179 ][ 302 ],
   alphaCSR[ 179 ][ 303 ],
   alphaCSR[ 179 ][ 304 ],
   alphaCSR[ 179 ][ 305 ],
   alphaCSR[ 179 ][ 306 ],
   alphaCSR[ 179 ][ 307 ],
   alphaCSR[ 179 ][ 308 ],
   alphaCSR[ 179 ][ 309 ],
   alphaCSR[ 179 ][ 310 ],
   alphaCSR[ 179 ][ 311 ],
   alphaCSR[ 179 ][ 312 ],
   alphaCSR[ 179 ][ 313 ],
   alphaCSR[ 179 ][ 314 ],
   alphaCSR[ 179 ][ 315 ],
   alphaCSR[ 179 ][ 316 ],
   alphaCSR[ 179 ][ 317 ],
   alphaCSR[ 179 ][ 318 ],
   alphaCSR[ 179 ][ 319 ],
   alphaCSR[ 179 ][ 320 ],
   alphaCSR[ 179 ][ 321 ],
   alphaCSR[ 179 ][ 322 ],
   alphaCSR[ 179 ][ 323 ],
   alphaCSR[ 179 ][ 324 ],
   alphaCSR[ 179 ][ 325 ],
   alphaCSR[ 179 ][ 326 ],
   alphaCSR[ 179 ][ 327 ],
   alphaCSR[ 179 ][ 328 ],
   alphaCSR[ 179 ][ 329 ],
   alphaCSR[ 179 ][ 330 ],
   alphaCSR[ 179 ][ 331 ],
   alphaCSR[ 179 ][ 332 ],
   alphaCSR[ 179 ][ 333 ],
   alphaCSR[ 179 ][ 334 ],
   alphaCSR[ 179 ][ 335 ],
   alphaCSR[ 179 ][ 336 ],
   alphaCSR[ 179 ][ 337 ],
   alphaCSR[ 179 ][ 338 ],
   alphaCSR[ 179 ][ 339 ],
   alphaCSR[ 179 ][ 340 ],
   alphaCSR[ 179 ][ 341 ],
   alphaCSR[ 179 ][ 342 ],
   alphaCSR[ 179 ][ 343 ],
   alphaCSR[ 179 ][ 344 ],
   alphaCSR[ 179 ][ 345 ],
   alphaCSR[ 179 ][ 346 ],
   alphaCSR[ 179 ][ 347 ],
   alphaCSR[ 179 ][ 348 ],
   alphaCSR[ 179 ][ 349 ],
   alphaCSR[ 179 ][ 350 ],
   alphaCSR[ 179 ][ 351 ],
   alphaCSR[ 179 ][ 352 ],
   alphaCSR[ 179 ][ 353 ],
   alphaCSR[ 179 ][ 354 ],
   alphaCSR[ 179 ][ 355 ],
   alphaCSR[ 179 ][ 356 ],
   alphaCSR[ 179 ][ 357 ],
   alphaCSR[ 179 ][ 358 ],
   alphaCSR[ 179 ][ 359 ],
   alphaCSR[ 179 ][ 360 ],
   alphaCSR[ 179 ][ 361 ],
   alphaCSR[ 179 ][ 362 ],
   alphaCSR[ 179 ][ 363 ],
   alphaCSR[ 179 ][ 364 ],
   alphaCSR[ 179 ][ 365 ],
   alphaCSR[ 179 ][ 366 ],
   alphaCSR[ 179 ][ 367 ],
   alphaCSR[ 179 ][ 368 ],
   alphaCSR[ 179 ][ 369 ],
   alphaCSR[ 179 ][ 370 ],
   alphaCSR[ 179 ][ 371 ],
   alphaCSR[ 179 ][ 372 ],
   alphaCSR[ 179 ][ 373 ],
   alphaCSR[ 179 ][ 374 ],
   alphaCSR[ 179 ][ 375 ],
   alphaCSR[ 179 ][ 376 ],
   alphaCSR[ 179 ][ 377 ],
   alphaCSR[ 179 ][ 378 ],
   alphaCSR[ 179 ][ 379 ],
   alphaCSR[ 179 ][ 380 ],
   alphaCSR[ 179 ][ 381 ],
   alphaCSR[ 179 ][ 382 ],
   alphaCSR[ 179 ][ 383 ],
   alphaCSR[ 180 ][ 0 ],
   alphaCSR[ 180 ][ 1 ],
   alphaCSR[ 180 ][ 2 ],
   alphaCSR[ 180 ][ 3 ],
   alphaCSR[ 180 ][ 4 ],
   alphaCSR[ 180 ][ 5 ],
   alphaCSR[ 180 ][ 6 ],
   alphaCSR[ 180 ][ 7 ],
   alphaCSR[ 180 ][ 8 ],
   alphaCSR[ 180 ][ 9 ],
   alphaCSR[ 180 ][ 10 ],
   alphaCSR[ 180 ][ 11 ],
   alphaCSR[ 180 ][ 12 ],
   alphaCSR[ 180 ][ 13 ],
   alphaCSR[ 180 ][ 14 ],
   alphaCSR[ 180 ][ 15 ],
   alphaCSR[ 180 ][ 16 ],
   alphaCSR[ 180 ][ 17 ],
   alphaCSR[ 180 ][ 18 ],
   alphaCSR[ 180 ][ 19 ],
   alphaCSR[ 180 ][ 20 ],
   alphaCSR[ 180 ][ 21 ],
   alphaCSR[ 180 ][ 22 ],
   alphaCSR[ 180 ][ 23 ],
   alphaCSR[ 180 ][ 24 ],
   alphaCSR[ 180 ][ 25 ],
   alphaCSR[ 180 ][ 26 ],
   alphaCSR[ 180 ][ 27 ],
   alphaCSR[ 180 ][ 28 ],
   alphaCSR[ 180 ][ 29 ],
   alphaCSR[ 180 ][ 30 ],
   alphaCSR[ 180 ][ 31 ],
   alphaCSR[ 180 ][ 32 ],
   alphaCSR[ 180 ][ 33 ],
   alphaCSR[ 180 ][ 34 ],
   alphaCSR[ 180 ][ 35 ],
   alphaCSR[ 180 ][ 36 ],
   alphaCSR[ 180 ][ 37 ],
   alphaCSR[ 180 ][ 38 ],
   alphaCSR[ 180 ][ 39 ],
   alphaCSR[ 180 ][ 40 ],
   alphaCSR[ 180 ][ 41 ],
   alphaCSR[ 180 ][ 42 ],
   alphaCSR[ 180 ][ 43 ],
   alphaCSR[ 180 ][ 44 ],
   alphaCSR[ 180 ][ 45 ],
   alphaCSR[ 180 ][ 46 ],
   alphaCSR[ 180 ][ 47 ],
   alphaCSR[ 180 ][ 48 ],
   alphaCSR[ 180 ][ 49 ],
   alphaCSR[ 180 ][ 50 ],
   alphaCSR[ 180 ][ 51 ],
   alphaCSR[ 180 ][ 52 ],
   alphaCSR[ 180 ][ 53 ],
   alphaCSR[ 180 ][ 54 ],
   alphaCSR[ 180 ][ 55 ],
   alphaCSR[ 180 ][ 56 ],
   alphaCSR[ 180 ][ 57 ],
   alphaCSR[ 180 ][ 58 ],
   alphaCSR[ 180 ][ 59 ],
   alphaCSR[ 180 ][ 60 ],
   alphaCSR[ 180 ][ 61 ],
   alphaCSR[ 180 ][ 62 ],
   alphaCSR[ 180 ][ 63 ],
   alphaCSR[ 180 ][ 64 ],
   alphaCSR[ 180 ][ 65 ],
   alphaCSR[ 180 ][ 66 ],
   alphaCSR[ 180 ][ 67 ],
   alphaCSR[ 180 ][ 68 ],
   alphaCSR[ 180 ][ 69 ],
   alphaCSR[ 180 ][ 70 ],
   alphaCSR[ 180 ][ 71 ],
   alphaCSR[ 180 ][ 72 ],
   alphaCSR[ 180 ][ 73 ],
   alphaCSR[ 180 ][ 74 ],
   alphaCSR[ 180 ][ 75 ],
   alphaCSR[ 180 ][ 76 ],
   alphaCSR[ 180 ][ 77 ],
   alphaCSR[ 180 ][ 78 ],
   alphaCSR[ 180 ][ 79 ],
   alphaCSR[ 180 ][ 80 ],
   alphaCSR[ 180 ][ 81 ],
   alphaCSR[ 180 ][ 82 ],
   alphaCSR[ 180 ][ 83 ],
   alphaCSR[ 180 ][ 84 ],
   alphaCSR[ 180 ][ 85 ],
   alphaCSR[ 180 ][ 86 ],
   alphaCSR[ 180 ][ 87 ],
   alphaCSR[ 180 ][ 88 ],
   alphaCSR[ 180 ][ 89 ],
   alphaCSR[ 180 ][ 90 ],
   alphaCSR[ 180 ][ 91 ],
   alphaCSR[ 180 ][ 92 ],
   alphaCSR[ 180 ][ 93 ],
   alphaCSR[ 180 ][ 94 ],
   alphaCSR[ 180 ][ 95 ],
   alphaCSR[ 180 ][ 96 ],
   alphaCSR[ 180 ][ 97 ],
   alphaCSR[ 180 ][ 98 ],
   alphaCSR[ 180 ][ 99 ],
   alphaCSR[ 180 ][ 100 ],
   alphaCSR[ 180 ][ 101 ],
   alphaCSR[ 180 ][ 102 ],
   alphaCSR[ 180 ][ 103 ],
   alphaCSR[ 180 ][ 104 ],
   alphaCSR[ 180 ][ 105 ],
   alphaCSR[ 180 ][ 106 ],
   alphaCSR[ 180 ][ 107 ],
   alphaCSR[ 180 ][ 108 ],
   alphaCSR[ 180 ][ 109 ],
   alphaCSR[ 180 ][ 110 ],
   alphaCSR[ 180 ][ 111 ],
   alphaCSR[ 180 ][ 112 ],
   alphaCSR[ 180 ][ 113 ],
   alphaCSR[ 180 ][ 114 ],
   alphaCSR[ 180 ][ 115 ],
   alphaCSR[ 180 ][ 116 ],
   alphaCSR[ 180 ][ 117 ],
   alphaCSR[ 180 ][ 118 ],
   alphaCSR[ 180 ][ 119 ],
   alphaCSR[ 180 ][ 120 ],
   alphaCSR[ 180 ][ 121 ],
   alphaCSR[ 180 ][ 122 ],
   alphaCSR[ 180 ][ 123 ],
   alphaCSR[ 180 ][ 124 ],
   alphaCSR[ 180 ][ 125 ],
   alphaCSR[ 180 ][ 126 ],
   alphaCSR[ 180 ][ 127 ],
   alphaCSR[ 180 ][ 128 ],
   alphaCSR[ 180 ][ 129 ],
   alphaCSR[ 180 ][ 130 ],
   alphaCSR[ 180 ][ 131 ],
   alphaCSR[ 180 ][ 132 ],
   alphaCSR[ 180 ][ 133 ],
   alphaCSR[ 180 ][ 134 ],
   alphaCSR[ 180 ][ 135 ],
   alphaCSR[ 180 ][ 136 ],
   alphaCSR[ 180 ][ 137 ],
   alphaCSR[ 180 ][ 138 ],
   alphaCSR[ 180 ][ 139 ],
   alphaCSR[ 180 ][ 140 ],
   alphaCSR[ 180 ][ 141 ],
   alphaCSR[ 180 ][ 142 ],
   alphaCSR[ 180 ][ 143 ],
   alphaCSR[ 180 ][ 144 ],
   alphaCSR[ 180 ][ 145 ],
   alphaCSR[ 180 ][ 146 ],
   alphaCSR[ 180 ][ 147 ],
   alphaCSR[ 180 ][ 148 ],
   alphaCSR[ 180 ][ 149 ],
   alphaCSR[ 180 ][ 150 ],
   alphaCSR[ 180 ][ 151 ],
   alphaCSR[ 180 ][ 152 ],
   alphaCSR[ 180 ][ 153 ],
   alphaCSR[ 180 ][ 154 ],
   alphaCSR[ 180 ][ 155 ],
   alphaCSR[ 180 ][ 156 ],
   alphaCSR[ 180 ][ 157 ],
   alphaCSR[ 180 ][ 158 ],
   alphaCSR[ 180 ][ 159 ],
   alphaCSR[ 180 ][ 160 ],
   alphaCSR[ 180 ][ 161 ],
   alphaCSR[ 180 ][ 162 ],
   alphaCSR[ 180 ][ 163 ],
   alphaCSR[ 180 ][ 164 ],
   alphaCSR[ 180 ][ 165 ],
   alphaCSR[ 180 ][ 166 ],
   alphaCSR[ 180 ][ 167 ],
   alphaCSR[ 180 ][ 168 ],
   alphaCSR[ 180 ][ 169 ],
   alphaCSR[ 180 ][ 170 ],
   alphaCSR[ 180 ][ 171 ],
   alphaCSR[ 180 ][ 172 ],
   alphaCSR[ 180 ][ 173 ],
   alphaCSR[ 180 ][ 174 ],
   alphaCSR[ 180 ][ 175 ],
   alphaCSR[ 180 ][ 176 ],
   alphaCSR[ 180 ][ 177 ],
   alphaCSR[ 180 ][ 178 ],
   alphaCSR[ 180 ][ 179 ],
   alphaCSR[ 180 ][ 180 ],
   alphaCSR[ 180 ][ 181 ],
   alphaCSR[ 180 ][ 182 ],
   alphaCSR[ 180 ][ 183 ],
   alphaCSR[ 180 ][ 184 ],
   alphaCSR[ 180 ][ 185 ],
   alphaCSR[ 180 ][ 186 ],
   alphaCSR[ 180 ][ 187 ],
   alphaCSR[ 180 ][ 188 ],
   alphaCSR[ 180 ][ 189 ],
   alphaCSR[ 180 ][ 190 ],
   alphaCSR[ 180 ][ 191 ],
   alphaCSR[ 180 ][ 192 ],
   alphaCSR[ 180 ][ 193 ],
   alphaCSR[ 180 ][ 194 ],
   alphaCSR[ 180 ][ 195 ],
   alphaCSR[ 180 ][ 196 ],
   alphaCSR[ 180 ][ 197 ],
   alphaCSR[ 180 ][ 198 ],
   alphaCSR[ 180 ][ 199 ],
   alphaCSR[ 180 ][ 200 ],
   alphaCSR[ 180 ][ 201 ],
   alphaCSR[ 180 ][ 202 ],
   alphaCSR[ 180 ][ 203 ],
   alphaCSR[ 180 ][ 204 ],
   alphaCSR[ 180 ][ 205 ],
   alphaCSR[ 180 ][ 206 ],
   alphaCSR[ 180 ][ 207 ],
   alphaCSR[ 180 ][ 208 ],
   alphaCSR[ 180 ][ 209 ],
   alphaCSR[ 180 ][ 210 ],
   alphaCSR[ 180 ][ 211 ],
   alphaCSR[ 180 ][ 212 ],
   alphaCSR[ 180 ][ 213 ],
   alphaCSR[ 180 ][ 214 ],
   alphaCSR[ 180 ][ 215 ],
   alphaCSR[ 180 ][ 216 ],
   alphaCSR[ 180 ][ 217 ],
   alphaCSR[ 180 ][ 218 ],
   alphaCSR[ 180 ][ 219 ],
   alphaCSR[ 180 ][ 220 ],
   alphaCSR[ 180 ][ 221 ],
   alphaCSR[ 180 ][ 222 ],
   alphaCSR[ 180 ][ 223 ],
   alphaCSR[ 180 ][ 224 ],
   alphaCSR[ 180 ][ 225 ],
   alphaCSR[ 180 ][ 226 ],
   alphaCSR[ 180 ][ 227 ],
   alphaCSR[ 180 ][ 228 ],
   alphaCSR[ 180 ][ 229 ],
   alphaCSR[ 180 ][ 230 ],
   alphaCSR[ 180 ][ 231 ],
   alphaCSR[ 180 ][ 232 ],
   alphaCSR[ 180 ][ 233 ],
   alphaCSR[ 180 ][ 234 ],
   alphaCSR[ 180 ][ 235 ],
   alphaCSR[ 180 ][ 236 ],
   alphaCSR[ 180 ][ 237 ],
   alphaCSR[ 180 ][ 238 ],
   alphaCSR[ 180 ][ 239 ],
   alphaCSR[ 180 ][ 240 ],
   alphaCSR[ 180 ][ 241 ],
   alphaCSR[ 180 ][ 242 ],
   alphaCSR[ 180 ][ 243 ],
   alphaCSR[ 180 ][ 244 ],
   alphaCSR[ 180 ][ 245 ],
   alphaCSR[ 180 ][ 246 ],
   alphaCSR[ 180 ][ 247 ],
   alphaCSR[ 180 ][ 248 ],
   alphaCSR[ 180 ][ 249 ],
   alphaCSR[ 180 ][ 250 ],
   alphaCSR[ 180 ][ 251 ],
   alphaCSR[ 180 ][ 252 ],
   alphaCSR[ 180 ][ 253 ],
   alphaCSR[ 180 ][ 254 ],
   alphaCSR[ 180 ][ 255 ],
   alphaCSR[ 180 ][ 256 ],
   alphaCSR[ 180 ][ 257 ],
   alphaCSR[ 180 ][ 258 ],
   alphaCSR[ 180 ][ 259 ],
   alphaCSR[ 180 ][ 260 ],
   alphaCSR[ 180 ][ 261 ],
   alphaCSR[ 180 ][ 262 ],
   alphaCSR[ 180 ][ 263 ],
   alphaCSR[ 180 ][ 264 ],
   alphaCSR[ 180 ][ 265 ],
   alphaCSR[ 180 ][ 266 ],
   alphaCSR[ 180 ][ 267 ],
   alphaCSR[ 180 ][ 268 ],
   alphaCSR[ 180 ][ 269 ],
   alphaCSR[ 180 ][ 270 ],
   alphaCSR[ 180 ][ 271 ],
   alphaCSR[ 180 ][ 272 ],
   alphaCSR[ 180 ][ 273 ],
   alphaCSR[ 180 ][ 274 ],
   alphaCSR[ 180 ][ 275 ],
   alphaCSR[ 180 ][ 276 ],
   alphaCSR[ 180 ][ 277 ],
   alphaCSR[ 180 ][ 278 ],
   alphaCSR[ 180 ][ 279 ],
   alphaCSR[ 180 ][ 280 ],
   alphaCSR[ 180 ][ 281 ],
   alphaCSR[ 180 ][ 282 ],
   alphaCSR[ 180 ][ 283 ],
   alphaCSR[ 180 ][ 284 ],
   alphaCSR[ 180 ][ 285 ],
   alphaCSR[ 180 ][ 286 ],
   alphaCSR[ 180 ][ 287 ],
   alphaCSR[ 180 ][ 288 ],
   alphaCSR[ 180 ][ 289 ],
   alphaCSR[ 180 ][ 290 ],
   alphaCSR[ 180 ][ 291 ],
   alphaCSR[ 180 ][ 292 ],
   alphaCSR[ 180 ][ 293 ],
   alphaCSR[ 180 ][ 294 ],
   alphaCSR[ 180 ][ 295 ],
   alphaCSR[ 180 ][ 296 ],
   alphaCSR[ 180 ][ 297 ],
   alphaCSR[ 180 ][ 298 ],
   alphaCSR[ 180 ][ 299 ],
   alphaCSR[ 180 ][ 300 ],
   alphaCSR[ 180 ][ 301 ],
   alphaCSR[ 180 ][ 302 ],
   alphaCSR[ 180 ][ 303 ],
   alphaCSR[ 180 ][ 304 ],
   alphaCSR[ 180 ][ 305 ],
   alphaCSR[ 180 ][ 306 ],
   alphaCSR[ 180 ][ 307 ],
   alphaCSR[ 180 ][ 308 ],
   alphaCSR[ 180 ][ 309 ],
   alphaCSR[ 180 ][ 310 ],
   alphaCSR[ 180 ][ 311 ],
   alphaCSR[ 180 ][ 312 ],
   alphaCSR[ 180 ][ 313 ],
   alphaCSR[ 180 ][ 314 ],
   alphaCSR[ 180 ][ 315 ],
   alphaCSR[ 180 ][ 316 ],
   alphaCSR[ 180 ][ 317 ],
   alphaCSR[ 180 ][ 318 ],
   alphaCSR[ 180 ][ 319 ],
   alphaCSR[ 180 ][ 320 ],
   alphaCSR[ 180 ][ 321 ],
   alphaCSR[ 180 ][ 322 ],
   alphaCSR[ 180 ][ 323 ],
   alphaCSR[ 180 ][ 324 ],
   alphaCSR[ 180 ][ 325 ],
   alphaCSR[ 180 ][ 326 ],
   alphaCSR[ 180 ][ 327 ],
   alphaCSR[ 180 ][ 328 ],
   alphaCSR[ 180 ][ 329 ],
   alphaCSR[ 180 ][ 330 ],
   alphaCSR[ 180 ][ 331 ],
   alphaCSR[ 180 ][ 332 ],
   alphaCSR[ 180 ][ 333 ],
   alphaCSR[ 180 ][ 334 ],
   alphaCSR[ 180 ][ 335 ],
   alphaCSR[ 180 ][ 336 ],
   alphaCSR[ 180 ][ 337 ],
   alphaCSR[ 180 ][ 338 ],
   alphaCSR[ 180 ][ 339 ],
   alphaCSR[ 180 ][ 340 ],
   alphaCSR[ 180 ][ 341 ],
   alphaCSR[ 180 ][ 342 ],
   alphaCSR[ 180 ][ 343 ],
   alphaCSR[ 180 ][ 344 ],
   alphaCSR[ 180 ][ 345 ],
   alphaCSR[ 180 ][ 346 ],
   alphaCSR[ 180 ][ 347 ],
   alphaCSR[ 180 ][ 348 ],
   alphaCSR[ 180 ][ 349 ],
   alphaCSR[ 180 ][ 350 ],
   alphaCSR[ 180 ][ 351 ],
   alphaCSR[ 180 ][ 352 ],
   alphaCSR[ 180 ][ 353 ],
   alphaCSR[ 180 ][ 354 ],
   alphaCSR[ 180 ][ 355 ],
   alphaCSR[ 180 ][ 356 ],
   alphaCSR[ 180 ][ 357 ],
   alphaCSR[ 180 ][ 358 ],
   alphaCSR[ 180 ][ 359 ],
   alphaCSR[ 180 ][ 360 ],
   alphaCSR[ 180 ][ 361 ],
   alphaCSR[ 180 ][ 362 ],
   alphaCSR[ 180 ][ 363 ],
   alphaCSR[ 180 ][ 364 ],
   alphaCSR[ 180 ][ 365 ],
   alphaCSR[ 180 ][ 366 ],
   alphaCSR[ 180 ][ 367 ],
   alphaCSR[ 180 ][ 368 ],
   alphaCSR[ 180 ][ 369 ],
   alphaCSR[ 180 ][ 370 ],
   alphaCSR[ 180 ][ 371 ],
   alphaCSR[ 180 ][ 372 ],
   alphaCSR[ 180 ][ 373 ],
   alphaCSR[ 180 ][ 374 ],
   alphaCSR[ 180 ][ 375 ],
   alphaCSR[ 180 ][ 376 ],
   alphaCSR[ 180 ][ 377 ],
   alphaCSR[ 180 ][ 378 ],
   alphaCSR[ 180 ][ 379 ],
   alphaCSR[ 180 ][ 380 ],
   alphaCSR[ 180 ][ 381 ],
   alphaCSR[ 180 ][ 382 ],
   alphaCSR[ 180 ][ 383 ],
   alphaCSR[ 181 ][ 0 ],
   alphaCSR[ 181 ][ 1 ],
   alphaCSR[ 181 ][ 2 ],
   alphaCSR[ 181 ][ 3 ],
   alphaCSR[ 181 ][ 4 ],
   alphaCSR[ 181 ][ 5 ],
   alphaCSR[ 181 ][ 6 ],
   alphaCSR[ 181 ][ 7 ],
   alphaCSR[ 181 ][ 8 ],
   alphaCSR[ 181 ][ 9 ],
   alphaCSR[ 181 ][ 10 ],
   alphaCSR[ 181 ][ 11 ],
   alphaCSR[ 181 ][ 12 ],
   alphaCSR[ 181 ][ 13 ],
   alphaCSR[ 181 ][ 14 ],
   alphaCSR[ 181 ][ 15 ],
   alphaCSR[ 181 ][ 16 ],
   alphaCSR[ 181 ][ 17 ],
   alphaCSR[ 181 ][ 18 ],
   alphaCSR[ 181 ][ 19 ],
   alphaCSR[ 181 ][ 20 ],
   alphaCSR[ 181 ][ 21 ],
   alphaCSR[ 181 ][ 22 ],
   alphaCSR[ 181 ][ 23 ],
   alphaCSR[ 181 ][ 24 ],
   alphaCSR[ 181 ][ 25 ],
   alphaCSR[ 181 ][ 26 ],
   alphaCSR[ 181 ][ 27 ],
   alphaCSR[ 181 ][ 28 ],
   alphaCSR[ 181 ][ 29 ],
   alphaCSR[ 181 ][ 30 ],
   alphaCSR[ 181 ][ 31 ],
   alphaCSR[ 181 ][ 32 ],
   alphaCSR[ 181 ][ 33 ],
   alphaCSR[ 181 ][ 34 ],
   alphaCSR[ 181 ][ 35 ],
   alphaCSR[ 181 ][ 36 ],
   alphaCSR[ 181 ][ 37 ],
   alphaCSR[ 181 ][ 38 ],
   alphaCSR[ 181 ][ 39 ],
   alphaCSR[ 181 ][ 40 ],
   alphaCSR[ 181 ][ 41 ],
   alphaCSR[ 181 ][ 42 ],
   alphaCSR[ 181 ][ 43 ],
   alphaCSR[ 181 ][ 44 ],
   alphaCSR[ 181 ][ 45 ],
   alphaCSR[ 181 ][ 46 ],
   alphaCSR[ 181 ][ 47 ],
   alphaCSR[ 181 ][ 48 ],
   alphaCSR[ 181 ][ 49 ],
   alphaCSR[ 181 ][ 50 ],
   alphaCSR[ 181 ][ 51 ],
   alphaCSR[ 181 ][ 52 ],
   alphaCSR[ 181 ][ 53 ],
   alphaCSR[ 181 ][ 54 ],
   alphaCSR[ 181 ][ 55 ],
   alphaCSR[ 181 ][ 56 ],
   alphaCSR[ 181 ][ 57 ],
   alphaCSR[ 181 ][ 58 ],
   alphaCSR[ 181 ][ 59 ],
   alphaCSR[ 181 ][ 60 ],
   alphaCSR[ 181 ][ 61 ],
   alphaCSR[ 181 ][ 62 ],
   alphaCSR[ 181 ][ 63 ],
   alphaCSR[ 181 ][ 64 ],
   alphaCSR[ 181 ][ 65 ],
   alphaCSR[ 181 ][ 66 ],
   alphaCSR[ 181 ][ 67 ],
   alphaCSR[ 181 ][ 68 ],
   alphaCSR[ 181 ][ 69 ],
   alphaCSR[ 181 ][ 70 ],
   alphaCSR[ 181 ][ 71 ],
   alphaCSR[ 181 ][ 72 ],
   alphaCSR[ 181 ][ 73 ],
   alphaCSR[ 181 ][ 74 ],
   alphaCSR[ 181 ][ 75 ],
   alphaCSR[ 181 ][ 76 ],
   alphaCSR[ 181 ][ 77 ],
   alphaCSR[ 181 ][ 78 ],
   alphaCSR[ 181 ][ 79 ],
   alphaCSR[ 181 ][ 80 ],
   alphaCSR[ 181 ][ 81 ],
   alphaCSR[ 181 ][ 82 ],
   alphaCSR[ 181 ][ 83 ],
   alphaCSR[ 181 ][ 84 ],
   alphaCSR[ 181 ][ 85 ],
   alphaCSR[ 181 ][ 86 ],
   alphaCSR[ 181 ][ 87 ],
   alphaCSR[ 181 ][ 88 ],
   alphaCSR[ 181 ][ 89 ],
   alphaCSR[ 181 ][ 90 ],
   alphaCSR[ 181 ][ 91 ],
   alphaCSR[ 181 ][ 92 ],
   alphaCSR[ 181 ][ 93 ],
   alphaCSR[ 181 ][ 94 ],
   alphaCSR[ 181 ][ 95 ],
   alphaCSR[ 181 ][ 96 ],
   alphaCSR[ 181 ][ 97 ],
   alphaCSR[ 181 ][ 98 ],
   alphaCSR[ 181 ][ 99 ],
   alphaCSR[ 181 ][ 100 ],
   alphaCSR[ 181 ][ 101 ],
   alphaCSR[ 181 ][ 102 ],
   alphaCSR[ 181 ][ 103 ],
   alphaCSR[ 181 ][ 104 ],
   alphaCSR[ 181 ][ 105 ],
   alphaCSR[ 181 ][ 106 ],
   alphaCSR[ 181 ][ 107 ],
   alphaCSR[ 181 ][ 108 ],
   alphaCSR[ 181 ][ 109 ],
   alphaCSR[ 181 ][ 110 ],
   alphaCSR[ 181 ][ 111 ],
   alphaCSR[ 181 ][ 112 ],
   alphaCSR[ 181 ][ 113 ],
   alphaCSR[ 181 ][ 114 ],
   alphaCSR[ 181 ][ 115 ],
   alphaCSR[ 181 ][ 116 ],
   alphaCSR[ 181 ][ 117 ],
   alphaCSR[ 181 ][ 118 ],
   alphaCSR[ 181 ][ 119 ],
   alphaCSR[ 181 ][ 120 ],
   alphaCSR[ 181 ][ 121 ],
   alphaCSR[ 181 ][ 122 ],
   alphaCSR[ 181 ][ 123 ],
   alphaCSR[ 181 ][ 124 ],
   alphaCSR[ 181 ][ 125 ],
   alphaCSR[ 181 ][ 126 ],
   alphaCSR[ 181 ][ 127 ],
   alphaCSR[ 181 ][ 128 ],
   alphaCSR[ 181 ][ 129 ],
   alphaCSR[ 181 ][ 130 ],
   alphaCSR[ 181 ][ 131 ],
   alphaCSR[ 181 ][ 132 ],
   alphaCSR[ 181 ][ 133 ],
   alphaCSR[ 181 ][ 134 ],
   alphaCSR[ 181 ][ 135 ],
   alphaCSR[ 181 ][ 136 ],
   alphaCSR[ 181 ][ 137 ],
   alphaCSR[ 181 ][ 138 ],
   alphaCSR[ 181 ][ 139 ],
   alphaCSR[ 181 ][ 140 ],
   alphaCSR[ 181 ][ 141 ],
   alphaCSR[ 181 ][ 142 ],
   alphaCSR[ 181 ][ 143 ],
   alphaCSR[ 181 ][ 144 ],
   alphaCSR[ 181 ][ 145 ],
   alphaCSR[ 181 ][ 146 ],
   alphaCSR[ 181 ][ 147 ],
   alphaCSR[ 181 ][ 148 ],
   alphaCSR[ 181 ][ 149 ],
   alphaCSR[ 181 ][ 150 ],
   alphaCSR[ 181 ][ 151 ],
   alphaCSR[ 181 ][ 152 ],
   alphaCSR[ 181 ][ 153 ],
   alphaCSR[ 181 ][ 154 ],
   alphaCSR[ 181 ][ 155 ],
   alphaCSR[ 181 ][ 156 ],
   alphaCSR[ 181 ][ 157 ],
   alphaCSR[ 181 ][ 158 ],
   alphaCSR[ 181 ][ 159 ],
   alphaCSR[ 181 ][ 160 ],
   alphaCSR[ 181 ][ 161 ],
   alphaCSR[ 181 ][ 162 ],
   alphaCSR[ 181 ][ 163 ],
   alphaCSR[ 181 ][ 164 ],
   alphaCSR[ 181 ][ 165 ],
   alphaCSR[ 181 ][ 166 ],
   alphaCSR[ 181 ][ 167 ],
   alphaCSR[ 181 ][ 168 ],
   alphaCSR[ 181 ][ 169 ],
   alphaCSR[ 181 ][ 170 ],
   alphaCSR[ 181 ][ 171 ],
   alphaCSR[ 181 ][ 172 ],
   alphaCSR[ 181 ][ 173 ],
   alphaCSR[ 181 ][ 174 ],
   alphaCSR[ 181 ][ 175 ],
   alphaCSR[ 181 ][ 176 ],
   alphaCSR[ 181 ][ 177 ],
   alphaCSR[ 181 ][ 178 ],
   alphaCSR[ 181 ][ 179 ],
   alphaCSR[ 181 ][ 180 ],
   alphaCSR[ 181 ][ 181 ],
   alphaCSR[ 181 ][ 182 ],
   alphaCSR[ 181 ][ 183 ],
   alphaCSR[ 181 ][ 184 ],
   alphaCSR[ 181 ][ 185 ],
   alphaCSR[ 181 ][ 186 ],
   alphaCSR[ 181 ][ 187 ],
   alphaCSR[ 181 ][ 188 ],
   alphaCSR[ 181 ][ 189 ],
   alphaCSR[ 181 ][ 190 ],
   alphaCSR[ 181 ][ 191 ],
   alphaCSR[ 181 ][ 192 ],
   alphaCSR[ 181 ][ 193 ],
   alphaCSR[ 181 ][ 194 ],
   alphaCSR[ 181 ][ 195 ],
   alphaCSR[ 181 ][ 196 ],
   alphaCSR[ 181 ][ 197 ],
   alphaCSR[ 181 ][ 198 ],
   alphaCSR[ 181 ][ 199 ],
   alphaCSR[ 181 ][ 200 ],
   alphaCSR[ 181 ][ 201 ],
   alphaCSR[ 181 ][ 202 ],
   alphaCSR[ 181 ][ 203 ],
   alphaCSR[ 181 ][ 204 ],
   alphaCSR[ 181 ][ 205 ],
   alphaCSR[ 181 ][ 206 ],
   alphaCSR[ 181 ][ 207 ],
   alphaCSR[ 181 ][ 208 ],
   alphaCSR[ 181 ][ 209 ],
   alphaCSR[ 181 ][ 210 ],
   alphaCSR[ 181 ][ 211 ],
   alphaCSR[ 181 ][ 212 ],
   alphaCSR[ 181 ][ 213 ],
   alphaCSR[ 181 ][ 214 ],
   alphaCSR[ 181 ][ 215 ],
   alphaCSR[ 181 ][ 216 ],
   alphaCSR[ 181 ][ 217 ],
   alphaCSR[ 181 ][ 218 ],
   alphaCSR[ 181 ][ 219 ],
   alphaCSR[ 181 ][ 220 ],
   alphaCSR[ 181 ][ 221 ],
   alphaCSR[ 181 ][ 222 ],
   alphaCSR[ 181 ][ 223 ],
   alphaCSR[ 181 ][ 224 ],
   alphaCSR[ 181 ][ 225 ],
   alphaCSR[ 181 ][ 226 ],
   alphaCSR[ 181 ][ 227 ],
   alphaCSR[ 181 ][ 228 ],
   alphaCSR[ 181 ][ 229 ],
   alphaCSR[ 181 ][ 230 ],
   alphaCSR[ 181 ][ 231 ],
   alphaCSR[ 181 ][ 232 ],
   alphaCSR[ 181 ][ 233 ],
   alphaCSR[ 181 ][ 234 ],
   alphaCSR[ 181 ][ 235 ],
   alphaCSR[ 181 ][ 236 ],
   alphaCSR[ 181 ][ 237 ],
   alphaCSR[ 181 ][ 238 ],
   alphaCSR[ 181 ][ 239 ],
   alphaCSR[ 181 ][ 240 ],
   alphaCSR[ 181 ][ 241 ],
   alphaCSR[ 181 ][ 242 ],
   alphaCSR[ 181 ][ 243 ],
   alphaCSR[ 181 ][ 244 ],
   alphaCSR[ 181 ][ 245 ],
   alphaCSR[ 181 ][ 246 ],
   alphaCSR[ 181 ][ 247 ],
   alphaCSR[ 181 ][ 248 ],
   alphaCSR[ 181 ][ 249 ],
   alphaCSR[ 181 ][ 250 ],
   alphaCSR[ 181 ][ 251 ],
   alphaCSR[ 181 ][ 252 ],
   alphaCSR[ 181 ][ 253 ],
   alphaCSR[ 181 ][ 254 ],
   alphaCSR[ 181 ][ 255 ],
   alphaCSR[ 181 ][ 256 ],
   alphaCSR[ 181 ][ 257 ],
   alphaCSR[ 181 ][ 258 ],
   alphaCSR[ 181 ][ 259 ],
   alphaCSR[ 181 ][ 260 ],
   alphaCSR[ 181 ][ 261 ],
   alphaCSR[ 181 ][ 262 ],
   alphaCSR[ 181 ][ 263 ],
   alphaCSR[ 181 ][ 264 ],
   alphaCSR[ 181 ][ 265 ],
   alphaCSR[ 181 ][ 266 ],
   alphaCSR[ 181 ][ 267 ],
   alphaCSR[ 181 ][ 268 ],
   alphaCSR[ 181 ][ 269 ],
   alphaCSR[ 181 ][ 270 ],
   alphaCSR[ 181 ][ 271 ],
   alphaCSR[ 181 ][ 272 ],
   alphaCSR[ 181 ][ 273 ],
   alphaCSR[ 181 ][ 274 ],
   alphaCSR[ 181 ][ 275 ],
   alphaCSR[ 181 ][ 276 ],
   alphaCSR[ 181 ][ 277 ],
   alphaCSR[ 181 ][ 278 ],
   alphaCSR[ 181 ][ 279 ],
   alphaCSR[ 181 ][ 280 ],
   alphaCSR[ 181 ][ 281 ],
   alphaCSR[ 181 ][ 282 ],
   alphaCSR[ 181 ][ 283 ],
   alphaCSR[ 181 ][ 284 ],
   alphaCSR[ 181 ][ 285 ],
   alphaCSR[ 181 ][ 286 ],
   alphaCSR[ 181 ][ 287 ],
   alphaCSR[ 181 ][ 288 ],
   alphaCSR[ 181 ][ 289 ],
   alphaCSR[ 181 ][ 290 ],
   alphaCSR[ 181 ][ 291 ],
   alphaCSR[ 181 ][ 292 ],
   alphaCSR[ 181 ][ 293 ],
   alphaCSR[ 181 ][ 294 ],
   alphaCSR[ 181 ][ 295 ],
   alphaCSR[ 181 ][ 296 ],
   alphaCSR[ 181 ][ 297 ],
   alphaCSR[ 181 ][ 298 ],
   alphaCSR[ 181 ][ 299 ],
   alphaCSR[ 181 ][ 300 ],
   alphaCSR[ 181 ][ 301 ],
   alphaCSR[ 181 ][ 302 ],
   alphaCSR[ 181 ][ 303 ],
   alphaCSR[ 181 ][ 304 ],
   alphaCSR[ 181 ][ 305 ],
   alphaCSR[ 181 ][ 306 ],
   alphaCSR[ 181 ][ 307 ],
   alphaCSR[ 181 ][ 308 ],
   alphaCSR[ 181 ][ 309 ],
   alphaCSR[ 181 ][ 310 ],
   alphaCSR[ 181 ][ 311 ],
   alphaCSR[ 181 ][ 312 ],
   alphaCSR[ 181 ][ 313 ],
   alphaCSR[ 181 ][ 314 ],
   alphaCSR[ 181 ][ 315 ],
   alphaCSR[ 181 ][ 316 ],
   alphaCSR[ 181 ][ 317 ],
   alphaCSR[ 181 ][ 318 ],
   alphaCSR[ 181 ][ 319 ],
   alphaCSR[ 181 ][ 320 ],
   alphaCSR[ 181 ][ 321 ],
   alphaCSR[ 181 ][ 322 ],
   alphaCSR[ 181 ][ 323 ],
   alphaCSR[ 181 ][ 324 ],
   alphaCSR[ 181 ][ 325 ],
   alphaCSR[ 181 ][ 326 ],
   alphaCSR[ 181 ][ 327 ],
   alphaCSR[ 181 ][ 328 ],
   alphaCSR[ 181 ][ 329 ],
   alphaCSR[ 181 ][ 330 ],
   alphaCSR[ 181 ][ 331 ],
   alphaCSR[ 181 ][ 332 ],
   alphaCSR[ 181 ][ 333 ],
   alphaCSR[ 181 ][ 334 ],
   alphaCSR[ 181 ][ 335 ],
   alphaCSR[ 181 ][ 336 ],
   alphaCSR[ 181 ][ 337 ],
   alphaCSR[ 181 ][ 338 ],
   alphaCSR[ 181 ][ 339 ],
   alphaCSR[ 181 ][ 340 ],
   alphaCSR[ 181 ][ 341 ],
   alphaCSR[ 181 ][ 342 ],
   alphaCSR[ 181 ][ 343 ],
   alphaCSR[ 181 ][ 344 ],
   alphaCSR[ 181 ][ 345 ],
   alphaCSR[ 181 ][ 346 ],
   alphaCSR[ 181 ][ 347 ],
   alphaCSR[ 181 ][ 348 ],
   alphaCSR[ 181 ][ 349 ],
   alphaCSR[ 181 ][ 350 ],
   alphaCSR[ 181 ][ 351 ],
   alphaCSR[ 181 ][ 352 ],
   alphaCSR[ 181 ][ 353 ],
   alphaCSR[ 181 ][ 354 ],
   alphaCSR[ 181 ][ 355 ],
   alphaCSR[ 181 ][ 356 ],
   alphaCSR[ 181 ][ 357 ],
   alphaCSR[ 181 ][ 358 ],
   alphaCSR[ 181 ][ 359 ],
   alphaCSR[ 181 ][ 360 ],
   alphaCSR[ 181 ][ 361 ],
   alphaCSR[ 181 ][ 362 ],
   alphaCSR[ 181 ][ 363 ],
   alphaCSR[ 181 ][ 364 ],
   alphaCSR[ 181 ][ 365 ],
   alphaCSR[ 181 ][ 366 ],
   alphaCSR[ 181 ][ 367 ],
   alphaCSR[ 181 ][ 368 ],
   alphaCSR[ 181 ][ 369 ],
   alphaCSR[ 181 ][ 370 ],
   alphaCSR[ 181 ][ 371 ],
   alphaCSR[ 181 ][ 372 ],
   alphaCSR[ 181 ][ 373 ],
   alphaCSR[ 181 ][ 374 ],
   alphaCSR[ 181 ][ 375 ],
   alphaCSR[ 181 ][ 376 ],
   alphaCSR[ 181 ][ 377 ],
   alphaCSR[ 181 ][ 378 ],
   alphaCSR[ 181 ][ 379 ],
   alphaCSR[ 181 ][ 380 ],
   alphaCSR[ 181 ][ 381 ],
   alphaCSR[ 181 ][ 382 ],
   alphaCSR[ 181 ][ 383 ],
   alphaCSR[ 182 ][ 0 ],
   alphaCSR[ 182 ][ 1 ],
   alphaCSR[ 182 ][ 2 ],
   alphaCSR[ 182 ][ 3 ],
   alphaCSR[ 182 ][ 4 ],
   alphaCSR[ 182 ][ 5 ],
   alphaCSR[ 182 ][ 6 ],
   alphaCSR[ 182 ][ 7 ],
   alphaCSR[ 182 ][ 8 ],
   alphaCSR[ 182 ][ 9 ],
   alphaCSR[ 182 ][ 10 ],
   alphaCSR[ 182 ][ 11 ],
   alphaCSR[ 182 ][ 12 ],
   alphaCSR[ 182 ][ 13 ],
   alphaCSR[ 182 ][ 14 ],
   alphaCSR[ 182 ][ 15 ],
   alphaCSR[ 182 ][ 16 ],
   alphaCSR[ 182 ][ 17 ],
   alphaCSR[ 182 ][ 18 ],
   alphaCSR[ 182 ][ 19 ],
   alphaCSR[ 182 ][ 20 ],
   alphaCSR[ 182 ][ 21 ],
   alphaCSR[ 182 ][ 22 ],
   alphaCSR[ 182 ][ 23 ],
   alphaCSR[ 182 ][ 24 ],
   alphaCSR[ 182 ][ 25 ],
   alphaCSR[ 182 ][ 26 ],
   alphaCSR[ 182 ][ 27 ],
   alphaCSR[ 182 ][ 28 ],
   alphaCSR[ 182 ][ 29 ],
   alphaCSR[ 182 ][ 30 ],
   alphaCSR[ 182 ][ 31 ],
   alphaCSR[ 182 ][ 32 ],
   alphaCSR[ 182 ][ 33 ],
   alphaCSR[ 182 ][ 34 ],
   alphaCSR[ 182 ][ 35 ],
   alphaCSR[ 182 ][ 36 ],
   alphaCSR[ 182 ][ 37 ],
   alphaCSR[ 182 ][ 38 ],
   alphaCSR[ 182 ][ 39 ],
   alphaCSR[ 182 ][ 40 ],
   alphaCSR[ 182 ][ 41 ],
   alphaCSR[ 182 ][ 42 ],
   alphaCSR[ 182 ][ 43 ],
   alphaCSR[ 182 ][ 44 ],
   alphaCSR[ 182 ][ 45 ],
   alphaCSR[ 182 ][ 46 ],
   alphaCSR[ 182 ][ 47 ],
   alphaCSR[ 182 ][ 48 ],
   alphaCSR[ 182 ][ 49 ],
   alphaCSR[ 182 ][ 50 ],
   alphaCSR[ 182 ][ 51 ],
   alphaCSR[ 182 ][ 52 ],
   alphaCSR[ 182 ][ 53 ],
   alphaCSR[ 182 ][ 54 ],
   alphaCSR[ 182 ][ 55 ],
   alphaCSR[ 182 ][ 56 ],
   alphaCSR[ 182 ][ 57 ],
   alphaCSR[ 182 ][ 58 ],
   alphaCSR[ 182 ][ 59 ],
   alphaCSR[ 182 ][ 60 ],
   alphaCSR[ 182 ][ 61 ],
   alphaCSR[ 182 ][ 62 ],
   alphaCSR[ 182 ][ 63 ],
   alphaCSR[ 182 ][ 64 ],
   alphaCSR[ 182 ][ 65 ],
   alphaCSR[ 182 ][ 66 ],
   alphaCSR[ 182 ][ 67 ],
   alphaCSR[ 182 ][ 68 ],
   alphaCSR[ 182 ][ 69 ],
   alphaCSR[ 182 ][ 70 ],
   alphaCSR[ 182 ][ 71 ],
   alphaCSR[ 182 ][ 72 ],
   alphaCSR[ 182 ][ 73 ],
   alphaCSR[ 182 ][ 74 ],
   alphaCSR[ 182 ][ 75 ],
   alphaCSR[ 182 ][ 76 ],
   alphaCSR[ 182 ][ 77 ],
   alphaCSR[ 182 ][ 78 ],
   alphaCSR[ 182 ][ 79 ],
   alphaCSR[ 182 ][ 80 ],
   alphaCSR[ 182 ][ 81 ],
   alphaCSR[ 182 ][ 82 ],
   alphaCSR[ 182 ][ 83 ],
   alphaCSR[ 182 ][ 84 ],
   alphaCSR[ 182 ][ 85 ],
   alphaCSR[ 182 ][ 86 ],
   alphaCSR[ 182 ][ 87 ],
   alphaCSR[ 182 ][ 88 ],
   alphaCSR[ 182 ][ 89 ],
   alphaCSR[ 182 ][ 90 ],
   alphaCSR[ 182 ][ 91 ],
   alphaCSR[ 182 ][ 92 ],
   alphaCSR[ 182 ][ 93 ],
   alphaCSR[ 182 ][ 94 ],
   alphaCSR[ 182 ][ 95 ],
   alphaCSR[ 182 ][ 96 ],
   alphaCSR[ 182 ][ 97 ],
   alphaCSR[ 182 ][ 98 ],
   alphaCSR[ 182 ][ 99 ],
   alphaCSR[ 182 ][ 100 ],
   alphaCSR[ 182 ][ 101 ],
   alphaCSR[ 182 ][ 102 ],
   alphaCSR[ 182 ][ 103 ],
   alphaCSR[ 182 ][ 104 ],
   alphaCSR[ 182 ][ 105 ],
   alphaCSR[ 182 ][ 106 ],
   alphaCSR[ 182 ][ 107 ],
   alphaCSR[ 182 ][ 108 ],
   alphaCSR[ 182 ][ 109 ],
   alphaCSR[ 182 ][ 110 ],
   alphaCSR[ 182 ][ 111 ],
   alphaCSR[ 182 ][ 112 ],
   alphaCSR[ 182 ][ 113 ],
   alphaCSR[ 182 ][ 114 ],
   alphaCSR[ 182 ][ 115 ],
   alphaCSR[ 182 ][ 116 ],
   alphaCSR[ 182 ][ 117 ],
   alphaCSR[ 182 ][ 118 ],
   alphaCSR[ 182 ][ 119 ],
   alphaCSR[ 182 ][ 120 ],
   alphaCSR[ 182 ][ 121 ],
   alphaCSR[ 182 ][ 122 ],
   alphaCSR[ 182 ][ 123 ],
   alphaCSR[ 182 ][ 124 ],
   alphaCSR[ 182 ][ 125 ],
   alphaCSR[ 182 ][ 126 ],
   alphaCSR[ 182 ][ 127 ],
   alphaCSR[ 182 ][ 128 ],
   alphaCSR[ 182 ][ 129 ],
   alphaCSR[ 182 ][ 130 ],
   alphaCSR[ 182 ][ 131 ],
   alphaCSR[ 182 ][ 132 ],
   alphaCSR[ 182 ][ 133 ],
   alphaCSR[ 182 ][ 134 ],
   alphaCSR[ 182 ][ 135 ],
   alphaCSR[ 182 ][ 136 ],
   alphaCSR[ 182 ][ 137 ],
   alphaCSR[ 182 ][ 138 ],
   alphaCSR[ 182 ][ 139 ],
   alphaCSR[ 182 ][ 140 ],
   alphaCSR[ 182 ][ 141 ],
   alphaCSR[ 182 ][ 142 ],
   alphaCSR[ 182 ][ 143 ],
   alphaCSR[ 182 ][ 144 ],
   alphaCSR[ 182 ][ 145 ],
   alphaCSR[ 182 ][ 146 ],
   alphaCSR[ 182 ][ 147 ],
   alphaCSR[ 182 ][ 148 ],
   alphaCSR[ 182 ][ 149 ],
   alphaCSR[ 182 ][ 150 ],
   alphaCSR[ 182 ][ 151 ],
   alphaCSR[ 182 ][ 152 ],
   alphaCSR[ 182 ][ 153 ],
   alphaCSR[ 182 ][ 154 ],
   alphaCSR[ 182 ][ 155 ],
   alphaCSR[ 182 ][ 156 ],
   alphaCSR[ 182 ][ 157 ],
   alphaCSR[ 182 ][ 158 ],
   alphaCSR[ 182 ][ 159 ],
   alphaCSR[ 182 ][ 160 ],
   alphaCSR[ 182 ][ 161 ],
   alphaCSR[ 182 ][ 162 ],
   alphaCSR[ 182 ][ 163 ],
   alphaCSR[ 182 ][ 164 ],
   alphaCSR[ 182 ][ 165 ],
   alphaCSR[ 182 ][ 166 ],
   alphaCSR[ 182 ][ 167 ],
   alphaCSR[ 182 ][ 168 ],
   alphaCSR[ 182 ][ 169 ],
   alphaCSR[ 182 ][ 170 ],
   alphaCSR[ 182 ][ 171 ],
   alphaCSR[ 182 ][ 172 ],
   alphaCSR[ 182 ][ 173 ],
   alphaCSR[ 182 ][ 174 ],
   alphaCSR[ 182 ][ 175 ],
   alphaCSR[ 182 ][ 176 ],
   alphaCSR[ 182 ][ 177 ],
   alphaCSR[ 182 ][ 178 ],
   alphaCSR[ 182 ][ 179 ],
   alphaCSR[ 182 ][ 180 ],
   alphaCSR[ 182 ][ 181 ],
   alphaCSR[ 182 ][ 182 ],
   alphaCSR[ 182 ][ 183 ],
   alphaCSR[ 182 ][ 184 ],
   alphaCSR[ 182 ][ 185 ],
   alphaCSR[ 182 ][ 186 ],
   alphaCSR[ 182 ][ 187 ],
   alphaCSR[ 182 ][ 188 ],
   alphaCSR[ 182 ][ 189 ],
   alphaCSR[ 182 ][ 190 ],
   alphaCSR[ 182 ][ 191 ],
   alphaCSR[ 182 ][ 192 ],
   alphaCSR[ 182 ][ 193 ],
   alphaCSR[ 182 ][ 194 ],
   alphaCSR[ 182 ][ 195 ],
   alphaCSR[ 182 ][ 196 ],
   alphaCSR[ 182 ][ 197 ],
   alphaCSR[ 182 ][ 198 ],
   alphaCSR[ 182 ][ 199 ],
   alphaCSR[ 182 ][ 200 ],
   alphaCSR[ 182 ][ 201 ],
   alphaCSR[ 182 ][ 202 ],
   alphaCSR[ 182 ][ 203 ],
   alphaCSR[ 182 ][ 204 ],
   alphaCSR[ 182 ][ 205 ],
   alphaCSR[ 182 ][ 206 ],
   alphaCSR[ 182 ][ 207 ],
   alphaCSR[ 182 ][ 208 ],
   alphaCSR[ 182 ][ 209 ],
   alphaCSR[ 182 ][ 210 ],
   alphaCSR[ 182 ][ 211 ],
   alphaCSR[ 182 ][ 212 ],
   alphaCSR[ 182 ][ 213 ],
   alphaCSR[ 182 ][ 214 ],
   alphaCSR[ 182 ][ 215 ],
   alphaCSR[ 182 ][ 216 ],
   alphaCSR[ 182 ][ 217 ],
   alphaCSR[ 182 ][ 218 ],
   alphaCSR[ 182 ][ 219 ],
   alphaCSR[ 182 ][ 220 ],
   alphaCSR[ 182 ][ 221 ],
   alphaCSR[ 182 ][ 222 ],
   alphaCSR[ 182 ][ 223 ],
   alphaCSR[ 182 ][ 224 ],
   alphaCSR[ 182 ][ 225 ],
   alphaCSR[ 182 ][ 226 ],
   alphaCSR[ 182 ][ 227 ],
   alphaCSR[ 182 ][ 228 ],
   alphaCSR[ 182 ][ 229 ],
   alphaCSR[ 182 ][ 230 ],
   alphaCSR[ 182 ][ 231 ],
   alphaCSR[ 182 ][ 232 ],
   alphaCSR[ 182 ][ 233 ],
   alphaCSR[ 182 ][ 234 ],
   alphaCSR[ 182 ][ 235 ],
   alphaCSR[ 182 ][ 236 ],
   alphaCSR[ 182 ][ 237 ],
   alphaCSR[ 182 ][ 238 ],
   alphaCSR[ 182 ][ 239 ],
   alphaCSR[ 182 ][ 240 ],
   alphaCSR[ 182 ][ 241 ],
   alphaCSR[ 182 ][ 242 ],
   alphaCSR[ 182 ][ 243 ],
   alphaCSR[ 182 ][ 244 ],
   alphaCSR[ 182 ][ 245 ],
   alphaCSR[ 182 ][ 246 ],
   alphaCSR[ 182 ][ 247 ],
   alphaCSR[ 182 ][ 248 ],
   alphaCSR[ 182 ][ 249 ],
   alphaCSR[ 182 ][ 250 ],
   alphaCSR[ 182 ][ 251 ],
   alphaCSR[ 182 ][ 252 ],
   alphaCSR[ 182 ][ 253 ],
   alphaCSR[ 182 ][ 254 ],
   alphaCSR[ 182 ][ 255 ],
   alphaCSR[ 182 ][ 256 ],
   alphaCSR[ 182 ][ 257 ],
   alphaCSR[ 182 ][ 258 ],
   alphaCSR[ 182 ][ 259 ],
   alphaCSR[ 182 ][ 260 ],
   alphaCSR[ 182 ][ 261 ],
   alphaCSR[ 182 ][ 262 ],
   alphaCSR[ 182 ][ 263 ],
   alphaCSR[ 182 ][ 264 ],
   alphaCSR[ 182 ][ 265 ],
   alphaCSR[ 182 ][ 266 ],
   alphaCSR[ 182 ][ 267 ],
   alphaCSR[ 182 ][ 268 ],
   alphaCSR[ 182 ][ 269 ],
   alphaCSR[ 182 ][ 270 ],
   alphaCSR[ 182 ][ 271 ],
   alphaCSR[ 182 ][ 272 ],
   alphaCSR[ 182 ][ 273 ],
   alphaCSR[ 182 ][ 274 ],
   alphaCSR[ 182 ][ 275 ],
   alphaCSR[ 182 ][ 276 ],
   alphaCSR[ 182 ][ 277 ],
   alphaCSR[ 182 ][ 278 ],
   alphaCSR[ 182 ][ 279 ],
   alphaCSR[ 182 ][ 280 ],
   alphaCSR[ 182 ][ 281 ],
   alphaCSR[ 182 ][ 282 ],
   alphaCSR[ 182 ][ 283 ],
   alphaCSR[ 182 ][ 284 ],
   alphaCSR[ 182 ][ 285 ],
   alphaCSR[ 182 ][ 286 ],
   alphaCSR[ 182 ][ 287 ],
   alphaCSR[ 182 ][ 288 ],
   alphaCSR[ 182 ][ 289 ],
   alphaCSR[ 182 ][ 290 ],
   alphaCSR[ 182 ][ 291 ],
   alphaCSR[ 182 ][ 292 ],
   alphaCSR[ 182 ][ 293 ],
   alphaCSR[ 182 ][ 294 ],
   alphaCSR[ 182 ][ 295 ],
   alphaCSR[ 182 ][ 296 ],
   alphaCSR[ 182 ][ 297 ],
   alphaCSR[ 182 ][ 298 ],
   alphaCSR[ 182 ][ 299 ],
   alphaCSR[ 182 ][ 300 ],
   alphaCSR[ 182 ][ 301 ],
   alphaCSR[ 182 ][ 302 ],
   alphaCSR[ 182 ][ 303 ],
   alphaCSR[ 182 ][ 304 ],
   alphaCSR[ 182 ][ 305 ],
   alphaCSR[ 182 ][ 306 ],
   alphaCSR[ 182 ][ 307 ],
   alphaCSR[ 182 ][ 308 ],
   alphaCSR[ 182 ][ 309 ],
   alphaCSR[ 182 ][ 310 ],
   alphaCSR[ 182 ][ 311 ],
   alphaCSR[ 182 ][ 312 ],
   alphaCSR[ 182 ][ 313 ],
   alphaCSR[ 182 ][ 314 ],
   alphaCSR[ 182 ][ 315 ],
   alphaCSR[ 182 ][ 316 ],
   alphaCSR[ 182 ][ 317 ],
   alphaCSR[ 182 ][ 318 ],
   alphaCSR[ 182 ][ 319 ],
   alphaCSR[ 182 ][ 320 ],
   alphaCSR[ 182 ][ 321 ],
   alphaCSR[ 182 ][ 322 ],
   alphaCSR[ 182 ][ 323 ],
   alphaCSR[ 182 ][ 324 ],
   alphaCSR[ 182 ][ 325 ],
   alphaCSR[ 182 ][ 326 ],
   alphaCSR[ 182 ][ 327 ],
   alphaCSR[ 182 ][ 328 ],
   alphaCSR[ 182 ][ 329 ],
   alphaCSR[ 182 ][ 330 ],
   alphaCSR[ 182 ][ 331 ],
   alphaCSR[ 182 ][ 332 ],
   alphaCSR[ 182 ][ 333 ],
   alphaCSR[ 182 ][ 334 ],
   alphaCSR[ 182 ][ 335 ],
   alphaCSR[ 182 ][ 336 ],
   alphaCSR[ 182 ][ 337 ],
   alphaCSR[ 182 ][ 338 ],
   alphaCSR[ 182 ][ 339 ],
   alphaCSR[ 182 ][ 340 ],
   alphaCSR[ 182 ][ 341 ],
   alphaCSR[ 182 ][ 342 ],
   alphaCSR[ 182 ][ 343 ],
   alphaCSR[ 182 ][ 344 ],
   alphaCSR[ 182 ][ 345 ],
   alphaCSR[ 182 ][ 346 ],
   alphaCSR[ 182 ][ 347 ],
   alphaCSR[ 182 ][ 348 ],
   alphaCSR[ 182 ][ 349 ],
   alphaCSR[ 182 ][ 350 ],
   alphaCSR[ 182 ][ 351 ],
   alphaCSR[ 182 ][ 352 ],
   alphaCSR[ 182 ][ 353 ],
   alphaCSR[ 182 ][ 354 ],
   alphaCSR[ 182 ][ 355 ],
   alphaCSR[ 182 ][ 356 ],
   alphaCSR[ 182 ][ 357 ],
   alphaCSR[ 182 ][ 358 ],
   alphaCSR[ 182 ][ 359 ],
   alphaCSR[ 182 ][ 360 ],
   alphaCSR[ 182 ][ 361 ],
   alphaCSR[ 182 ][ 362 ],
   alphaCSR[ 182 ][ 363 ],
   alphaCSR[ 182 ][ 364 ],
   alphaCSR[ 182 ][ 365 ],
   alphaCSR[ 182 ][ 366 ],
   alphaCSR[ 182 ][ 367 ],
   alphaCSR[ 182 ][ 368 ],
   alphaCSR[ 182 ][ 369 ],
   alphaCSR[ 182 ][ 370 ],
   alphaCSR[ 182 ][ 371 ],
   alphaCSR[ 182 ][ 372 ],
   alphaCSR[ 182 ][ 373 ],
   alphaCSR[ 182 ][ 374 ],
   alphaCSR[ 182 ][ 375 ],
   alphaCSR[ 182 ][ 376 ],
   alphaCSR[ 182 ][ 377 ],
   alphaCSR[ 182 ][ 378 ],
   alphaCSR[ 182 ][ 379 ],
   alphaCSR[ 182 ][ 380 ],
   alphaCSR[ 182 ][ 381 ],
   alphaCSR[ 182 ][ 382 ],
   alphaCSR[ 182 ][ 383 ],
   alphaCSR[ 183 ][ 0 ],
   alphaCSR[ 183 ][ 1 ],
   alphaCSR[ 183 ][ 2 ],
   alphaCSR[ 183 ][ 3 ],
   alphaCSR[ 183 ][ 4 ],
   alphaCSR[ 183 ][ 5 ],
   alphaCSR[ 183 ][ 6 ],
   alphaCSR[ 183 ][ 7 ],
   alphaCSR[ 183 ][ 8 ],
   alphaCSR[ 183 ][ 9 ],
   alphaCSR[ 183 ][ 10 ],
   alphaCSR[ 183 ][ 11 ],
   alphaCSR[ 183 ][ 12 ],
   alphaCSR[ 183 ][ 13 ],
   alphaCSR[ 183 ][ 14 ],
   alphaCSR[ 183 ][ 15 ],
   alphaCSR[ 183 ][ 16 ],
   alphaCSR[ 183 ][ 17 ],
   alphaCSR[ 183 ][ 18 ],
   alphaCSR[ 183 ][ 19 ],
   alphaCSR[ 183 ][ 20 ],
   alphaCSR[ 183 ][ 21 ],
   alphaCSR[ 183 ][ 22 ],
   alphaCSR[ 183 ][ 23 ],
   alphaCSR[ 183 ][ 24 ],
   alphaCSR[ 183 ][ 25 ],
   alphaCSR[ 183 ][ 26 ],
   alphaCSR[ 183 ][ 27 ],
   alphaCSR[ 183 ][ 28 ],
   alphaCSR[ 183 ][ 29 ],
   alphaCSR[ 183 ][ 30 ],
   alphaCSR[ 183 ][ 31 ],
   alphaCSR[ 183 ][ 32 ],
   alphaCSR[ 183 ][ 33 ],
   alphaCSR[ 183 ][ 34 ],
   alphaCSR[ 183 ][ 35 ],
   alphaCSR[ 183 ][ 36 ],
   alphaCSR[ 183 ][ 37 ],
   alphaCSR[ 183 ][ 38 ],
   alphaCSR[ 183 ][ 39 ],
   alphaCSR[ 183 ][ 40 ],
   alphaCSR[ 183 ][ 41 ],
   alphaCSR[ 183 ][ 42 ],
   alphaCSR[ 183 ][ 43 ],
   alphaCSR[ 183 ][ 44 ],
   alphaCSR[ 183 ][ 45 ],
   alphaCSR[ 183 ][ 46 ],
   alphaCSR[ 183 ][ 47 ],
   alphaCSR[ 183 ][ 48 ],
   alphaCSR[ 183 ][ 49 ],
   alphaCSR[ 183 ][ 50 ],
   alphaCSR[ 183 ][ 51 ],
   alphaCSR[ 183 ][ 52 ],
   alphaCSR[ 183 ][ 53 ],
   alphaCSR[ 183 ][ 54 ],
   alphaCSR[ 183 ][ 55 ],
   alphaCSR[ 183 ][ 56 ],
   alphaCSR[ 183 ][ 57 ],
   alphaCSR[ 183 ][ 58 ],
   alphaCSR[ 183 ][ 59 ],
   alphaCSR[ 183 ][ 60 ],
   alphaCSR[ 183 ][ 61 ],
   alphaCSR[ 183 ][ 62 ],
   alphaCSR[ 183 ][ 63 ],
   alphaCSR[ 183 ][ 64 ],
   alphaCSR[ 183 ][ 65 ],
   alphaCSR[ 183 ][ 66 ],
   alphaCSR[ 183 ][ 67 ],
   alphaCSR[ 183 ][ 68 ],
   alphaCSR[ 183 ][ 69 ],
   alphaCSR[ 183 ][ 70 ],
   alphaCSR[ 183 ][ 71 ],
   alphaCSR[ 183 ][ 72 ],
   alphaCSR[ 183 ][ 73 ],
   alphaCSR[ 183 ][ 74 ],
   alphaCSR[ 183 ][ 75 ],
   alphaCSR[ 183 ][ 76 ],
   alphaCSR[ 183 ][ 77 ],
   alphaCSR[ 183 ][ 78 ],
   alphaCSR[ 183 ][ 79 ],
   alphaCSR[ 183 ][ 80 ],
   alphaCSR[ 183 ][ 81 ],
   alphaCSR[ 183 ][ 82 ],
   alphaCSR[ 183 ][ 83 ],
   alphaCSR[ 183 ][ 84 ],
   alphaCSR[ 183 ][ 85 ],
   alphaCSR[ 183 ][ 86 ],
   alphaCSR[ 183 ][ 87 ],
   alphaCSR[ 183 ][ 88 ],
   alphaCSR[ 183 ][ 89 ],
   alphaCSR[ 183 ][ 90 ],
   alphaCSR[ 183 ][ 91 ],
   alphaCSR[ 183 ][ 92 ],
   alphaCSR[ 183 ][ 93 ],
   alphaCSR[ 183 ][ 94 ],
   alphaCSR[ 183 ][ 95 ],
   alphaCSR[ 183 ][ 96 ],
   alphaCSR[ 183 ][ 97 ],
   alphaCSR[ 183 ][ 98 ],
   alphaCSR[ 183 ][ 99 ],
   alphaCSR[ 183 ][ 100 ],
   alphaCSR[ 183 ][ 101 ],
   alphaCSR[ 183 ][ 102 ],
   alphaCSR[ 183 ][ 103 ],
   alphaCSR[ 183 ][ 104 ],
   alphaCSR[ 183 ][ 105 ],
   alphaCSR[ 183 ][ 106 ],
   alphaCSR[ 183 ][ 107 ],
   alphaCSR[ 183 ][ 108 ],
   alphaCSR[ 183 ][ 109 ],
   alphaCSR[ 183 ][ 110 ],
   alphaCSR[ 183 ][ 111 ],
   alphaCSR[ 183 ][ 112 ],
   alphaCSR[ 183 ][ 113 ],
   alphaCSR[ 183 ][ 114 ],
   alphaCSR[ 183 ][ 115 ],
   alphaCSR[ 183 ][ 116 ],
   alphaCSR[ 183 ][ 117 ],
   alphaCSR[ 183 ][ 118 ],
   alphaCSR[ 183 ][ 119 ],
   alphaCSR[ 183 ][ 120 ],
   alphaCSR[ 183 ][ 121 ],
   alphaCSR[ 183 ][ 122 ],
   alphaCSR[ 183 ][ 123 ],
   alphaCSR[ 183 ][ 124 ],
   alphaCSR[ 183 ][ 125 ],
   alphaCSR[ 183 ][ 126 ],
   alphaCSR[ 183 ][ 127 ],
   alphaCSR[ 183 ][ 128 ],
   alphaCSR[ 183 ][ 129 ],
   alphaCSR[ 183 ][ 130 ],
   alphaCSR[ 183 ][ 131 ],
   alphaCSR[ 183 ][ 132 ],
   alphaCSR[ 183 ][ 133 ],
   alphaCSR[ 183 ][ 134 ],
   alphaCSR[ 183 ][ 135 ],
   alphaCSR[ 183 ][ 136 ],
   alphaCSR[ 183 ][ 137 ],
   alphaCSR[ 183 ][ 138 ],
   alphaCSR[ 183 ][ 139 ],
   alphaCSR[ 183 ][ 140 ],
   alphaCSR[ 183 ][ 141 ],
   alphaCSR[ 183 ][ 142 ],
   alphaCSR[ 183 ][ 143 ],
   alphaCSR[ 183 ][ 144 ],
   alphaCSR[ 183 ][ 145 ],
   alphaCSR[ 183 ][ 146 ],
   alphaCSR[ 183 ][ 147 ],
   alphaCSR[ 183 ][ 148 ],
   alphaCSR[ 183 ][ 149 ],
   alphaCSR[ 183 ][ 150 ],
   alphaCSR[ 183 ][ 151 ],
   alphaCSR[ 183 ][ 152 ],
   alphaCSR[ 183 ][ 153 ],
   alphaCSR[ 183 ][ 154 ],
   alphaCSR[ 183 ][ 155 ],
   alphaCSR[ 183 ][ 156 ],
   alphaCSR[ 183 ][ 157 ],
   alphaCSR[ 183 ][ 158 ],
   alphaCSR[ 183 ][ 159 ],
   alphaCSR[ 183 ][ 160 ],
   alphaCSR[ 183 ][ 161 ],
   alphaCSR[ 183 ][ 162 ],
   alphaCSR[ 183 ][ 163 ],
   alphaCSR[ 183 ][ 164 ],
   alphaCSR[ 183 ][ 165 ],
   alphaCSR[ 183 ][ 166 ],
   alphaCSR[ 183 ][ 167 ],
   alphaCSR[ 183 ][ 168 ],
   alphaCSR[ 183 ][ 169 ],
   alphaCSR[ 183 ][ 170 ],
   alphaCSR[ 183 ][ 171 ],
   alphaCSR[ 183 ][ 172 ],
   alphaCSR[ 183 ][ 173 ],
   alphaCSR[ 183 ][ 174 ],
   alphaCSR[ 183 ][ 175 ],
   alphaCSR[ 183 ][ 176 ],
   alphaCSR[ 183 ][ 177 ],
   alphaCSR[ 183 ][ 178 ],
   alphaCSR[ 183 ][ 179 ],
   alphaCSR[ 183 ][ 180 ],
   alphaCSR[ 183 ][ 181 ],
   alphaCSR[ 183 ][ 182 ],
   alphaCSR[ 183 ][ 183 ],
   alphaCSR[ 183 ][ 184 ],
   alphaCSR[ 183 ][ 185 ],
   alphaCSR[ 183 ][ 186 ],
   alphaCSR[ 183 ][ 187 ],
   alphaCSR[ 183 ][ 188 ],
   alphaCSR[ 183 ][ 189 ],
   alphaCSR[ 183 ][ 190 ],
   alphaCSR[ 183 ][ 191 ],
   alphaCSR[ 183 ][ 192 ],
   alphaCSR[ 183 ][ 193 ],
   alphaCSR[ 183 ][ 194 ],
   alphaCSR[ 183 ][ 195 ],
   alphaCSR[ 183 ][ 196 ],
   alphaCSR[ 183 ][ 197 ],
   alphaCSR[ 183 ][ 198 ],
   alphaCSR[ 183 ][ 199 ],
   alphaCSR[ 183 ][ 200 ],
   alphaCSR[ 183 ][ 201 ],
   alphaCSR[ 183 ][ 202 ],
   alphaCSR[ 183 ][ 203 ],
   alphaCSR[ 183 ][ 204 ],
   alphaCSR[ 183 ][ 205 ],
   alphaCSR[ 183 ][ 206 ],
   alphaCSR[ 183 ][ 207 ],
   alphaCSR[ 183 ][ 208 ],
   alphaCSR[ 183 ][ 209 ],
   alphaCSR[ 183 ][ 210 ],
   alphaCSR[ 183 ][ 211 ],
   alphaCSR[ 183 ][ 212 ],
   alphaCSR[ 183 ][ 213 ],
   alphaCSR[ 183 ][ 214 ],
   alphaCSR[ 183 ][ 215 ],
   alphaCSR[ 183 ][ 216 ],
   alphaCSR[ 183 ][ 217 ],
   alphaCSR[ 183 ][ 218 ],
   alphaCSR[ 183 ][ 219 ],
   alphaCSR[ 183 ][ 220 ],
   alphaCSR[ 183 ][ 221 ],
   alphaCSR[ 183 ][ 222 ],
   alphaCSR[ 183 ][ 223 ],
   alphaCSR[ 183 ][ 224 ],
   alphaCSR[ 183 ][ 225 ],
   alphaCSR[ 183 ][ 226 ],
   alphaCSR[ 183 ][ 227 ],
   alphaCSR[ 183 ][ 228 ],
   alphaCSR[ 183 ][ 229 ],
   alphaCSR[ 183 ][ 230 ],
   alphaCSR[ 183 ][ 231 ],
   alphaCSR[ 183 ][ 232 ],
   alphaCSR[ 183 ][ 233 ],
   alphaCSR[ 183 ][ 234 ],
   alphaCSR[ 183 ][ 235 ],
   alphaCSR[ 183 ][ 236 ],
   alphaCSR[ 183 ][ 237 ],
   alphaCSR[ 183 ][ 238 ],
   alphaCSR[ 183 ][ 239 ],
   alphaCSR[ 183 ][ 240 ],
   alphaCSR[ 183 ][ 241 ],
   alphaCSR[ 183 ][ 242 ],
   alphaCSR[ 183 ][ 243 ],
   alphaCSR[ 183 ][ 244 ],
   alphaCSR[ 183 ][ 245 ],
   alphaCSR[ 183 ][ 246 ],
   alphaCSR[ 183 ][ 247 ],
   alphaCSR[ 183 ][ 248 ],
   alphaCSR[ 183 ][ 249 ],
   alphaCSR[ 183 ][ 250 ],
   alphaCSR[ 183 ][ 251 ],
   alphaCSR[ 183 ][ 252 ],
   alphaCSR[ 183 ][ 253 ],
   alphaCSR[ 183 ][ 254 ],
   alphaCSR[ 183 ][ 255 ],
   alphaCSR[ 183 ][ 256 ],
   alphaCSR[ 183 ][ 257 ],
   alphaCSR[ 183 ][ 258 ],
   alphaCSR[ 183 ][ 259 ],
   alphaCSR[ 183 ][ 260 ],
   alphaCSR[ 183 ][ 261 ],
   alphaCSR[ 183 ][ 262 ],
   alphaCSR[ 183 ][ 263 ],
   alphaCSR[ 183 ][ 264 ],
   alphaCSR[ 183 ][ 265 ],
   alphaCSR[ 183 ][ 266 ],
   alphaCSR[ 183 ][ 267 ],
   alphaCSR[ 183 ][ 268 ],
   alphaCSR[ 183 ][ 269 ],
   alphaCSR[ 183 ][ 270 ],
   alphaCSR[ 183 ][ 271 ],
   alphaCSR[ 183 ][ 272 ],
   alphaCSR[ 183 ][ 273 ],
   alphaCSR[ 183 ][ 274 ],
   alphaCSR[ 183 ][ 275 ],
   alphaCSR[ 183 ][ 276 ],
   alphaCSR[ 183 ][ 277 ],
   alphaCSR[ 183 ][ 278 ],
   alphaCSR[ 183 ][ 279 ],
   alphaCSR[ 183 ][ 280 ],
   alphaCSR[ 183 ][ 281 ],
   alphaCSR[ 183 ][ 282 ],
   alphaCSR[ 183 ][ 283 ],
   alphaCSR[ 183 ][ 284 ],
   alphaCSR[ 183 ][ 285 ],
   alphaCSR[ 183 ][ 286 ],
   alphaCSR[ 183 ][ 287 ],
   alphaCSR[ 183 ][ 288 ],
   alphaCSR[ 183 ][ 289 ],
   alphaCSR[ 183 ][ 290 ],
   alphaCSR[ 183 ][ 291 ],
   alphaCSR[ 183 ][ 292 ],
   alphaCSR[ 183 ][ 293 ],
   alphaCSR[ 183 ][ 294 ],
   alphaCSR[ 183 ][ 295 ],
   alphaCSR[ 183 ][ 296 ],
   alphaCSR[ 183 ][ 297 ],
   alphaCSR[ 183 ][ 298 ],
   alphaCSR[ 183 ][ 299 ],
   alphaCSR[ 183 ][ 300 ],
   alphaCSR[ 183 ][ 301 ],
   alphaCSR[ 183 ][ 302 ],
   alphaCSR[ 183 ][ 303 ],
   alphaCSR[ 183 ][ 304 ],
   alphaCSR[ 183 ][ 305 ],
   alphaCSR[ 183 ][ 306 ],
   alphaCSR[ 183 ][ 307 ],
   alphaCSR[ 183 ][ 308 ],
   alphaCSR[ 183 ][ 309 ],
   alphaCSR[ 183 ][ 310 ],
   alphaCSR[ 183 ][ 311 ],
   alphaCSR[ 183 ][ 312 ],
   alphaCSR[ 183 ][ 313 ],
   alphaCSR[ 183 ][ 314 ],
   alphaCSR[ 183 ][ 315 ],
   alphaCSR[ 183 ][ 316 ],
   alphaCSR[ 183 ][ 317 ],
   alphaCSR[ 183 ][ 318 ],
   alphaCSR[ 183 ][ 319 ],
   alphaCSR[ 183 ][ 320 ],
   alphaCSR[ 183 ][ 321 ],
   alphaCSR[ 183 ][ 322 ],
   alphaCSR[ 183 ][ 323 ],
   alphaCSR[ 183 ][ 324 ],
   alphaCSR[ 183 ][ 325 ],
   alphaCSR[ 183 ][ 326 ],
   alphaCSR[ 183 ][ 327 ],
   alphaCSR[ 183 ][ 328 ],
   alphaCSR[ 183 ][ 329 ],
   alphaCSR[ 183 ][ 330 ],
   alphaCSR[ 183 ][ 331 ],
   alphaCSR[ 183 ][ 332 ],
   alphaCSR[ 183 ][ 333 ],
   alphaCSR[ 183 ][ 334 ],
   alphaCSR[ 183 ][ 335 ],
   alphaCSR[ 183 ][ 336 ],
   alphaCSR[ 183 ][ 337 ],
   alphaCSR[ 183 ][ 338 ],
   alphaCSR[ 183 ][ 339 ],
   alphaCSR[ 183 ][ 340 ],
   alphaCSR[ 183 ][ 341 ],
   alphaCSR[ 183 ][ 342 ],
   alphaCSR[ 183 ][ 343 ],
   alphaCSR[ 183 ][ 344 ],
   alphaCSR[ 183 ][ 345 ],
   alphaCSR[ 183 ][ 346 ],
   alphaCSR[ 183 ][ 347 ],
   alphaCSR[ 183 ][ 348 ],
   alphaCSR[ 183 ][ 349 ],
   alphaCSR[ 183 ][ 350 ],
   alphaCSR[ 183 ][ 351 ],
   alphaCSR[ 183 ][ 352 ],
   alphaCSR[ 183 ][ 353 ],
   alphaCSR[ 183 ][ 354 ],
   alphaCSR[ 183 ][ 355 ],
   alphaCSR[ 183 ][ 356 ],
   alphaCSR[ 183 ][ 357 ],
   alphaCSR[ 183 ][ 358 ],
   alphaCSR[ 183 ][ 359 ],
   alphaCSR[ 183 ][ 360 ],
   alphaCSR[ 183 ][ 361 ],
   alphaCSR[ 183 ][ 362 ],
   alphaCSR[ 183 ][ 363 ],
   alphaCSR[ 183 ][ 364 ],
   alphaCSR[ 183 ][ 365 ],
   alphaCSR[ 183 ][ 366 ],
   alphaCSR[ 183 ][ 367 ],
   alphaCSR[ 183 ][ 368 ],
   alphaCSR[ 183 ][ 369 ],
   alphaCSR[ 183 ][ 370 ],
   alphaCSR[ 183 ][ 371 ],
   alphaCSR[ 183 ][ 372 ],
   alphaCSR[ 183 ][ 373 ],
   alphaCSR[ 183 ][ 374 ],
   alphaCSR[ 183 ][ 375 ],
   alphaCSR[ 183 ][ 376 ],
   alphaCSR[ 183 ][ 377 ],
   alphaCSR[ 183 ][ 378 ],
   alphaCSR[ 183 ][ 379 ],
   alphaCSR[ 183 ][ 380 ],
   alphaCSR[ 183 ][ 381 ],
   alphaCSR[ 183 ][ 382 ],
   alphaCSR[ 183 ][ 383 ],
   alphaCSR[ 184 ][ 0 ],
   alphaCSR[ 184 ][ 1 ],
   alphaCSR[ 184 ][ 2 ],
   alphaCSR[ 184 ][ 3 ],
   alphaCSR[ 184 ][ 4 ],
   alphaCSR[ 184 ][ 5 ],
   alphaCSR[ 184 ][ 6 ],
   alphaCSR[ 184 ][ 7 ],
   alphaCSR[ 184 ][ 8 ],
   alphaCSR[ 184 ][ 9 ],
   alphaCSR[ 184 ][ 10 ],
   alphaCSR[ 184 ][ 11 ],
   alphaCSR[ 184 ][ 12 ],
   alphaCSR[ 184 ][ 13 ],
   alphaCSR[ 184 ][ 14 ],
   alphaCSR[ 184 ][ 15 ],
   alphaCSR[ 184 ][ 16 ],
   alphaCSR[ 184 ][ 17 ],
   alphaCSR[ 184 ][ 18 ],
   alphaCSR[ 184 ][ 19 ],
   alphaCSR[ 184 ][ 20 ],
   alphaCSR[ 184 ][ 21 ],
   alphaCSR[ 184 ][ 22 ],
   alphaCSR[ 184 ][ 23 ],
   alphaCSR[ 184 ][ 24 ],
   alphaCSR[ 184 ][ 25 ],
   alphaCSR[ 184 ][ 26 ],
   alphaCSR[ 184 ][ 27 ],
   alphaCSR[ 184 ][ 28 ],
   alphaCSR[ 184 ][ 29 ],
   alphaCSR[ 184 ][ 30 ],
   alphaCSR[ 184 ][ 31 ],
   alphaCSR[ 184 ][ 32 ],
   alphaCSR[ 184 ][ 33 ],
   alphaCSR[ 184 ][ 34 ],
   alphaCSR[ 184 ][ 35 ],
   alphaCSR[ 184 ][ 36 ],
   alphaCSR[ 184 ][ 37 ],
   alphaCSR[ 184 ][ 38 ],
   alphaCSR[ 184 ][ 39 ],
   alphaCSR[ 184 ][ 40 ],
   alphaCSR[ 184 ][ 41 ],
   alphaCSR[ 184 ][ 42 ],
   alphaCSR[ 184 ][ 43 ],
   alphaCSR[ 184 ][ 44 ],
   alphaCSR[ 184 ][ 45 ],
   alphaCSR[ 184 ][ 46 ],
   alphaCSR[ 184 ][ 47 ],
   alphaCSR[ 184 ][ 48 ],
   alphaCSR[ 184 ][ 49 ],
   alphaCSR[ 184 ][ 50 ],
   alphaCSR[ 184 ][ 51 ],
   alphaCSR[ 184 ][ 52 ],
   alphaCSR[ 184 ][ 53 ],
   alphaCSR[ 184 ][ 54 ],
   alphaCSR[ 184 ][ 55 ],
   alphaCSR[ 184 ][ 56 ],
   alphaCSR[ 184 ][ 57 ],
   alphaCSR[ 184 ][ 58 ],
   alphaCSR[ 184 ][ 59 ],
   alphaCSR[ 184 ][ 60 ],
   alphaCSR[ 184 ][ 61 ],
   alphaCSR[ 184 ][ 62 ],
   alphaCSR[ 184 ][ 63 ],
   alphaCSR[ 184 ][ 64 ],
   alphaCSR[ 184 ][ 65 ],
   alphaCSR[ 184 ][ 66 ],
   alphaCSR[ 184 ][ 67 ],
   alphaCSR[ 184 ][ 68 ],
   alphaCSR[ 184 ][ 69 ],
   alphaCSR[ 184 ][ 70 ],
   alphaCSR[ 184 ][ 71 ],
   alphaCSR[ 184 ][ 72 ],
   alphaCSR[ 184 ][ 73 ],
   alphaCSR[ 184 ][ 74 ],
   alphaCSR[ 184 ][ 75 ],
   alphaCSR[ 184 ][ 76 ],
   alphaCSR[ 184 ][ 77 ],
   alphaCSR[ 184 ][ 78 ],
   alphaCSR[ 184 ][ 79 ],
   alphaCSR[ 184 ][ 80 ],
   alphaCSR[ 184 ][ 81 ],
   alphaCSR[ 184 ][ 82 ],
   alphaCSR[ 184 ][ 83 ],
   alphaCSR[ 184 ][ 84 ],
   alphaCSR[ 184 ][ 85 ],
   alphaCSR[ 184 ][ 86 ],
   alphaCSR[ 184 ][ 87 ],
   alphaCSR[ 184 ][ 88 ],
   alphaCSR[ 184 ][ 89 ],
   alphaCSR[ 184 ][ 90 ],
   alphaCSR[ 184 ][ 91 ],
   alphaCSR[ 184 ][ 92 ],
   alphaCSR[ 184 ][ 93 ],
   alphaCSR[ 184 ][ 94 ],
   alphaCSR[ 184 ][ 95 ],
   alphaCSR[ 184 ][ 96 ],
   alphaCSR[ 184 ][ 97 ],
   alphaCSR[ 184 ][ 98 ],
   alphaCSR[ 184 ][ 99 ],
   alphaCSR[ 184 ][ 100 ],
   alphaCSR[ 184 ][ 101 ],
   alphaCSR[ 184 ][ 102 ],
   alphaCSR[ 184 ][ 103 ],
   alphaCSR[ 184 ][ 104 ],
   alphaCSR[ 184 ][ 105 ],
   alphaCSR[ 184 ][ 106 ],
   alphaCSR[ 184 ][ 107 ],
   alphaCSR[ 184 ][ 108 ],
   alphaCSR[ 184 ][ 109 ],
   alphaCSR[ 184 ][ 110 ],
   alphaCSR[ 184 ][ 111 ],
   alphaCSR[ 184 ][ 112 ],
   alphaCSR[ 184 ][ 113 ],
   alphaCSR[ 184 ][ 114 ],
   alphaCSR[ 184 ][ 115 ],
   alphaCSR[ 184 ][ 116 ],
   alphaCSR[ 184 ][ 117 ],
   alphaCSR[ 184 ][ 118 ],
   alphaCSR[ 184 ][ 119 ],
   alphaCSR[ 184 ][ 120 ],
   alphaCSR[ 184 ][ 121 ],
   alphaCSR[ 184 ][ 122 ],
   alphaCSR[ 184 ][ 123 ],
   alphaCSR[ 184 ][ 124 ],
   alphaCSR[ 184 ][ 125 ],
   alphaCSR[ 184 ][ 126 ],
   alphaCSR[ 184 ][ 127 ],
   alphaCSR[ 184 ][ 128 ],
   alphaCSR[ 184 ][ 129 ],
   alphaCSR[ 184 ][ 130 ],
   alphaCSR[ 184 ][ 131 ],
   alphaCSR[ 184 ][ 132 ],
   alphaCSR[ 184 ][ 133 ],
   alphaCSR[ 184 ][ 134 ],
   alphaCSR[ 184 ][ 135 ],
   alphaCSR[ 184 ][ 136 ],
   alphaCSR[ 184 ][ 137 ],
   alphaCSR[ 184 ][ 138 ],
   alphaCSR[ 184 ][ 139 ],
   alphaCSR[ 184 ][ 140 ],
   alphaCSR[ 184 ][ 141 ],
   alphaCSR[ 184 ][ 142 ],
   alphaCSR[ 184 ][ 143 ],
   alphaCSR[ 184 ][ 144 ],
   alphaCSR[ 184 ][ 145 ],
   alphaCSR[ 184 ][ 146 ],
   alphaCSR[ 184 ][ 147 ],
   alphaCSR[ 184 ][ 148 ],
   alphaCSR[ 184 ][ 149 ],
   alphaCSR[ 184 ][ 150 ],
   alphaCSR[ 184 ][ 151 ],
   alphaCSR[ 184 ][ 152 ],
   alphaCSR[ 184 ][ 153 ],
   alphaCSR[ 184 ][ 154 ],
   alphaCSR[ 184 ][ 155 ],
   alphaCSR[ 184 ][ 156 ],
   alphaCSR[ 184 ][ 157 ],
   alphaCSR[ 184 ][ 158 ],
   alphaCSR[ 184 ][ 159 ],
   alphaCSR[ 184 ][ 160 ],
   alphaCSR[ 184 ][ 161 ],
   alphaCSR[ 184 ][ 162 ],
   alphaCSR[ 184 ][ 163 ],
   alphaCSR[ 184 ][ 164 ],
   alphaCSR[ 184 ][ 165 ],
   alphaCSR[ 184 ][ 166 ],
   alphaCSR[ 184 ][ 167 ],
   alphaCSR[ 184 ][ 168 ],
   alphaCSR[ 184 ][ 169 ],
   alphaCSR[ 184 ][ 170 ],
   alphaCSR[ 184 ][ 171 ],
   alphaCSR[ 184 ][ 172 ],
   alphaCSR[ 184 ][ 173 ],
   alphaCSR[ 184 ][ 174 ],
   alphaCSR[ 184 ][ 175 ],
   alphaCSR[ 184 ][ 176 ],
   alphaCSR[ 184 ][ 177 ],
   alphaCSR[ 184 ][ 178 ],
   alphaCSR[ 184 ][ 179 ],
   alphaCSR[ 184 ][ 180 ],
   alphaCSR[ 184 ][ 181 ],
   alphaCSR[ 184 ][ 182 ],
   alphaCSR[ 184 ][ 183 ],
   alphaCSR[ 184 ][ 184 ],
   alphaCSR[ 184 ][ 185 ],
   alphaCSR[ 184 ][ 186 ],
   alphaCSR[ 184 ][ 187 ],
   alphaCSR[ 184 ][ 188 ],
   alphaCSR[ 184 ][ 189 ],
   alphaCSR[ 184 ][ 190 ],
   alphaCSR[ 184 ][ 191 ],
   alphaCSR[ 184 ][ 192 ],
   alphaCSR[ 184 ][ 193 ],
   alphaCSR[ 184 ][ 194 ],
   alphaCSR[ 184 ][ 195 ],
   alphaCSR[ 184 ][ 196 ],
   alphaCSR[ 184 ][ 197 ],
   alphaCSR[ 184 ][ 198 ],
   alphaCSR[ 184 ][ 199 ],
   alphaCSR[ 184 ][ 200 ],
   alphaCSR[ 184 ][ 201 ],
   alphaCSR[ 184 ][ 202 ],
   alphaCSR[ 184 ][ 203 ],
   alphaCSR[ 184 ][ 204 ],
   alphaCSR[ 184 ][ 205 ],
   alphaCSR[ 184 ][ 206 ],
   alphaCSR[ 184 ][ 207 ],
   alphaCSR[ 184 ][ 208 ],
   alphaCSR[ 184 ][ 209 ],
   alphaCSR[ 184 ][ 210 ],
   alphaCSR[ 184 ][ 211 ],
   alphaCSR[ 184 ][ 212 ],
   alphaCSR[ 184 ][ 213 ],
   alphaCSR[ 184 ][ 214 ],
   alphaCSR[ 184 ][ 215 ],
   alphaCSR[ 184 ][ 216 ],
   alphaCSR[ 184 ][ 217 ],
   alphaCSR[ 184 ][ 218 ],
   alphaCSR[ 184 ][ 219 ],
   alphaCSR[ 184 ][ 220 ],
   alphaCSR[ 184 ][ 221 ],
   alphaCSR[ 184 ][ 222 ],
   alphaCSR[ 184 ][ 223 ],
   alphaCSR[ 184 ][ 224 ],
   alphaCSR[ 184 ][ 225 ],
   alphaCSR[ 184 ][ 226 ],
   alphaCSR[ 184 ][ 227 ],
   alphaCSR[ 184 ][ 228 ],
   alphaCSR[ 184 ][ 229 ],
   alphaCSR[ 184 ][ 230 ],
   alphaCSR[ 184 ][ 231 ],
   alphaCSR[ 184 ][ 232 ],
   alphaCSR[ 184 ][ 233 ],
   alphaCSR[ 184 ][ 234 ],
   alphaCSR[ 184 ][ 235 ],
   alphaCSR[ 184 ][ 236 ],
   alphaCSR[ 184 ][ 237 ],
   alphaCSR[ 184 ][ 238 ],
   alphaCSR[ 184 ][ 239 ],
   alphaCSR[ 184 ][ 240 ],
   alphaCSR[ 184 ][ 241 ],
   alphaCSR[ 184 ][ 242 ],
   alphaCSR[ 184 ][ 243 ],
   alphaCSR[ 184 ][ 244 ],
   alphaCSR[ 184 ][ 245 ],
   alphaCSR[ 184 ][ 246 ],
   alphaCSR[ 184 ][ 247 ],
   alphaCSR[ 184 ][ 248 ],
   alphaCSR[ 184 ][ 249 ],
   alphaCSR[ 184 ][ 250 ],
   alphaCSR[ 184 ][ 251 ],
   alphaCSR[ 184 ][ 252 ],
   alphaCSR[ 184 ][ 253 ],
   alphaCSR[ 184 ][ 254 ],
   alphaCSR[ 184 ][ 255 ],
   alphaCSR[ 184 ][ 256 ],
   alphaCSR[ 184 ][ 257 ],
   alphaCSR[ 184 ][ 258 ],
   alphaCSR[ 184 ][ 259 ],
   alphaCSR[ 184 ][ 260 ],
   alphaCSR[ 184 ][ 261 ],
   alphaCSR[ 184 ][ 262 ],
   alphaCSR[ 184 ][ 263 ],
   alphaCSR[ 184 ][ 264 ],
   alphaCSR[ 184 ][ 265 ],
   alphaCSR[ 184 ][ 266 ],
   alphaCSR[ 184 ][ 267 ],
   alphaCSR[ 184 ][ 268 ],
   alphaCSR[ 184 ][ 269 ],
   alphaCSR[ 184 ][ 270 ],
   alphaCSR[ 184 ][ 271 ],
   alphaCSR[ 184 ][ 272 ],
   alphaCSR[ 184 ][ 273 ],
   alphaCSR[ 184 ][ 274 ],
   alphaCSR[ 184 ][ 275 ],
   alphaCSR[ 184 ][ 276 ],
   alphaCSR[ 184 ][ 277 ],
   alphaCSR[ 184 ][ 278 ],
   alphaCSR[ 184 ][ 279 ],
   alphaCSR[ 184 ][ 280 ],
   alphaCSR[ 184 ][ 281 ],
   alphaCSR[ 184 ][ 282 ],
   alphaCSR[ 184 ][ 283 ],
   alphaCSR[ 184 ][ 284 ],
   alphaCSR[ 184 ][ 285 ],
   alphaCSR[ 184 ][ 286 ],
   alphaCSR[ 184 ][ 287 ],
   alphaCSR[ 184 ][ 288 ],
   alphaCSR[ 184 ][ 289 ],
   alphaCSR[ 184 ][ 290 ],
   alphaCSR[ 184 ][ 291 ],
   alphaCSR[ 184 ][ 292 ],
   alphaCSR[ 184 ][ 293 ],
   alphaCSR[ 184 ][ 294 ],
   alphaCSR[ 184 ][ 295 ],
   alphaCSR[ 184 ][ 296 ],
   alphaCSR[ 184 ][ 297 ],
   alphaCSR[ 184 ][ 298 ],
   alphaCSR[ 184 ][ 299 ],
   alphaCSR[ 184 ][ 300 ],
   alphaCSR[ 184 ][ 301 ],
   alphaCSR[ 184 ][ 302 ],
   alphaCSR[ 184 ][ 303 ],
   alphaCSR[ 184 ][ 304 ],
   alphaCSR[ 184 ][ 305 ],
   alphaCSR[ 184 ][ 306 ],
   alphaCSR[ 184 ][ 307 ],
   alphaCSR[ 184 ][ 308 ],
   alphaCSR[ 184 ][ 309 ],
   alphaCSR[ 184 ][ 310 ],
   alphaCSR[ 184 ][ 311 ],
   alphaCSR[ 184 ][ 312 ],
   alphaCSR[ 184 ][ 313 ],
   alphaCSR[ 184 ][ 314 ],
   alphaCSR[ 184 ][ 315 ],
   alphaCSR[ 184 ][ 316 ],
   alphaCSR[ 184 ][ 317 ],
   alphaCSR[ 184 ][ 318 ],
   alphaCSR[ 184 ][ 319 ],
   alphaCSR[ 184 ][ 320 ],
   alphaCSR[ 184 ][ 321 ],
   alphaCSR[ 184 ][ 322 ],
   alphaCSR[ 184 ][ 323 ],
   alphaCSR[ 184 ][ 324 ],
   alphaCSR[ 184 ][ 325 ],
   alphaCSR[ 184 ][ 326 ],
   alphaCSR[ 184 ][ 327 ],
   alphaCSR[ 184 ][ 328 ],
   alphaCSR[ 184 ][ 329 ],
   alphaCSR[ 184 ][ 330 ],
   alphaCSR[ 184 ][ 331 ],
   alphaCSR[ 184 ][ 332 ],
   alphaCSR[ 184 ][ 333 ],
   alphaCSR[ 184 ][ 334 ],
   alphaCSR[ 184 ][ 335 ],
   alphaCSR[ 184 ][ 336 ],
   alphaCSR[ 184 ][ 337 ],
   alphaCSR[ 184 ][ 338 ],
   alphaCSR[ 184 ][ 339 ],
   alphaCSR[ 184 ][ 340 ],
   alphaCSR[ 184 ][ 341 ],
   alphaCSR[ 184 ][ 342 ],
   alphaCSR[ 184 ][ 343 ],
   alphaCSR[ 184 ][ 344 ],
   alphaCSR[ 184 ][ 345 ],
   alphaCSR[ 184 ][ 346 ],
   alphaCSR[ 184 ][ 347 ],
   alphaCSR[ 184 ][ 348 ],
   alphaCSR[ 184 ][ 349 ],
   alphaCSR[ 184 ][ 350 ],
   alphaCSR[ 184 ][ 351 ],
   alphaCSR[ 184 ][ 352 ],
   alphaCSR[ 184 ][ 353 ],
   alphaCSR[ 184 ][ 354 ],
   alphaCSR[ 184 ][ 355 ],
   alphaCSR[ 184 ][ 356 ],
   alphaCSR[ 184 ][ 357 ],
   alphaCSR[ 184 ][ 358 ],
   alphaCSR[ 184 ][ 359 ],
   alphaCSR[ 184 ][ 360 ],
   alphaCSR[ 184 ][ 361 ],
   alphaCSR[ 184 ][ 362 ],
   alphaCSR[ 184 ][ 363 ],
   alphaCSR[ 184 ][ 364 ],
   alphaCSR[ 184 ][ 365 ],
   alphaCSR[ 184 ][ 366 ],
   alphaCSR[ 184 ][ 367 ],
   alphaCSR[ 184 ][ 368 ],
   alphaCSR[ 184 ][ 369 ],
   alphaCSR[ 184 ][ 370 ],
   alphaCSR[ 184 ][ 371 ],
   alphaCSR[ 184 ][ 372 ],
   alphaCSR[ 184 ][ 373 ],
   alphaCSR[ 184 ][ 374 ],
   alphaCSR[ 184 ][ 375 ],
   alphaCSR[ 184 ][ 376 ],
   alphaCSR[ 184 ][ 377 ],
   alphaCSR[ 184 ][ 378 ],
   alphaCSR[ 184 ][ 379 ],
   alphaCSR[ 184 ][ 380 ],
   alphaCSR[ 184 ][ 381 ],
   alphaCSR[ 184 ][ 382 ],
   alphaCSR[ 184 ][ 383 ],
   alphaCSR[ 185 ][ 0 ],
   alphaCSR[ 185 ][ 1 ],
   alphaCSR[ 185 ][ 2 ],
   alphaCSR[ 185 ][ 3 ],
   alphaCSR[ 185 ][ 4 ],
   alphaCSR[ 185 ][ 5 ],
   alphaCSR[ 185 ][ 6 ],
   alphaCSR[ 185 ][ 7 ],
   alphaCSR[ 185 ][ 8 ],
   alphaCSR[ 185 ][ 9 ],
   alphaCSR[ 185 ][ 10 ],
   alphaCSR[ 185 ][ 11 ],
   alphaCSR[ 185 ][ 12 ],
   alphaCSR[ 185 ][ 13 ],
   alphaCSR[ 185 ][ 14 ],
   alphaCSR[ 185 ][ 15 ],
   alphaCSR[ 185 ][ 16 ],
   alphaCSR[ 185 ][ 17 ],
   alphaCSR[ 185 ][ 18 ],
   alphaCSR[ 185 ][ 19 ],
   alphaCSR[ 185 ][ 20 ],
   alphaCSR[ 185 ][ 21 ],
   alphaCSR[ 185 ][ 22 ],
   alphaCSR[ 185 ][ 23 ],
   alphaCSR[ 185 ][ 24 ],
   alphaCSR[ 185 ][ 25 ],
   alphaCSR[ 185 ][ 26 ],
   alphaCSR[ 185 ][ 27 ],
   alphaCSR[ 185 ][ 28 ],
   alphaCSR[ 185 ][ 29 ],
   alphaCSR[ 185 ][ 30 ],
   alphaCSR[ 185 ][ 31 ],
   alphaCSR[ 185 ][ 32 ],
   alphaCSR[ 185 ][ 33 ],
   alphaCSR[ 185 ][ 34 ],
   alphaCSR[ 185 ][ 35 ],
   alphaCSR[ 185 ][ 36 ],
   alphaCSR[ 185 ][ 37 ],
   alphaCSR[ 185 ][ 38 ],
   alphaCSR[ 185 ][ 39 ],
   alphaCSR[ 185 ][ 40 ],
   alphaCSR[ 185 ][ 41 ],
   alphaCSR[ 185 ][ 42 ],
   alphaCSR[ 185 ][ 43 ],
   alphaCSR[ 185 ][ 44 ],
   alphaCSR[ 185 ][ 45 ],
   alphaCSR[ 185 ][ 46 ],
   alphaCSR[ 185 ][ 47 ],
   alphaCSR[ 185 ][ 48 ],
   alphaCSR[ 185 ][ 49 ],
   alphaCSR[ 185 ][ 50 ],
   alphaCSR[ 185 ][ 51 ],
   alphaCSR[ 185 ][ 52 ],
   alphaCSR[ 185 ][ 53 ],
   alphaCSR[ 185 ][ 54 ],
   alphaCSR[ 185 ][ 55 ],
   alphaCSR[ 185 ][ 56 ],
   alphaCSR[ 185 ][ 57 ],
   alphaCSR[ 185 ][ 58 ],
   alphaCSR[ 185 ][ 59 ],
   alphaCSR[ 185 ][ 60 ],
   alphaCSR[ 185 ][ 61 ],
   alphaCSR[ 185 ][ 62 ],
   alphaCSR[ 185 ][ 63 ],
   alphaCSR[ 185 ][ 64 ],
   alphaCSR[ 185 ][ 65 ],
   alphaCSR[ 185 ][ 66 ],
   alphaCSR[ 185 ][ 67 ],
   alphaCSR[ 185 ][ 68 ],
   alphaCSR[ 185 ][ 69 ],
   alphaCSR[ 185 ][ 70 ],
   alphaCSR[ 185 ][ 71 ],
   alphaCSR[ 185 ][ 72 ],
   alphaCSR[ 185 ][ 73 ],
   alphaCSR[ 185 ][ 74 ],
   alphaCSR[ 185 ][ 75 ],
   alphaCSR[ 185 ][ 76 ],
   alphaCSR[ 185 ][ 77 ],
   alphaCSR[ 185 ][ 78 ],
   alphaCSR[ 185 ][ 79 ],
   alphaCSR[ 185 ][ 80 ],
   alphaCSR[ 185 ][ 81 ],
   alphaCSR[ 185 ][ 82 ],
   alphaCSR[ 185 ][ 83 ],
   alphaCSR[ 185 ][ 84 ],
   alphaCSR[ 185 ][ 85 ],
   alphaCSR[ 185 ][ 86 ],
   alphaCSR[ 185 ][ 87 ],
   alphaCSR[ 185 ][ 88 ],
   alphaCSR[ 185 ][ 89 ],
   alphaCSR[ 185 ][ 90 ],
   alphaCSR[ 185 ][ 91 ],
   alphaCSR[ 185 ][ 92 ],
   alphaCSR[ 185 ][ 93 ],
   alphaCSR[ 185 ][ 94 ],
   alphaCSR[ 185 ][ 95 ],
   alphaCSR[ 185 ][ 96 ],
   alphaCSR[ 185 ][ 97 ],
   alphaCSR[ 185 ][ 98 ],
   alphaCSR[ 185 ][ 99 ],
   alphaCSR[ 185 ][ 100 ],
   alphaCSR[ 185 ][ 101 ],
   alphaCSR[ 185 ][ 102 ],
   alphaCSR[ 185 ][ 103 ],
   alphaCSR[ 185 ][ 104 ],
   alphaCSR[ 185 ][ 105 ],
   alphaCSR[ 185 ][ 106 ],
   alphaCSR[ 185 ][ 107 ],
   alphaCSR[ 185 ][ 108 ],
   alphaCSR[ 185 ][ 109 ],
   alphaCSR[ 185 ][ 110 ],
   alphaCSR[ 185 ][ 111 ],
   alphaCSR[ 185 ][ 112 ],
   alphaCSR[ 185 ][ 113 ],
   alphaCSR[ 185 ][ 114 ],
   alphaCSR[ 185 ][ 115 ],
   alphaCSR[ 185 ][ 116 ],
   alphaCSR[ 185 ][ 117 ],
   alphaCSR[ 185 ][ 118 ],
   alphaCSR[ 185 ][ 119 ],
   alphaCSR[ 185 ][ 120 ],
   alphaCSR[ 185 ][ 121 ],
   alphaCSR[ 185 ][ 122 ],
   alphaCSR[ 185 ][ 123 ],
   alphaCSR[ 185 ][ 124 ],
   alphaCSR[ 185 ][ 125 ],
   alphaCSR[ 185 ][ 126 ],
   alphaCSR[ 185 ][ 127 ],
   alphaCSR[ 185 ][ 128 ],
   alphaCSR[ 185 ][ 129 ],
   alphaCSR[ 185 ][ 130 ],
   alphaCSR[ 185 ][ 131 ],
   alphaCSR[ 185 ][ 132 ],
   alphaCSR[ 185 ][ 133 ],
   alphaCSR[ 185 ][ 134 ],
   alphaCSR[ 185 ][ 135 ],
   alphaCSR[ 185 ][ 136 ],
   alphaCSR[ 185 ][ 137 ],
   alphaCSR[ 185 ][ 138 ],
   alphaCSR[ 185 ][ 139 ],
   alphaCSR[ 185 ][ 140 ],
   alphaCSR[ 185 ][ 141 ],
   alphaCSR[ 185 ][ 142 ],
   alphaCSR[ 185 ][ 143 ],
   alphaCSR[ 185 ][ 144 ],
   alphaCSR[ 185 ][ 145 ],
   alphaCSR[ 185 ][ 146 ],
   alphaCSR[ 185 ][ 147 ],
   alphaCSR[ 185 ][ 148 ],
   alphaCSR[ 185 ][ 149 ],
   alphaCSR[ 185 ][ 150 ],
   alphaCSR[ 185 ][ 151 ],
   alphaCSR[ 185 ][ 152 ],
   alphaCSR[ 185 ][ 153 ],
   alphaCSR[ 185 ][ 154 ],
   alphaCSR[ 185 ][ 155 ],
   alphaCSR[ 185 ][ 156 ],
   alphaCSR[ 185 ][ 157 ],
   alphaCSR[ 185 ][ 158 ],
   alphaCSR[ 185 ][ 159 ],
   alphaCSR[ 185 ][ 160 ],
   alphaCSR[ 185 ][ 161 ],
   alphaCSR[ 185 ][ 162 ],
   alphaCSR[ 185 ][ 163 ],
   alphaCSR[ 185 ][ 164 ],
   alphaCSR[ 185 ][ 165 ],
   alphaCSR[ 185 ][ 166 ],
   alphaCSR[ 185 ][ 167 ],
   alphaCSR[ 185 ][ 168 ],
   alphaCSR[ 185 ][ 169 ],
   alphaCSR[ 185 ][ 170 ],
   alphaCSR[ 185 ][ 171 ],
   alphaCSR[ 185 ][ 172 ],
   alphaCSR[ 185 ][ 173 ],
   alphaCSR[ 185 ][ 174 ],
   alphaCSR[ 185 ][ 175 ],
   alphaCSR[ 185 ][ 176 ],
   alphaCSR[ 185 ][ 177 ],
   alphaCSR[ 185 ][ 178 ],
   alphaCSR[ 185 ][ 179 ],
   alphaCSR[ 185 ][ 180 ],
   alphaCSR[ 185 ][ 181 ],
   alphaCSR[ 185 ][ 182 ],
   alphaCSR[ 185 ][ 183 ],
   alphaCSR[ 185 ][ 184 ],
   alphaCSR[ 185 ][ 185 ],
   alphaCSR[ 185 ][ 186 ],
   alphaCSR[ 185 ][ 187 ],
   alphaCSR[ 185 ][ 188 ],
   alphaCSR[ 185 ][ 189 ],
   alphaCSR[ 185 ][ 190 ],
   alphaCSR[ 185 ][ 191 ],
   alphaCSR[ 185 ][ 192 ],
   alphaCSR[ 185 ][ 193 ],
   alphaCSR[ 185 ][ 194 ],
   alphaCSR[ 185 ][ 195 ],
   alphaCSR[ 185 ][ 196 ],
   alphaCSR[ 185 ][ 197 ],
   alphaCSR[ 185 ][ 198 ],
   alphaCSR[ 185 ][ 199 ],
   alphaCSR[ 185 ][ 200 ],
   alphaCSR[ 185 ][ 201 ],
   alphaCSR[ 185 ][ 202 ],
   alphaCSR[ 185 ][ 203 ],
   alphaCSR[ 185 ][ 204 ],
   alphaCSR[ 185 ][ 205 ],
   alphaCSR[ 185 ][ 206 ],
   alphaCSR[ 185 ][ 207 ],
   alphaCSR[ 185 ][ 208 ],
   alphaCSR[ 185 ][ 209 ],
   alphaCSR[ 185 ][ 210 ],
   alphaCSR[ 185 ][ 211 ],
   alphaCSR[ 185 ][ 212 ],
   alphaCSR[ 185 ][ 213 ],
   alphaCSR[ 185 ][ 214 ],
   alphaCSR[ 185 ][ 215 ],
   alphaCSR[ 185 ][ 216 ],
   alphaCSR[ 185 ][ 217 ],
   alphaCSR[ 185 ][ 218 ],
   alphaCSR[ 185 ][ 219 ],
   alphaCSR[ 185 ][ 220 ],
   alphaCSR[ 185 ][ 221 ],
   alphaCSR[ 185 ][ 222 ],
   alphaCSR[ 185 ][ 223 ],
   alphaCSR[ 185 ][ 224 ],
   alphaCSR[ 185 ][ 225 ],
   alphaCSR[ 185 ][ 226 ],
   alphaCSR[ 185 ][ 227 ],
   alphaCSR[ 185 ][ 228 ],
   alphaCSR[ 185 ][ 229 ],
   alphaCSR[ 185 ][ 230 ],
   alphaCSR[ 185 ][ 231 ],
   alphaCSR[ 185 ][ 232 ],
   alphaCSR[ 185 ][ 233 ],
   alphaCSR[ 185 ][ 234 ],
   alphaCSR[ 185 ][ 235 ],
   alphaCSR[ 185 ][ 236 ],
   alphaCSR[ 185 ][ 237 ],
   alphaCSR[ 185 ][ 238 ],
   alphaCSR[ 185 ][ 239 ],
   alphaCSR[ 185 ][ 240 ],
   alphaCSR[ 185 ][ 241 ],
   alphaCSR[ 185 ][ 242 ],
   alphaCSR[ 185 ][ 243 ],
   alphaCSR[ 185 ][ 244 ],
   alphaCSR[ 185 ][ 245 ],
   alphaCSR[ 185 ][ 246 ],
   alphaCSR[ 185 ][ 247 ],
   alphaCSR[ 185 ][ 248 ],
   alphaCSR[ 185 ][ 249 ],
   alphaCSR[ 185 ][ 250 ],
   alphaCSR[ 185 ][ 251 ],
   alphaCSR[ 185 ][ 252 ],
   alphaCSR[ 185 ][ 253 ],
   alphaCSR[ 185 ][ 254 ],
   alphaCSR[ 185 ][ 255 ],
   alphaCSR[ 185 ][ 256 ],
   alphaCSR[ 185 ][ 257 ],
   alphaCSR[ 185 ][ 258 ],
   alphaCSR[ 185 ][ 259 ],
   alphaCSR[ 185 ][ 260 ],
   alphaCSR[ 185 ][ 261 ],
   alphaCSR[ 185 ][ 262 ],
   alphaCSR[ 185 ][ 263 ],
   alphaCSR[ 185 ][ 264 ],
   alphaCSR[ 185 ][ 265 ],
   alphaCSR[ 185 ][ 266 ],
   alphaCSR[ 185 ][ 267 ],
   alphaCSR[ 185 ][ 268 ],
   alphaCSR[ 185 ][ 269 ],
   alphaCSR[ 185 ][ 270 ],
   alphaCSR[ 185 ][ 271 ],
   alphaCSR[ 185 ][ 272 ],
   alphaCSR[ 185 ][ 273 ],
   alphaCSR[ 185 ][ 274 ],
   alphaCSR[ 185 ][ 275 ],
   alphaCSR[ 185 ][ 276 ],
   alphaCSR[ 185 ][ 277 ],
   alphaCSR[ 185 ][ 278 ],
   alphaCSR[ 185 ][ 279 ],
   alphaCSR[ 185 ][ 280 ],
   alphaCSR[ 185 ][ 281 ],
   alphaCSR[ 185 ][ 282 ],
   alphaCSR[ 185 ][ 283 ],
   alphaCSR[ 185 ][ 284 ],
   alphaCSR[ 185 ][ 285 ],
   alphaCSR[ 185 ][ 286 ],
   alphaCSR[ 185 ][ 287 ],
   alphaCSR[ 185 ][ 288 ],
   alphaCSR[ 185 ][ 289 ],
   alphaCSR[ 185 ][ 290 ],
   alphaCSR[ 185 ][ 291 ],
   alphaCSR[ 185 ][ 292 ],
   alphaCSR[ 185 ][ 293 ],
   alphaCSR[ 185 ][ 294 ],
   alphaCSR[ 185 ][ 295 ],
   alphaCSR[ 185 ][ 296 ],
   alphaCSR[ 185 ][ 297 ],
   alphaCSR[ 185 ][ 298 ],
   alphaCSR[ 185 ][ 299 ],
   alphaCSR[ 185 ][ 300 ],
   alphaCSR[ 185 ][ 301 ],
   alphaCSR[ 185 ][ 302 ],
   alphaCSR[ 185 ][ 303 ],
   alphaCSR[ 185 ][ 304 ],
   alphaCSR[ 185 ][ 305 ],
   alphaCSR[ 185 ][ 306 ],
   alphaCSR[ 185 ][ 307 ],
   alphaCSR[ 185 ][ 308 ],
   alphaCSR[ 185 ][ 309 ],
   alphaCSR[ 185 ][ 310 ],
   alphaCSR[ 185 ][ 311 ],
   alphaCSR[ 185 ][ 312 ],
   alphaCSR[ 185 ][ 313 ],
   alphaCSR[ 185 ][ 314 ],
   alphaCSR[ 185 ][ 315 ],
   alphaCSR[ 185 ][ 316 ],
   alphaCSR[ 185 ][ 317 ],
   alphaCSR[ 185 ][ 318 ],
   alphaCSR[ 185 ][ 319 ],
   alphaCSR[ 185 ][ 320 ],
   alphaCSR[ 185 ][ 321 ],
   alphaCSR[ 185 ][ 322 ],
   alphaCSR[ 185 ][ 323 ],
   alphaCSR[ 185 ][ 324 ],
   alphaCSR[ 185 ][ 325 ],
   alphaCSR[ 185 ][ 326 ],
   alphaCSR[ 185 ][ 327 ],
   alphaCSR[ 185 ][ 328 ],
   alphaCSR[ 185 ][ 329 ],
   alphaCSR[ 185 ][ 330 ],
   alphaCSR[ 185 ][ 331 ],
   alphaCSR[ 185 ][ 332 ],
   alphaCSR[ 185 ][ 333 ],
   alphaCSR[ 185 ][ 334 ],
   alphaCSR[ 185 ][ 335 ],
   alphaCSR[ 185 ][ 336 ],
   alphaCSR[ 185 ][ 337 ],
   alphaCSR[ 185 ][ 338 ],
   alphaCSR[ 185 ][ 339 ],
   alphaCSR[ 185 ][ 340 ],
   alphaCSR[ 185 ][ 341 ],
   alphaCSR[ 185 ][ 342 ],
   alphaCSR[ 185 ][ 343 ],
   alphaCSR[ 185 ][ 344 ],
   alphaCSR[ 185 ][ 345 ],
   alphaCSR[ 185 ][ 346 ],
   alphaCSR[ 185 ][ 347 ],
   alphaCSR[ 185 ][ 348 ],
   alphaCSR[ 185 ][ 349 ],
   alphaCSR[ 185 ][ 350 ],
   alphaCSR[ 185 ][ 351 ],
   alphaCSR[ 185 ][ 352 ],
   alphaCSR[ 185 ][ 353 ],
   alphaCSR[ 185 ][ 354 ],
   alphaCSR[ 185 ][ 355 ],
   alphaCSR[ 185 ][ 356 ],
   alphaCSR[ 185 ][ 357 ],
   alphaCSR[ 185 ][ 358 ],
   alphaCSR[ 185 ][ 359 ],
   alphaCSR[ 185 ][ 360 ],
   alphaCSR[ 185 ][ 361 ],
   alphaCSR[ 185 ][ 362 ],
   alphaCSR[ 185 ][ 363 ],
   alphaCSR[ 185 ][ 364 ],
   alphaCSR[ 185 ][ 365 ],
   alphaCSR[ 185 ][ 366 ],
   alphaCSR[ 185 ][ 367 ],
   alphaCSR[ 185 ][ 368 ],
   alphaCSR[ 185 ][ 369 ],
   alphaCSR[ 185 ][ 370 ],
   alphaCSR[ 185 ][ 371 ],
   alphaCSR[ 185 ][ 372 ],
   alphaCSR[ 185 ][ 373 ],
   alphaCSR[ 185 ][ 374 ],
   alphaCSR[ 185 ][ 375 ],
   alphaCSR[ 185 ][ 376 ],
   alphaCSR[ 185 ][ 377 ],
   alphaCSR[ 185 ][ 378 ],
   alphaCSR[ 185 ][ 379 ],
   alphaCSR[ 185 ][ 380 ],
   alphaCSR[ 185 ][ 381 ],
   alphaCSR[ 185 ][ 382 ],
   alphaCSR[ 185 ][ 383 ],
   alphaCSR[ 186 ][ 0 ],
   alphaCSR[ 186 ][ 1 ],
   alphaCSR[ 186 ][ 2 ],
   alphaCSR[ 186 ][ 3 ],
   alphaCSR[ 186 ][ 4 ],
   alphaCSR[ 186 ][ 5 ],
   alphaCSR[ 186 ][ 6 ],
   alphaCSR[ 186 ][ 7 ],
   alphaCSR[ 186 ][ 8 ],
   alphaCSR[ 186 ][ 9 ],
   alphaCSR[ 186 ][ 10 ],
   alphaCSR[ 186 ][ 11 ],
   alphaCSR[ 186 ][ 12 ],
   alphaCSR[ 186 ][ 13 ],
   alphaCSR[ 186 ][ 14 ],
   alphaCSR[ 186 ][ 15 ],
   alphaCSR[ 186 ][ 16 ],
   alphaCSR[ 186 ][ 17 ],
   alphaCSR[ 186 ][ 18 ],
   alphaCSR[ 186 ][ 19 ],
   alphaCSR[ 186 ][ 20 ],
   alphaCSR[ 186 ][ 21 ],
   alphaCSR[ 186 ][ 22 ],
   alphaCSR[ 186 ][ 23 ],
   alphaCSR[ 186 ][ 24 ],
   alphaCSR[ 186 ][ 25 ],
   alphaCSR[ 186 ][ 26 ],
   alphaCSR[ 186 ][ 27 ],
   alphaCSR[ 186 ][ 28 ],
   alphaCSR[ 186 ][ 29 ],
   alphaCSR[ 186 ][ 30 ],
   alphaCSR[ 186 ][ 31 ],
   alphaCSR[ 186 ][ 32 ],
   alphaCSR[ 186 ][ 33 ],
   alphaCSR[ 186 ][ 34 ],
   alphaCSR[ 186 ][ 35 ],
   alphaCSR[ 186 ][ 36 ],
   alphaCSR[ 186 ][ 37 ],
   alphaCSR[ 186 ][ 38 ],
   alphaCSR[ 186 ][ 39 ],
   alphaCSR[ 186 ][ 40 ],
   alphaCSR[ 186 ][ 41 ],
   alphaCSR[ 186 ][ 42 ],
   alphaCSR[ 186 ][ 43 ],
   alphaCSR[ 186 ][ 44 ],
   alphaCSR[ 186 ][ 45 ],
   alphaCSR[ 186 ][ 46 ],
   alphaCSR[ 186 ][ 47 ],
   alphaCSR[ 186 ][ 48 ],
   alphaCSR[ 186 ][ 49 ],
   alphaCSR[ 186 ][ 50 ],
   alphaCSR[ 186 ][ 51 ],
   alphaCSR[ 186 ][ 52 ],
   alphaCSR[ 186 ][ 53 ],
   alphaCSR[ 186 ][ 54 ],
   alphaCSR[ 186 ][ 55 ],
   alphaCSR[ 186 ][ 56 ],
   alphaCSR[ 186 ][ 57 ],
   alphaCSR[ 186 ][ 58 ],
   alphaCSR[ 186 ][ 59 ],
   alphaCSR[ 186 ][ 60 ],
   alphaCSR[ 186 ][ 61 ],
   alphaCSR[ 186 ][ 62 ],
   alphaCSR[ 186 ][ 63 ],
   alphaCSR[ 186 ][ 64 ],
   alphaCSR[ 186 ][ 65 ],
   alphaCSR[ 186 ][ 66 ],
   alphaCSR[ 186 ][ 67 ],
   alphaCSR[ 186 ][ 68 ],
   alphaCSR[ 186 ][ 69 ],
   alphaCSR[ 186 ][ 70 ],
   alphaCSR[ 186 ][ 71 ],
   alphaCSR[ 186 ][ 72 ],
   alphaCSR[ 186 ][ 73 ],
   alphaCSR[ 186 ][ 74 ],
   alphaCSR[ 186 ][ 75 ],
   alphaCSR[ 186 ][ 76 ],
   alphaCSR[ 186 ][ 77 ],
   alphaCSR[ 186 ][ 78 ],
   alphaCSR[ 186 ][ 79 ],
   alphaCSR[ 186 ][ 80 ],
   alphaCSR[ 186 ][ 81 ],
   alphaCSR[ 186 ][ 82 ],
   alphaCSR[ 186 ][ 83 ],
   alphaCSR[ 186 ][ 84 ],
   alphaCSR[ 186 ][ 85 ],
   alphaCSR[ 186 ][ 86 ],
   alphaCSR[ 186 ][ 87 ],
   alphaCSR[ 186 ][ 88 ],
   alphaCSR[ 186 ][ 89 ],
   alphaCSR[ 186 ][ 90 ],
   alphaCSR[ 186 ][ 91 ],
   alphaCSR[ 186 ][ 92 ],
   alphaCSR[ 186 ][ 93 ],
   alphaCSR[ 186 ][ 94 ],
   alphaCSR[ 186 ][ 95 ],
   alphaCSR[ 186 ][ 96 ],
   alphaCSR[ 186 ][ 97 ],
   alphaCSR[ 186 ][ 98 ],
   alphaCSR[ 186 ][ 99 ],
   alphaCSR[ 186 ][ 100 ],
   alphaCSR[ 186 ][ 101 ],
   alphaCSR[ 186 ][ 102 ],
   alphaCSR[ 186 ][ 103 ],
   alphaCSR[ 186 ][ 104 ],
   alphaCSR[ 186 ][ 105 ],
   alphaCSR[ 186 ][ 106 ],
   alphaCSR[ 186 ][ 107 ],
   alphaCSR[ 186 ][ 108 ],
   alphaCSR[ 186 ][ 109 ],
   alphaCSR[ 186 ][ 110 ],
   alphaCSR[ 186 ][ 111 ],
   alphaCSR[ 186 ][ 112 ],
   alphaCSR[ 186 ][ 113 ],
   alphaCSR[ 186 ][ 114 ],
   alphaCSR[ 186 ][ 115 ],
   alphaCSR[ 186 ][ 116 ],
   alphaCSR[ 186 ][ 117 ],
   alphaCSR[ 186 ][ 118 ],
   alphaCSR[ 186 ][ 119 ],
   alphaCSR[ 186 ][ 120 ],
   alphaCSR[ 186 ][ 121 ],
   alphaCSR[ 186 ][ 122 ],
   alphaCSR[ 186 ][ 123 ],
   alphaCSR[ 186 ][ 124 ],
   alphaCSR[ 186 ][ 125 ],
   alphaCSR[ 186 ][ 126 ],
   alphaCSR[ 186 ][ 127 ],
   alphaCSR[ 186 ][ 128 ],
   alphaCSR[ 186 ][ 129 ],
   alphaCSR[ 186 ][ 130 ],
   alphaCSR[ 186 ][ 131 ],
   alphaCSR[ 186 ][ 132 ],
   alphaCSR[ 186 ][ 133 ],
   alphaCSR[ 186 ][ 134 ],
   alphaCSR[ 186 ][ 135 ],
   alphaCSR[ 186 ][ 136 ],
   alphaCSR[ 186 ][ 137 ],
   alphaCSR[ 186 ][ 138 ],
   alphaCSR[ 186 ][ 139 ],
   alphaCSR[ 186 ][ 140 ],
   alphaCSR[ 186 ][ 141 ],
   alphaCSR[ 186 ][ 142 ],
   alphaCSR[ 186 ][ 143 ],
   alphaCSR[ 186 ][ 144 ],
   alphaCSR[ 186 ][ 145 ],
   alphaCSR[ 186 ][ 146 ],
   alphaCSR[ 186 ][ 147 ],
   alphaCSR[ 186 ][ 148 ],
   alphaCSR[ 186 ][ 149 ],
   alphaCSR[ 186 ][ 150 ],
   alphaCSR[ 186 ][ 151 ],
   alphaCSR[ 186 ][ 152 ],
   alphaCSR[ 186 ][ 153 ],
   alphaCSR[ 186 ][ 154 ],
   alphaCSR[ 186 ][ 155 ],
   alphaCSR[ 186 ][ 156 ],
   alphaCSR[ 186 ][ 157 ],
   alphaCSR[ 186 ][ 158 ],
   alphaCSR[ 186 ][ 159 ],
   alphaCSR[ 186 ][ 160 ],
   alphaCSR[ 186 ][ 161 ],
   alphaCSR[ 186 ][ 162 ],
   alphaCSR[ 186 ][ 163 ],
   alphaCSR[ 186 ][ 164 ],
   alphaCSR[ 186 ][ 165 ],
   alphaCSR[ 186 ][ 166 ],
   alphaCSR[ 186 ][ 167 ],
   alphaCSR[ 186 ][ 168 ],
   alphaCSR[ 186 ][ 169 ],
   alphaCSR[ 186 ][ 170 ],
   alphaCSR[ 186 ][ 171 ],
   alphaCSR[ 186 ][ 172 ],
   alphaCSR[ 186 ][ 173 ],
   alphaCSR[ 186 ][ 174 ],
   alphaCSR[ 186 ][ 175 ],
   alphaCSR[ 186 ][ 176 ],
   alphaCSR[ 186 ][ 177 ],
   alphaCSR[ 186 ][ 178 ],
   alphaCSR[ 186 ][ 179 ],
   alphaCSR[ 186 ][ 180 ],
   alphaCSR[ 186 ][ 181 ],
   alphaCSR[ 186 ][ 182 ],
   alphaCSR[ 186 ][ 183 ],
   alphaCSR[ 186 ][ 184 ],
   alphaCSR[ 186 ][ 185 ],
   alphaCSR[ 186 ][ 186 ],
   alphaCSR[ 186 ][ 187 ],
   alphaCSR[ 186 ][ 188 ],
   alphaCSR[ 186 ][ 189 ],
   alphaCSR[ 186 ][ 190 ],
   alphaCSR[ 186 ][ 191 ],
   alphaCSR[ 186 ][ 192 ],
   alphaCSR[ 186 ][ 193 ],
   alphaCSR[ 186 ][ 194 ],
   alphaCSR[ 186 ][ 195 ],
   alphaCSR[ 186 ][ 196 ],
   alphaCSR[ 186 ][ 197 ],
   alphaCSR[ 186 ][ 198 ],
   alphaCSR[ 186 ][ 199 ],
   alphaCSR[ 186 ][ 200 ],
   alphaCSR[ 186 ][ 201 ],
   alphaCSR[ 186 ][ 202 ],
   alphaCSR[ 186 ][ 203 ],
   alphaCSR[ 186 ][ 204 ],
   alphaCSR[ 186 ][ 205 ],
   alphaCSR[ 186 ][ 206 ],
   alphaCSR[ 186 ][ 207 ],
   alphaCSR[ 186 ][ 208 ],
   alphaCSR[ 186 ][ 209 ],
   alphaCSR[ 186 ][ 210 ],
   alphaCSR[ 186 ][ 211 ],
   alphaCSR[ 186 ][ 212 ],
   alphaCSR[ 186 ][ 213 ],
   alphaCSR[ 186 ][ 214 ],
   alphaCSR[ 186 ][ 215 ],
   alphaCSR[ 186 ][ 216 ],
   alphaCSR[ 186 ][ 217 ],
   alphaCSR[ 186 ][ 218 ],
   alphaCSR[ 186 ][ 219 ],
   alphaCSR[ 186 ][ 220 ],
   alphaCSR[ 186 ][ 221 ],
   alphaCSR[ 186 ][ 222 ],
   alphaCSR[ 186 ][ 223 ],
   alphaCSR[ 186 ][ 224 ],
   alphaCSR[ 186 ][ 225 ],
   alphaCSR[ 186 ][ 226 ],
   alphaCSR[ 186 ][ 227 ],
   alphaCSR[ 186 ][ 228 ],
   alphaCSR[ 186 ][ 229 ],
   alphaCSR[ 186 ][ 230 ],
   alphaCSR[ 186 ][ 231 ],
   alphaCSR[ 186 ][ 232 ],
   alphaCSR[ 186 ][ 233 ],
   alphaCSR[ 186 ][ 234 ],
   alphaCSR[ 186 ][ 235 ],
   alphaCSR[ 186 ][ 236 ],
   alphaCSR[ 186 ][ 237 ],
   alphaCSR[ 186 ][ 238 ],
   alphaCSR[ 186 ][ 239 ],
   alphaCSR[ 186 ][ 240 ],
   alphaCSR[ 186 ][ 241 ],
   alphaCSR[ 186 ][ 242 ],
   alphaCSR[ 186 ][ 243 ],
   alphaCSR[ 186 ][ 244 ],
   alphaCSR[ 186 ][ 245 ],
   alphaCSR[ 186 ][ 246 ],
   alphaCSR[ 186 ][ 247 ],
   alphaCSR[ 186 ][ 248 ],
   alphaCSR[ 186 ][ 249 ],
   alphaCSR[ 186 ][ 250 ],
   alphaCSR[ 186 ][ 251 ],
   alphaCSR[ 186 ][ 252 ],
   alphaCSR[ 186 ][ 253 ],
   alphaCSR[ 186 ][ 254 ],
   alphaCSR[ 186 ][ 255 ],
   alphaCSR[ 186 ][ 256 ],
   alphaCSR[ 186 ][ 257 ],
   alphaCSR[ 186 ][ 258 ],
   alphaCSR[ 186 ][ 259 ],
   alphaCSR[ 186 ][ 260 ],
   alphaCSR[ 186 ][ 261 ],
   alphaCSR[ 186 ][ 262 ],
   alphaCSR[ 186 ][ 263 ],
   alphaCSR[ 186 ][ 264 ],
   alphaCSR[ 186 ][ 265 ],
   alphaCSR[ 186 ][ 266 ],
   alphaCSR[ 186 ][ 267 ],
   alphaCSR[ 186 ][ 268 ],
   alphaCSR[ 186 ][ 269 ],
   alphaCSR[ 186 ][ 270 ],
   alphaCSR[ 186 ][ 271 ],
   alphaCSR[ 186 ][ 272 ],
   alphaCSR[ 186 ][ 273 ],
   alphaCSR[ 186 ][ 274 ],
   alphaCSR[ 186 ][ 275 ],
   alphaCSR[ 186 ][ 276 ],
   alphaCSR[ 186 ][ 277 ],
   alphaCSR[ 186 ][ 278 ],
   alphaCSR[ 186 ][ 279 ],
   alphaCSR[ 186 ][ 280 ],
   alphaCSR[ 186 ][ 281 ],
   alphaCSR[ 186 ][ 282 ],
   alphaCSR[ 186 ][ 283 ],
   alphaCSR[ 186 ][ 284 ],
   alphaCSR[ 186 ][ 285 ],
   alphaCSR[ 186 ][ 286 ],
   alphaCSR[ 186 ][ 287 ],
   alphaCSR[ 186 ][ 288 ],
   alphaCSR[ 186 ][ 289 ],
   alphaCSR[ 186 ][ 290 ],
   alphaCSR[ 186 ][ 291 ],
   alphaCSR[ 186 ][ 292 ],
   alphaCSR[ 186 ][ 293 ],
   alphaCSR[ 186 ][ 294 ],
   alphaCSR[ 186 ][ 295 ],
   alphaCSR[ 186 ][ 296 ],
   alphaCSR[ 186 ][ 297 ],
   alphaCSR[ 186 ][ 298 ],
   alphaCSR[ 186 ][ 299 ],
   alphaCSR[ 186 ][ 300 ],
   alphaCSR[ 186 ][ 301 ],
   alphaCSR[ 186 ][ 302 ],
   alphaCSR[ 186 ][ 303 ],
   alphaCSR[ 186 ][ 304 ],
   alphaCSR[ 186 ][ 305 ],
   alphaCSR[ 186 ][ 306 ],
   alphaCSR[ 186 ][ 307 ],
   alphaCSR[ 186 ][ 308 ],
   alphaCSR[ 186 ][ 309 ],
   alphaCSR[ 186 ][ 310 ],
   alphaCSR[ 186 ][ 311 ],
   alphaCSR[ 186 ][ 312 ],
   alphaCSR[ 186 ][ 313 ],
   alphaCSR[ 186 ][ 314 ],
   alphaCSR[ 186 ][ 315 ],
   alphaCSR[ 186 ][ 316 ],
   alphaCSR[ 186 ][ 317 ],
   alphaCSR[ 186 ][ 318 ],
   alphaCSR[ 186 ][ 319 ],
   alphaCSR[ 186 ][ 320 ],
   alphaCSR[ 186 ][ 321 ],
   alphaCSR[ 186 ][ 322 ],
   alphaCSR[ 186 ][ 323 ],
   alphaCSR[ 186 ][ 324 ],
   alphaCSR[ 186 ][ 325 ],
   alphaCSR[ 186 ][ 326 ],
   alphaCSR[ 186 ][ 327 ],
   alphaCSR[ 186 ][ 328 ],
   alphaCSR[ 186 ][ 329 ],
   alphaCSR[ 186 ][ 330 ],
   alphaCSR[ 186 ][ 331 ],
   alphaCSR[ 186 ][ 332 ],
   alphaCSR[ 186 ][ 333 ],
   alphaCSR[ 186 ][ 334 ],
   alphaCSR[ 186 ][ 335 ],
   alphaCSR[ 186 ][ 336 ],
   alphaCSR[ 186 ][ 337 ],
   alphaCSR[ 186 ][ 338 ],
   alphaCSR[ 186 ][ 339 ],
   alphaCSR[ 186 ][ 340 ],
   alphaCSR[ 186 ][ 341 ],
   alphaCSR[ 186 ][ 342 ],
   alphaCSR[ 186 ][ 343 ],
   alphaCSR[ 186 ][ 344 ],
   alphaCSR[ 186 ][ 345 ],
   alphaCSR[ 186 ][ 346 ],
   alphaCSR[ 186 ][ 347 ],
   alphaCSR[ 186 ][ 348 ],
   alphaCSR[ 186 ][ 349 ],
   alphaCSR[ 186 ][ 350 ],
   alphaCSR[ 186 ][ 351 ],
   alphaCSR[ 186 ][ 352 ],
   alphaCSR[ 186 ][ 353 ],
   alphaCSR[ 186 ][ 354 ],
   alphaCSR[ 186 ][ 355 ],
   alphaCSR[ 186 ][ 356 ],
   alphaCSR[ 186 ][ 357 ],
   alphaCSR[ 186 ][ 358 ],
   alphaCSR[ 186 ][ 359 ],
   alphaCSR[ 186 ][ 360 ],
   alphaCSR[ 186 ][ 361 ],
   alphaCSR[ 186 ][ 362 ],
   alphaCSR[ 186 ][ 363 ],
   alphaCSR[ 186 ][ 364 ],
   alphaCSR[ 186 ][ 365 ],
   alphaCSR[ 186 ][ 366 ],
   alphaCSR[ 186 ][ 367 ],
   alphaCSR[ 186 ][ 368 ],
   alphaCSR[ 186 ][ 369 ],
   alphaCSR[ 186 ][ 370 ],
   alphaCSR[ 186 ][ 371 ],
   alphaCSR[ 186 ][ 372 ],
   alphaCSR[ 186 ][ 373 ],
   alphaCSR[ 186 ][ 374 ],
   alphaCSR[ 186 ][ 375 ],
   alphaCSR[ 186 ][ 376 ],
   alphaCSR[ 186 ][ 377 ],
   alphaCSR[ 186 ][ 378 ],
   alphaCSR[ 186 ][ 379 ],
   alphaCSR[ 186 ][ 380 ],
   alphaCSR[ 186 ][ 381 ],
   alphaCSR[ 186 ][ 382 ],
   alphaCSR[ 186 ][ 383 ],
   alphaCSR[ 187 ][ 0 ],
   alphaCSR[ 187 ][ 1 ],
   alphaCSR[ 187 ][ 2 ],
   alphaCSR[ 187 ][ 3 ],
   alphaCSR[ 187 ][ 4 ],
   alphaCSR[ 187 ][ 5 ],
   alphaCSR[ 187 ][ 6 ],
   alphaCSR[ 187 ][ 7 ],
   alphaCSR[ 187 ][ 8 ],
   alphaCSR[ 187 ][ 9 ],
   alphaCSR[ 187 ][ 10 ],
   alphaCSR[ 187 ][ 11 ],
   alphaCSR[ 187 ][ 12 ],
   alphaCSR[ 187 ][ 13 ],
   alphaCSR[ 187 ][ 14 ],
   alphaCSR[ 187 ][ 15 ],
   alphaCSR[ 187 ][ 16 ],
   alphaCSR[ 187 ][ 17 ],
   alphaCSR[ 187 ][ 18 ],
   alphaCSR[ 187 ][ 19 ],
   alphaCSR[ 187 ][ 20 ],
   alphaCSR[ 187 ][ 21 ],
   alphaCSR[ 187 ][ 22 ],
   alphaCSR[ 187 ][ 23 ],
   alphaCSR[ 187 ][ 24 ],
   alphaCSR[ 187 ][ 25 ],
   alphaCSR[ 187 ][ 26 ],
   alphaCSR[ 187 ][ 27 ],
   alphaCSR[ 187 ][ 28 ],
   alphaCSR[ 187 ][ 29 ],
   alphaCSR[ 187 ][ 30 ],
   alphaCSR[ 187 ][ 31 ],
   alphaCSR[ 187 ][ 32 ],
   alphaCSR[ 187 ][ 33 ],
   alphaCSR[ 187 ][ 34 ],
   alphaCSR[ 187 ][ 35 ],
   alphaCSR[ 187 ][ 36 ],
   alphaCSR[ 187 ][ 37 ],
   alphaCSR[ 187 ][ 38 ],
   alphaCSR[ 187 ][ 39 ],
   alphaCSR[ 187 ][ 40 ],
   alphaCSR[ 187 ][ 41 ],
   alphaCSR[ 187 ][ 42 ],
   alphaCSR[ 187 ][ 43 ],
   alphaCSR[ 187 ][ 44 ],
   alphaCSR[ 187 ][ 45 ],
   alphaCSR[ 187 ][ 46 ],
   alphaCSR[ 187 ][ 47 ],
   alphaCSR[ 187 ][ 48 ],
   alphaCSR[ 187 ][ 49 ],
   alphaCSR[ 187 ][ 50 ],
   alphaCSR[ 187 ][ 51 ],
   alphaCSR[ 187 ][ 52 ],
   alphaCSR[ 187 ][ 53 ],
   alphaCSR[ 187 ][ 54 ],
   alphaCSR[ 187 ][ 55 ],
   alphaCSR[ 187 ][ 56 ],
   alphaCSR[ 187 ][ 57 ],
   alphaCSR[ 187 ][ 58 ],
   alphaCSR[ 187 ][ 59 ],
   alphaCSR[ 187 ][ 60 ],
   alphaCSR[ 187 ][ 61 ],
   alphaCSR[ 187 ][ 62 ],
   alphaCSR[ 187 ][ 63 ],
   alphaCSR[ 187 ][ 64 ],
   alphaCSR[ 187 ][ 65 ],
   alphaCSR[ 187 ][ 66 ],
   alphaCSR[ 187 ][ 67 ],
   alphaCSR[ 187 ][ 68 ],
   alphaCSR[ 187 ][ 69 ],
   alphaCSR[ 187 ][ 70 ],
   alphaCSR[ 187 ][ 71 ],
   alphaCSR[ 187 ][ 72 ],
   alphaCSR[ 187 ][ 73 ],
   alphaCSR[ 187 ][ 74 ],
   alphaCSR[ 187 ][ 75 ],
   alphaCSR[ 187 ][ 76 ],
   alphaCSR[ 187 ][ 77 ],
   alphaCSR[ 187 ][ 78 ],
   alphaCSR[ 187 ][ 79 ],
   alphaCSR[ 187 ][ 80 ],
   alphaCSR[ 187 ][ 81 ],
   alphaCSR[ 187 ][ 82 ],
   alphaCSR[ 187 ][ 83 ],
   alphaCSR[ 187 ][ 84 ],
   alphaCSR[ 187 ][ 85 ],
   alphaCSR[ 187 ][ 86 ],
   alphaCSR[ 187 ][ 87 ],
   alphaCSR[ 187 ][ 88 ],
   alphaCSR[ 187 ][ 89 ],
   alphaCSR[ 187 ][ 90 ],
   alphaCSR[ 187 ][ 91 ],
   alphaCSR[ 187 ][ 92 ],
   alphaCSR[ 187 ][ 93 ],
   alphaCSR[ 187 ][ 94 ],
   alphaCSR[ 187 ][ 95 ],
   alphaCSR[ 187 ][ 96 ],
   alphaCSR[ 187 ][ 97 ],
   alphaCSR[ 187 ][ 98 ],
   alphaCSR[ 187 ][ 99 ],
   alphaCSR[ 187 ][ 100 ],
   alphaCSR[ 187 ][ 101 ],
   alphaCSR[ 187 ][ 102 ],
   alphaCSR[ 187 ][ 103 ],
   alphaCSR[ 187 ][ 104 ],
   alphaCSR[ 187 ][ 105 ],
   alphaCSR[ 187 ][ 106 ],
   alphaCSR[ 187 ][ 107 ],
   alphaCSR[ 187 ][ 108 ],
   alphaCSR[ 187 ][ 109 ],
   alphaCSR[ 187 ][ 110 ],
   alphaCSR[ 187 ][ 111 ],
   alphaCSR[ 187 ][ 112 ],
   alphaCSR[ 187 ][ 113 ],
   alphaCSR[ 187 ][ 114 ],
   alphaCSR[ 187 ][ 115 ],
   alphaCSR[ 187 ][ 116 ],
   alphaCSR[ 187 ][ 117 ],
   alphaCSR[ 187 ][ 118 ],
   alphaCSR[ 187 ][ 119 ],
   alphaCSR[ 187 ][ 120 ],
   alphaCSR[ 187 ][ 121 ],
   alphaCSR[ 187 ][ 122 ],
   alphaCSR[ 187 ][ 123 ],
   alphaCSR[ 187 ][ 124 ],
   alphaCSR[ 187 ][ 125 ],
   alphaCSR[ 187 ][ 126 ],
   alphaCSR[ 187 ][ 127 ],
   alphaCSR[ 187 ][ 128 ],
   alphaCSR[ 187 ][ 129 ],
   alphaCSR[ 187 ][ 130 ],
   alphaCSR[ 187 ][ 131 ],
   alphaCSR[ 187 ][ 132 ],
   alphaCSR[ 187 ][ 133 ],
   alphaCSR[ 187 ][ 134 ],
   alphaCSR[ 187 ][ 135 ],
   alphaCSR[ 187 ][ 136 ],
   alphaCSR[ 187 ][ 137 ],
   alphaCSR[ 187 ][ 138 ],
   alphaCSR[ 187 ][ 139 ],
   alphaCSR[ 187 ][ 140 ],
   alphaCSR[ 187 ][ 141 ],
   alphaCSR[ 187 ][ 142 ],
   alphaCSR[ 187 ][ 143 ],
   alphaCSR[ 187 ][ 144 ],
   alphaCSR[ 187 ][ 145 ],
   alphaCSR[ 187 ][ 146 ],
   alphaCSR[ 187 ][ 147 ],
   alphaCSR[ 187 ][ 148 ],
   alphaCSR[ 187 ][ 149 ],
   alphaCSR[ 187 ][ 150 ],
   alphaCSR[ 187 ][ 151 ],
   alphaCSR[ 187 ][ 152 ],
   alphaCSR[ 187 ][ 153 ],
   alphaCSR[ 187 ][ 154 ],
   alphaCSR[ 187 ][ 155 ],
   alphaCSR[ 187 ][ 156 ],
   alphaCSR[ 187 ][ 157 ],
   alphaCSR[ 187 ][ 158 ],
   alphaCSR[ 187 ][ 159 ],
   alphaCSR[ 187 ][ 160 ],
   alphaCSR[ 187 ][ 161 ],
   alphaCSR[ 187 ][ 162 ],
   alphaCSR[ 187 ][ 163 ],
   alphaCSR[ 187 ][ 164 ],
   alphaCSR[ 187 ][ 165 ],
   alphaCSR[ 187 ][ 166 ],
   alphaCSR[ 187 ][ 167 ],
   alphaCSR[ 187 ][ 168 ],
   alphaCSR[ 187 ][ 169 ],
   alphaCSR[ 187 ][ 170 ],
   alphaCSR[ 187 ][ 171 ],
   alphaCSR[ 187 ][ 172 ],
   alphaCSR[ 187 ][ 173 ],
   alphaCSR[ 187 ][ 174 ],
   alphaCSR[ 187 ][ 175 ],
   alphaCSR[ 187 ][ 176 ],
   alphaCSR[ 187 ][ 177 ],
   alphaCSR[ 187 ][ 178 ],
   alphaCSR[ 187 ][ 179 ],
   alphaCSR[ 187 ][ 180 ],
   alphaCSR[ 187 ][ 181 ],
   alphaCSR[ 187 ][ 182 ],
   alphaCSR[ 187 ][ 183 ],
   alphaCSR[ 187 ][ 184 ],
   alphaCSR[ 187 ][ 185 ],
   alphaCSR[ 187 ][ 186 ],
   alphaCSR[ 187 ][ 187 ],
   alphaCSR[ 187 ][ 188 ],
   alphaCSR[ 187 ][ 189 ],
   alphaCSR[ 187 ][ 190 ],
   alphaCSR[ 187 ][ 191 ],
   alphaCSR[ 187 ][ 192 ],
   alphaCSR[ 187 ][ 193 ],
   alphaCSR[ 187 ][ 194 ],
   alphaCSR[ 187 ][ 195 ],
   alphaCSR[ 187 ][ 196 ],
   alphaCSR[ 187 ][ 197 ],
   alphaCSR[ 187 ][ 198 ],
   alphaCSR[ 187 ][ 199 ],
   alphaCSR[ 187 ][ 200 ],
   alphaCSR[ 187 ][ 201 ],
   alphaCSR[ 187 ][ 202 ],
   alphaCSR[ 187 ][ 203 ],
   alphaCSR[ 187 ][ 204 ],
   alphaCSR[ 187 ][ 205 ],
   alphaCSR[ 187 ][ 206 ],
   alphaCSR[ 187 ][ 207 ],
   alphaCSR[ 187 ][ 208 ],
   alphaCSR[ 187 ][ 209 ],
   alphaCSR[ 187 ][ 210 ],
   alphaCSR[ 187 ][ 211 ],
   alphaCSR[ 187 ][ 212 ],
   alphaCSR[ 187 ][ 213 ],
   alphaCSR[ 187 ][ 214 ],
   alphaCSR[ 187 ][ 215 ],
   alphaCSR[ 187 ][ 216 ],
   alphaCSR[ 187 ][ 217 ],
   alphaCSR[ 187 ][ 218 ],
   alphaCSR[ 187 ][ 219 ],
   alphaCSR[ 187 ][ 220 ],
   alphaCSR[ 187 ][ 221 ],
   alphaCSR[ 187 ][ 222 ],
   alphaCSR[ 187 ][ 223 ],
   alphaCSR[ 187 ][ 224 ],
   alphaCSR[ 187 ][ 225 ],
   alphaCSR[ 187 ][ 226 ],
   alphaCSR[ 187 ][ 227 ],
   alphaCSR[ 187 ][ 228 ],
   alphaCSR[ 187 ][ 229 ],
   alphaCSR[ 187 ][ 230 ],
   alphaCSR[ 187 ][ 231 ],
   alphaCSR[ 187 ][ 232 ],
   alphaCSR[ 187 ][ 233 ],
   alphaCSR[ 187 ][ 234 ],
   alphaCSR[ 187 ][ 235 ],
   alphaCSR[ 187 ][ 236 ],
   alphaCSR[ 187 ][ 237 ],
   alphaCSR[ 187 ][ 238 ],
   alphaCSR[ 187 ][ 239 ],
   alphaCSR[ 187 ][ 240 ],
   alphaCSR[ 187 ][ 241 ],
   alphaCSR[ 187 ][ 242 ],
   alphaCSR[ 187 ][ 243 ],
   alphaCSR[ 187 ][ 244 ],
   alphaCSR[ 187 ][ 245 ],
   alphaCSR[ 187 ][ 246 ],
   alphaCSR[ 187 ][ 247 ],
   alphaCSR[ 187 ][ 248 ],
   alphaCSR[ 187 ][ 249 ],
   alphaCSR[ 187 ][ 250 ],
   alphaCSR[ 187 ][ 251 ],
   alphaCSR[ 187 ][ 252 ],
   alphaCSR[ 187 ][ 253 ],
   alphaCSR[ 187 ][ 254 ],
   alphaCSR[ 187 ][ 255 ],
   alphaCSR[ 187 ][ 256 ],
   alphaCSR[ 187 ][ 257 ],
   alphaCSR[ 187 ][ 258 ],
   alphaCSR[ 187 ][ 259 ],
   alphaCSR[ 187 ][ 260 ],
   alphaCSR[ 187 ][ 261 ],
   alphaCSR[ 187 ][ 262 ],
   alphaCSR[ 187 ][ 263 ],
   alphaCSR[ 187 ][ 264 ],
   alphaCSR[ 187 ][ 265 ],
   alphaCSR[ 187 ][ 266 ],
   alphaCSR[ 187 ][ 267 ],
   alphaCSR[ 187 ][ 268 ],
   alphaCSR[ 187 ][ 269 ],
   alphaCSR[ 187 ][ 270 ],
   alphaCSR[ 187 ][ 271 ],
   alphaCSR[ 187 ][ 272 ],
   alphaCSR[ 187 ][ 273 ],
   alphaCSR[ 187 ][ 274 ],
   alphaCSR[ 187 ][ 275 ],
   alphaCSR[ 187 ][ 276 ],
   alphaCSR[ 187 ][ 277 ],
   alphaCSR[ 187 ][ 278 ],
   alphaCSR[ 187 ][ 279 ],
   alphaCSR[ 187 ][ 280 ],
   alphaCSR[ 187 ][ 281 ],
   alphaCSR[ 187 ][ 282 ],
   alphaCSR[ 187 ][ 283 ],
   alphaCSR[ 187 ][ 284 ],
   alphaCSR[ 187 ][ 285 ],
   alphaCSR[ 187 ][ 286 ],
   alphaCSR[ 187 ][ 287 ],
   alphaCSR[ 187 ][ 288 ],
   alphaCSR[ 187 ][ 289 ],
   alphaCSR[ 187 ][ 290 ],
   alphaCSR[ 187 ][ 291 ],
   alphaCSR[ 187 ][ 292 ],
   alphaCSR[ 187 ][ 293 ],
   alphaCSR[ 187 ][ 294 ],
   alphaCSR[ 187 ][ 295 ],
   alphaCSR[ 187 ][ 296 ],
   alphaCSR[ 187 ][ 297 ],
   alphaCSR[ 187 ][ 298 ],
   alphaCSR[ 187 ][ 299 ],
   alphaCSR[ 187 ][ 300 ],
   alphaCSR[ 187 ][ 301 ],
   alphaCSR[ 187 ][ 302 ],
   alphaCSR[ 187 ][ 303 ],
   alphaCSR[ 187 ][ 304 ],
   alphaCSR[ 187 ][ 305 ],
   alphaCSR[ 187 ][ 306 ],
   alphaCSR[ 187 ][ 307 ],
   alphaCSR[ 187 ][ 308 ],
   alphaCSR[ 187 ][ 309 ],
   alphaCSR[ 187 ][ 310 ],
   alphaCSR[ 187 ][ 311 ],
   alphaCSR[ 187 ][ 312 ],
   alphaCSR[ 187 ][ 313 ],
   alphaCSR[ 187 ][ 314 ],
   alphaCSR[ 187 ][ 315 ],
   alphaCSR[ 187 ][ 316 ],
   alphaCSR[ 187 ][ 317 ],
   alphaCSR[ 187 ][ 318 ],
   alphaCSR[ 187 ][ 319 ],
   alphaCSR[ 187 ][ 320 ],
   alphaCSR[ 187 ][ 321 ],
   alphaCSR[ 187 ][ 322 ],
   alphaCSR[ 187 ][ 323 ],
   alphaCSR[ 187 ][ 324 ],
   alphaCSR[ 187 ][ 325 ],
   alphaCSR[ 187 ][ 326 ],
   alphaCSR[ 187 ][ 327 ],
   alphaCSR[ 187 ][ 328 ],
   alphaCSR[ 187 ][ 329 ],
   alphaCSR[ 187 ][ 330 ],
   alphaCSR[ 187 ][ 331 ],
   alphaCSR[ 187 ][ 332 ],
   alphaCSR[ 187 ][ 333 ],
   alphaCSR[ 187 ][ 334 ],
   alphaCSR[ 187 ][ 335 ],
   alphaCSR[ 187 ][ 336 ],
   alphaCSR[ 187 ][ 337 ],
   alphaCSR[ 187 ][ 338 ],
   alphaCSR[ 187 ][ 339 ],
   alphaCSR[ 187 ][ 340 ],
   alphaCSR[ 187 ][ 341 ],
   alphaCSR[ 187 ][ 342 ],
   alphaCSR[ 187 ][ 343 ],
   alphaCSR[ 187 ][ 344 ],
   alphaCSR[ 187 ][ 345 ],
   alphaCSR[ 187 ][ 346 ],
   alphaCSR[ 187 ][ 347 ],
   alphaCSR[ 187 ][ 348 ],
   alphaCSR[ 187 ][ 349 ],
   alphaCSR[ 187 ][ 350 ],
   alphaCSR[ 187 ][ 351 ],
   alphaCSR[ 187 ][ 352 ],
   alphaCSR[ 187 ][ 353 ],
   alphaCSR[ 187 ][ 354 ],
   alphaCSR[ 187 ][ 355 ],
   alphaCSR[ 187 ][ 356 ],
   alphaCSR[ 187 ][ 357 ],
   alphaCSR[ 187 ][ 358 ],
   alphaCSR[ 187 ][ 359 ],
   alphaCSR[ 187 ][ 360 ],
   alphaCSR[ 187 ][ 361 ],
   alphaCSR[ 187 ][ 362 ],
   alphaCSR[ 187 ][ 363 ],
   alphaCSR[ 187 ][ 364 ],
   alphaCSR[ 187 ][ 365 ],
   alphaCSR[ 187 ][ 366 ],
   alphaCSR[ 187 ][ 367 ],
   alphaCSR[ 187 ][ 368 ],
   alphaCSR[ 187 ][ 369 ],
   alphaCSR[ 187 ][ 370 ],
   alphaCSR[ 187 ][ 371 ],
   alphaCSR[ 187 ][ 372 ],
   alphaCSR[ 187 ][ 373 ],
   alphaCSR[ 187 ][ 374 ],
   alphaCSR[ 187 ][ 375 ],
   alphaCSR[ 187 ][ 376 ],
   alphaCSR[ 187 ][ 377 ],
   alphaCSR[ 187 ][ 378 ],
   alphaCSR[ 187 ][ 379 ],
   alphaCSR[ 187 ][ 380 ],
   alphaCSR[ 187 ][ 381 ],
   alphaCSR[ 187 ][ 382 ],
   alphaCSR[ 187 ][ 383 ],
   alphaCSR[ 188 ][ 0 ],
   alphaCSR[ 188 ][ 1 ],
   alphaCSR[ 188 ][ 2 ],
   alphaCSR[ 188 ][ 3 ],
   alphaCSR[ 188 ][ 4 ],
   alphaCSR[ 188 ][ 5 ],
   alphaCSR[ 188 ][ 6 ],
   alphaCSR[ 188 ][ 7 ],
   alphaCSR[ 188 ][ 8 ],
   alphaCSR[ 188 ][ 9 ],
   alphaCSR[ 188 ][ 10 ],
   alphaCSR[ 188 ][ 11 ],
   alphaCSR[ 188 ][ 12 ],
   alphaCSR[ 188 ][ 13 ],
   alphaCSR[ 188 ][ 14 ],
   alphaCSR[ 188 ][ 15 ],
   alphaCSR[ 188 ][ 16 ],
   alphaCSR[ 188 ][ 17 ],
   alphaCSR[ 188 ][ 18 ],
   alphaCSR[ 188 ][ 19 ],
   alphaCSR[ 188 ][ 20 ],
   alphaCSR[ 188 ][ 21 ],
   alphaCSR[ 188 ][ 22 ],
   alphaCSR[ 188 ][ 23 ],
   alphaCSR[ 188 ][ 24 ],
   alphaCSR[ 188 ][ 25 ],
   alphaCSR[ 188 ][ 26 ],
   alphaCSR[ 188 ][ 27 ],
   alphaCSR[ 188 ][ 28 ],
   alphaCSR[ 188 ][ 29 ],
   alphaCSR[ 188 ][ 30 ],
   alphaCSR[ 188 ][ 31 ],
   alphaCSR[ 188 ][ 32 ],
   alphaCSR[ 188 ][ 33 ],
   alphaCSR[ 188 ][ 34 ],
   alphaCSR[ 188 ][ 35 ],
   alphaCSR[ 188 ][ 36 ],
   alphaCSR[ 188 ][ 37 ],
   alphaCSR[ 188 ][ 38 ],
   alphaCSR[ 188 ][ 39 ],
   alphaCSR[ 188 ][ 40 ],
   alphaCSR[ 188 ][ 41 ],
   alphaCSR[ 188 ][ 42 ],
   alphaCSR[ 188 ][ 43 ],
   alphaCSR[ 188 ][ 44 ],
   alphaCSR[ 188 ][ 45 ],
   alphaCSR[ 188 ][ 46 ],
   alphaCSR[ 188 ][ 47 ],
   alphaCSR[ 188 ][ 48 ],
   alphaCSR[ 188 ][ 49 ],
   alphaCSR[ 188 ][ 50 ],
   alphaCSR[ 188 ][ 51 ],
   alphaCSR[ 188 ][ 52 ],
   alphaCSR[ 188 ][ 53 ],
   alphaCSR[ 188 ][ 54 ],
   alphaCSR[ 188 ][ 55 ],
   alphaCSR[ 188 ][ 56 ],
   alphaCSR[ 188 ][ 57 ],
   alphaCSR[ 188 ][ 58 ],
   alphaCSR[ 188 ][ 59 ],
   alphaCSR[ 188 ][ 60 ],
   alphaCSR[ 188 ][ 61 ],
   alphaCSR[ 188 ][ 62 ],
   alphaCSR[ 188 ][ 63 ],
   alphaCSR[ 188 ][ 64 ],
   alphaCSR[ 188 ][ 65 ],
   alphaCSR[ 188 ][ 66 ],
   alphaCSR[ 188 ][ 67 ],
   alphaCSR[ 188 ][ 68 ],
   alphaCSR[ 188 ][ 69 ],
   alphaCSR[ 188 ][ 70 ],
   alphaCSR[ 188 ][ 71 ],
   alphaCSR[ 188 ][ 72 ],
   alphaCSR[ 188 ][ 73 ],
   alphaCSR[ 188 ][ 74 ],
   alphaCSR[ 188 ][ 75 ],
   alphaCSR[ 188 ][ 76 ],
   alphaCSR[ 188 ][ 77 ],
   alphaCSR[ 188 ][ 78 ],
   alphaCSR[ 188 ][ 79 ],
   alphaCSR[ 188 ][ 80 ],
   alphaCSR[ 188 ][ 81 ],
   alphaCSR[ 188 ][ 82 ],
   alphaCSR[ 188 ][ 83 ],
   alphaCSR[ 188 ][ 84 ],
   alphaCSR[ 188 ][ 85 ],
   alphaCSR[ 188 ][ 86 ],
   alphaCSR[ 188 ][ 87 ],
   alphaCSR[ 188 ][ 88 ],
   alphaCSR[ 188 ][ 89 ],
   alphaCSR[ 188 ][ 90 ],
   alphaCSR[ 188 ][ 91 ],
   alphaCSR[ 188 ][ 92 ],
   alphaCSR[ 188 ][ 93 ],
   alphaCSR[ 188 ][ 94 ],
   alphaCSR[ 188 ][ 95 ],
   alphaCSR[ 188 ][ 96 ],
   alphaCSR[ 188 ][ 97 ],
   alphaCSR[ 188 ][ 98 ],
   alphaCSR[ 188 ][ 99 ],
   alphaCSR[ 188 ][ 100 ],
   alphaCSR[ 188 ][ 101 ],
   alphaCSR[ 188 ][ 102 ],
   alphaCSR[ 188 ][ 103 ],
   alphaCSR[ 188 ][ 104 ],
   alphaCSR[ 188 ][ 105 ],
   alphaCSR[ 188 ][ 106 ],
   alphaCSR[ 188 ][ 107 ],
   alphaCSR[ 188 ][ 108 ],
   alphaCSR[ 188 ][ 109 ],
   alphaCSR[ 188 ][ 110 ],
   alphaCSR[ 188 ][ 111 ],
   alphaCSR[ 188 ][ 112 ],
   alphaCSR[ 188 ][ 113 ],
   alphaCSR[ 188 ][ 114 ],
   alphaCSR[ 188 ][ 115 ],
   alphaCSR[ 188 ][ 116 ],
   alphaCSR[ 188 ][ 117 ],
   alphaCSR[ 188 ][ 118 ],
   alphaCSR[ 188 ][ 119 ],
   alphaCSR[ 188 ][ 120 ],
   alphaCSR[ 188 ][ 121 ],
   alphaCSR[ 188 ][ 122 ],
   alphaCSR[ 188 ][ 123 ],
   alphaCSR[ 188 ][ 124 ],
   alphaCSR[ 188 ][ 125 ],
   alphaCSR[ 188 ][ 126 ],
   alphaCSR[ 188 ][ 127 ],
   alphaCSR[ 188 ][ 128 ],
   alphaCSR[ 188 ][ 129 ],
   alphaCSR[ 188 ][ 130 ],
   alphaCSR[ 188 ][ 131 ],
   alphaCSR[ 188 ][ 132 ],
   alphaCSR[ 188 ][ 133 ],
   alphaCSR[ 188 ][ 134 ],
   alphaCSR[ 188 ][ 135 ],
   alphaCSR[ 188 ][ 136 ],
   alphaCSR[ 188 ][ 137 ],
   alphaCSR[ 188 ][ 138 ],
   alphaCSR[ 188 ][ 139 ],
   alphaCSR[ 188 ][ 140 ],
   alphaCSR[ 188 ][ 141 ],
   alphaCSR[ 188 ][ 142 ],
   alphaCSR[ 188 ][ 143 ],
   alphaCSR[ 188 ][ 144 ],
   alphaCSR[ 188 ][ 145 ],
   alphaCSR[ 188 ][ 146 ],
   alphaCSR[ 188 ][ 147 ],
   alphaCSR[ 188 ][ 148 ],
   alphaCSR[ 188 ][ 149 ],
   alphaCSR[ 188 ][ 150 ],
   alphaCSR[ 188 ][ 151 ],
   alphaCSR[ 188 ][ 152 ],
   alphaCSR[ 188 ][ 153 ],
   alphaCSR[ 188 ][ 154 ],
   alphaCSR[ 188 ][ 155 ],
   alphaCSR[ 188 ][ 156 ],
   alphaCSR[ 188 ][ 157 ],
   alphaCSR[ 188 ][ 158 ],
   alphaCSR[ 188 ][ 159 ],
   alphaCSR[ 188 ][ 160 ],
   alphaCSR[ 188 ][ 161 ],
   alphaCSR[ 188 ][ 162 ],
   alphaCSR[ 188 ][ 163 ],
   alphaCSR[ 188 ][ 164 ],
   alphaCSR[ 188 ][ 165 ],
   alphaCSR[ 188 ][ 166 ],
   alphaCSR[ 188 ][ 167 ],
   alphaCSR[ 188 ][ 168 ],
   alphaCSR[ 188 ][ 169 ],
   alphaCSR[ 188 ][ 170 ],
   alphaCSR[ 188 ][ 171 ],
   alphaCSR[ 188 ][ 172 ],
   alphaCSR[ 188 ][ 173 ],
   alphaCSR[ 188 ][ 174 ],
   alphaCSR[ 188 ][ 175 ],
   alphaCSR[ 188 ][ 176 ],
   alphaCSR[ 188 ][ 177 ],
   alphaCSR[ 188 ][ 178 ],
   alphaCSR[ 188 ][ 179 ],
   alphaCSR[ 188 ][ 180 ],
   alphaCSR[ 188 ][ 181 ],
   alphaCSR[ 188 ][ 182 ],
   alphaCSR[ 188 ][ 183 ],
   alphaCSR[ 188 ][ 184 ],
   alphaCSR[ 188 ][ 185 ],
   alphaCSR[ 188 ][ 186 ],
   alphaCSR[ 188 ][ 187 ],
   alphaCSR[ 188 ][ 188 ],
   alphaCSR[ 188 ][ 189 ],
   alphaCSR[ 188 ][ 190 ],
   alphaCSR[ 188 ][ 191 ],
   alphaCSR[ 188 ][ 192 ],
   alphaCSR[ 188 ][ 193 ],
   alphaCSR[ 188 ][ 194 ],
   alphaCSR[ 188 ][ 195 ],
   alphaCSR[ 188 ][ 196 ],
   alphaCSR[ 188 ][ 197 ],
   alphaCSR[ 188 ][ 198 ],
   alphaCSR[ 188 ][ 199 ],
   alphaCSR[ 188 ][ 200 ],
   alphaCSR[ 188 ][ 201 ],
   alphaCSR[ 188 ][ 202 ],
   alphaCSR[ 188 ][ 203 ],
   alphaCSR[ 188 ][ 204 ],
   alphaCSR[ 188 ][ 205 ],
   alphaCSR[ 188 ][ 206 ],
   alphaCSR[ 188 ][ 207 ],
   alphaCSR[ 188 ][ 208 ],
   alphaCSR[ 188 ][ 209 ],
   alphaCSR[ 188 ][ 210 ],
   alphaCSR[ 188 ][ 211 ],
   alphaCSR[ 188 ][ 212 ],
   alphaCSR[ 188 ][ 213 ],
   alphaCSR[ 188 ][ 214 ],
   alphaCSR[ 188 ][ 215 ],
   alphaCSR[ 188 ][ 216 ],
   alphaCSR[ 188 ][ 217 ],
   alphaCSR[ 188 ][ 218 ],
   alphaCSR[ 188 ][ 219 ],
   alphaCSR[ 188 ][ 220 ],
   alphaCSR[ 188 ][ 221 ],
   alphaCSR[ 188 ][ 222 ],
   alphaCSR[ 188 ][ 223 ],
   alphaCSR[ 188 ][ 224 ],
   alphaCSR[ 188 ][ 225 ],
   alphaCSR[ 188 ][ 226 ],
   alphaCSR[ 188 ][ 227 ],
   alphaCSR[ 188 ][ 228 ],
   alphaCSR[ 188 ][ 229 ],
   alphaCSR[ 188 ][ 230 ],
   alphaCSR[ 188 ][ 231 ],
   alphaCSR[ 188 ][ 232 ],
   alphaCSR[ 188 ][ 233 ],
   alphaCSR[ 188 ][ 234 ],
   alphaCSR[ 188 ][ 235 ],
   alphaCSR[ 188 ][ 236 ],
   alphaCSR[ 188 ][ 237 ],
   alphaCSR[ 188 ][ 238 ],
   alphaCSR[ 188 ][ 239 ],
   alphaCSR[ 188 ][ 240 ],
   alphaCSR[ 188 ][ 241 ],
   alphaCSR[ 188 ][ 242 ],
   alphaCSR[ 188 ][ 243 ],
   alphaCSR[ 188 ][ 244 ],
   alphaCSR[ 188 ][ 245 ],
   alphaCSR[ 188 ][ 246 ],
   alphaCSR[ 188 ][ 247 ],
   alphaCSR[ 188 ][ 248 ],
   alphaCSR[ 188 ][ 249 ],
   alphaCSR[ 188 ][ 250 ],
   alphaCSR[ 188 ][ 251 ],
   alphaCSR[ 188 ][ 252 ],
   alphaCSR[ 188 ][ 253 ],
   alphaCSR[ 188 ][ 254 ],
   alphaCSR[ 188 ][ 255 ],
   alphaCSR[ 188 ][ 256 ],
   alphaCSR[ 188 ][ 257 ],
   alphaCSR[ 188 ][ 258 ],
   alphaCSR[ 188 ][ 259 ],
   alphaCSR[ 188 ][ 260 ],
   alphaCSR[ 188 ][ 261 ],
   alphaCSR[ 188 ][ 262 ],
   alphaCSR[ 188 ][ 263 ],
   alphaCSR[ 188 ][ 264 ],
   alphaCSR[ 188 ][ 265 ],
   alphaCSR[ 188 ][ 266 ],
   alphaCSR[ 188 ][ 267 ],
   alphaCSR[ 188 ][ 268 ],
   alphaCSR[ 188 ][ 269 ],
   alphaCSR[ 188 ][ 270 ],
   alphaCSR[ 188 ][ 271 ],
   alphaCSR[ 188 ][ 272 ],
   alphaCSR[ 188 ][ 273 ],
   alphaCSR[ 188 ][ 274 ],
   alphaCSR[ 188 ][ 275 ],
   alphaCSR[ 188 ][ 276 ],
   alphaCSR[ 188 ][ 277 ],
   alphaCSR[ 188 ][ 278 ],
   alphaCSR[ 188 ][ 279 ],
   alphaCSR[ 188 ][ 280 ],
   alphaCSR[ 188 ][ 281 ],
   alphaCSR[ 188 ][ 282 ],
   alphaCSR[ 188 ][ 283 ],
   alphaCSR[ 188 ][ 284 ],
   alphaCSR[ 188 ][ 285 ],
   alphaCSR[ 188 ][ 286 ],
   alphaCSR[ 188 ][ 287 ],
   alphaCSR[ 188 ][ 288 ],
   alphaCSR[ 188 ][ 289 ],
   alphaCSR[ 188 ][ 290 ],
   alphaCSR[ 188 ][ 291 ],
   alphaCSR[ 188 ][ 292 ],
   alphaCSR[ 188 ][ 293 ],
   alphaCSR[ 188 ][ 294 ],
   alphaCSR[ 188 ][ 295 ],
   alphaCSR[ 188 ][ 296 ],
   alphaCSR[ 188 ][ 297 ],
   alphaCSR[ 188 ][ 298 ],
   alphaCSR[ 188 ][ 299 ],
   alphaCSR[ 188 ][ 300 ],
   alphaCSR[ 188 ][ 301 ],
   alphaCSR[ 188 ][ 302 ],
   alphaCSR[ 188 ][ 303 ],
   alphaCSR[ 188 ][ 304 ],
   alphaCSR[ 188 ][ 305 ],
   alphaCSR[ 188 ][ 306 ],
   alphaCSR[ 188 ][ 307 ],
   alphaCSR[ 188 ][ 308 ],
   alphaCSR[ 188 ][ 309 ],
   alphaCSR[ 188 ][ 310 ],
   alphaCSR[ 188 ][ 311 ],
   alphaCSR[ 188 ][ 312 ],
   alphaCSR[ 188 ][ 313 ],
   alphaCSR[ 188 ][ 314 ],
   alphaCSR[ 188 ][ 315 ],
   alphaCSR[ 188 ][ 316 ],
   alphaCSR[ 188 ][ 317 ],
   alphaCSR[ 188 ][ 318 ],
   alphaCSR[ 188 ][ 319 ],
   alphaCSR[ 188 ][ 320 ],
   alphaCSR[ 188 ][ 321 ],
   alphaCSR[ 188 ][ 322 ],
   alphaCSR[ 188 ][ 323 ],
   alphaCSR[ 188 ][ 324 ],
   alphaCSR[ 188 ][ 325 ],
   alphaCSR[ 188 ][ 326 ],
   alphaCSR[ 188 ][ 327 ],
   alphaCSR[ 188 ][ 328 ],
   alphaCSR[ 188 ][ 329 ],
   alphaCSR[ 188 ][ 330 ],
   alphaCSR[ 188 ][ 331 ],
   alphaCSR[ 188 ][ 332 ],
   alphaCSR[ 188 ][ 333 ],
   alphaCSR[ 188 ][ 334 ],
   alphaCSR[ 188 ][ 335 ],
   alphaCSR[ 188 ][ 336 ],
   alphaCSR[ 188 ][ 337 ],
   alphaCSR[ 188 ][ 338 ],
   alphaCSR[ 188 ][ 339 ],
   alphaCSR[ 188 ][ 340 ],
   alphaCSR[ 188 ][ 341 ],
   alphaCSR[ 188 ][ 342 ],
   alphaCSR[ 188 ][ 343 ],
   alphaCSR[ 188 ][ 344 ],
   alphaCSR[ 188 ][ 345 ],
   alphaCSR[ 188 ][ 346 ],
   alphaCSR[ 188 ][ 347 ],
   alphaCSR[ 188 ][ 348 ],
   alphaCSR[ 188 ][ 349 ],
   alphaCSR[ 188 ][ 350 ],
   alphaCSR[ 188 ][ 351 ],
   alphaCSR[ 188 ][ 352 ],
   alphaCSR[ 188 ][ 353 ],
   alphaCSR[ 188 ][ 354 ],
   alphaCSR[ 188 ][ 355 ],
   alphaCSR[ 188 ][ 356 ],
   alphaCSR[ 188 ][ 357 ],
   alphaCSR[ 188 ][ 358 ],
   alphaCSR[ 188 ][ 359 ],
   alphaCSR[ 188 ][ 360 ],
   alphaCSR[ 188 ][ 361 ],
   alphaCSR[ 188 ][ 362 ],
   alphaCSR[ 188 ][ 363 ],
   alphaCSR[ 188 ][ 364 ],
   alphaCSR[ 188 ][ 365 ],
   alphaCSR[ 188 ][ 366 ],
   alphaCSR[ 188 ][ 367 ],
   alphaCSR[ 188 ][ 368 ],
   alphaCSR[ 188 ][ 369 ],
   alphaCSR[ 188 ][ 370 ],
   alphaCSR[ 188 ][ 371 ],
   alphaCSR[ 188 ][ 372 ],
   alphaCSR[ 188 ][ 373 ],
   alphaCSR[ 188 ][ 374 ],
   alphaCSR[ 188 ][ 375 ],
   alphaCSR[ 188 ][ 376 ],
   alphaCSR[ 188 ][ 377 ],
   alphaCSR[ 188 ][ 378 ],
   alphaCSR[ 188 ][ 379 ],
   alphaCSR[ 188 ][ 380 ],
   alphaCSR[ 188 ][ 381 ],
   alphaCSR[ 188 ][ 382 ],
   alphaCSR[ 188 ][ 383 ],
   alphaCSR[ 189 ][ 0 ],
   alphaCSR[ 189 ][ 1 ],
   alphaCSR[ 189 ][ 2 ],
   alphaCSR[ 189 ][ 3 ],
   alphaCSR[ 189 ][ 4 ],
   alphaCSR[ 189 ][ 5 ],
   alphaCSR[ 189 ][ 6 ],
   alphaCSR[ 189 ][ 7 ],
   alphaCSR[ 189 ][ 8 ],
   alphaCSR[ 189 ][ 9 ],
   alphaCSR[ 189 ][ 10 ],
   alphaCSR[ 189 ][ 11 ],
   alphaCSR[ 189 ][ 12 ],
   alphaCSR[ 189 ][ 13 ],
   alphaCSR[ 189 ][ 14 ],
   alphaCSR[ 189 ][ 15 ],
   alphaCSR[ 189 ][ 16 ],
   alphaCSR[ 189 ][ 17 ],
   alphaCSR[ 189 ][ 18 ],
   alphaCSR[ 189 ][ 19 ],
   alphaCSR[ 189 ][ 20 ],
   alphaCSR[ 189 ][ 21 ],
   alphaCSR[ 189 ][ 22 ],
   alphaCSR[ 189 ][ 23 ],
   alphaCSR[ 189 ][ 24 ],
   alphaCSR[ 189 ][ 25 ],
   alphaCSR[ 189 ][ 26 ],
   alphaCSR[ 189 ][ 27 ],
   alphaCSR[ 189 ][ 28 ],
   alphaCSR[ 189 ][ 29 ],
   alphaCSR[ 189 ][ 30 ],
   alphaCSR[ 189 ][ 31 ],
   alphaCSR[ 189 ][ 32 ],
   alphaCSR[ 189 ][ 33 ],
   alphaCSR[ 189 ][ 34 ],
   alphaCSR[ 189 ][ 35 ],
   alphaCSR[ 189 ][ 36 ],
   alphaCSR[ 189 ][ 37 ],
   alphaCSR[ 189 ][ 38 ],
   alphaCSR[ 189 ][ 39 ],
   alphaCSR[ 189 ][ 40 ],
   alphaCSR[ 189 ][ 41 ],
   alphaCSR[ 189 ][ 42 ],
   alphaCSR[ 189 ][ 43 ],
   alphaCSR[ 189 ][ 44 ],
   alphaCSR[ 189 ][ 45 ],
   alphaCSR[ 189 ][ 46 ],
   alphaCSR[ 189 ][ 47 ],
   alphaCSR[ 189 ][ 48 ],
   alphaCSR[ 189 ][ 49 ],
   alphaCSR[ 189 ][ 50 ],
   alphaCSR[ 189 ][ 51 ],
   alphaCSR[ 189 ][ 52 ],
   alphaCSR[ 189 ][ 53 ],
   alphaCSR[ 189 ][ 54 ],
   alphaCSR[ 189 ][ 55 ],
   alphaCSR[ 189 ][ 56 ],
   alphaCSR[ 189 ][ 57 ],
   alphaCSR[ 189 ][ 58 ],
   alphaCSR[ 189 ][ 59 ],
   alphaCSR[ 189 ][ 60 ],
   alphaCSR[ 189 ][ 61 ],
   alphaCSR[ 189 ][ 62 ],
   alphaCSR[ 189 ][ 63 ],
   alphaCSR[ 189 ][ 64 ],
   alphaCSR[ 189 ][ 65 ],
   alphaCSR[ 189 ][ 66 ],
   alphaCSR[ 189 ][ 67 ],
   alphaCSR[ 189 ][ 68 ],
   alphaCSR[ 189 ][ 69 ],
   alphaCSR[ 189 ][ 70 ],
   alphaCSR[ 189 ][ 71 ],
   alphaCSR[ 189 ][ 72 ],
   alphaCSR[ 189 ][ 73 ],
   alphaCSR[ 189 ][ 74 ],
   alphaCSR[ 189 ][ 75 ],
   alphaCSR[ 189 ][ 76 ],
   alphaCSR[ 189 ][ 77 ],
   alphaCSR[ 189 ][ 78 ],
   alphaCSR[ 189 ][ 79 ],
   alphaCSR[ 189 ][ 80 ],
   alphaCSR[ 189 ][ 81 ],
   alphaCSR[ 189 ][ 82 ],
   alphaCSR[ 189 ][ 83 ],
   alphaCSR[ 189 ][ 84 ],
   alphaCSR[ 189 ][ 85 ],
   alphaCSR[ 189 ][ 86 ],
   alphaCSR[ 189 ][ 87 ],
   alphaCSR[ 189 ][ 88 ],
   alphaCSR[ 189 ][ 89 ],
   alphaCSR[ 189 ][ 90 ],
   alphaCSR[ 189 ][ 91 ],
   alphaCSR[ 189 ][ 92 ],
   alphaCSR[ 189 ][ 93 ],
   alphaCSR[ 189 ][ 94 ],
   alphaCSR[ 189 ][ 95 ],
   alphaCSR[ 189 ][ 96 ],
   alphaCSR[ 189 ][ 97 ],
   alphaCSR[ 189 ][ 98 ],
   alphaCSR[ 189 ][ 99 ],
   alphaCSR[ 189 ][ 100 ],
   alphaCSR[ 189 ][ 101 ],
   alphaCSR[ 189 ][ 102 ],
   alphaCSR[ 189 ][ 103 ],
   alphaCSR[ 189 ][ 104 ],
   alphaCSR[ 189 ][ 105 ],
   alphaCSR[ 189 ][ 106 ],
   alphaCSR[ 189 ][ 107 ],
   alphaCSR[ 189 ][ 108 ],
   alphaCSR[ 189 ][ 109 ],
   alphaCSR[ 189 ][ 110 ],
   alphaCSR[ 189 ][ 111 ],
   alphaCSR[ 189 ][ 112 ],
   alphaCSR[ 189 ][ 113 ],
   alphaCSR[ 189 ][ 114 ],
   alphaCSR[ 189 ][ 115 ],
   alphaCSR[ 189 ][ 116 ],
   alphaCSR[ 189 ][ 117 ],
   alphaCSR[ 189 ][ 118 ],
   alphaCSR[ 189 ][ 119 ],
   alphaCSR[ 189 ][ 120 ],
   alphaCSR[ 189 ][ 121 ],
   alphaCSR[ 189 ][ 122 ],
   alphaCSR[ 189 ][ 123 ],
   alphaCSR[ 189 ][ 124 ],
   alphaCSR[ 189 ][ 125 ],
   alphaCSR[ 189 ][ 126 ],
   alphaCSR[ 189 ][ 127 ],
   alphaCSR[ 189 ][ 128 ],
   alphaCSR[ 189 ][ 129 ],
   alphaCSR[ 189 ][ 130 ],
   alphaCSR[ 189 ][ 131 ],
   alphaCSR[ 189 ][ 132 ],
   alphaCSR[ 189 ][ 133 ],
   alphaCSR[ 189 ][ 134 ],
   alphaCSR[ 189 ][ 135 ],
   alphaCSR[ 189 ][ 136 ],
   alphaCSR[ 189 ][ 137 ],
   alphaCSR[ 189 ][ 138 ],
   alphaCSR[ 189 ][ 139 ],
   alphaCSR[ 189 ][ 140 ],
   alphaCSR[ 189 ][ 141 ],
   alphaCSR[ 189 ][ 142 ],
   alphaCSR[ 189 ][ 143 ],
   alphaCSR[ 189 ][ 144 ],
   alphaCSR[ 189 ][ 145 ],
   alphaCSR[ 189 ][ 146 ],
   alphaCSR[ 189 ][ 147 ],
   alphaCSR[ 189 ][ 148 ],
   alphaCSR[ 189 ][ 149 ],
   alphaCSR[ 189 ][ 150 ],
   alphaCSR[ 189 ][ 151 ],
   alphaCSR[ 189 ][ 152 ],
   alphaCSR[ 189 ][ 153 ],
   alphaCSR[ 189 ][ 154 ],
   alphaCSR[ 189 ][ 155 ],
   alphaCSR[ 189 ][ 156 ],
   alphaCSR[ 189 ][ 157 ],
   alphaCSR[ 189 ][ 158 ],
   alphaCSR[ 189 ][ 159 ],
   alphaCSR[ 189 ][ 160 ],
   alphaCSR[ 189 ][ 161 ],
   alphaCSR[ 189 ][ 162 ],
   alphaCSR[ 189 ][ 163 ],
   alphaCSR[ 189 ][ 164 ],
   alphaCSR[ 189 ][ 165 ],
   alphaCSR[ 189 ][ 166 ],
   alphaCSR[ 189 ][ 167 ],
   alphaCSR[ 189 ][ 168 ],
   alphaCSR[ 189 ][ 169 ],
   alphaCSR[ 189 ][ 170 ],
   alphaCSR[ 189 ][ 171 ],
   alphaCSR[ 189 ][ 172 ],
   alphaCSR[ 189 ][ 173 ],
   alphaCSR[ 189 ][ 174 ],
   alphaCSR[ 189 ][ 175 ],
   alphaCSR[ 189 ][ 176 ],
   alphaCSR[ 189 ][ 177 ],
   alphaCSR[ 189 ][ 178 ],
   alphaCSR[ 189 ][ 179 ],
   alphaCSR[ 189 ][ 180 ],
   alphaCSR[ 189 ][ 181 ],
   alphaCSR[ 189 ][ 182 ],
   alphaCSR[ 189 ][ 183 ],
   alphaCSR[ 189 ][ 184 ],
   alphaCSR[ 189 ][ 185 ],
   alphaCSR[ 189 ][ 186 ],
   alphaCSR[ 189 ][ 187 ],
   alphaCSR[ 189 ][ 188 ],
   alphaCSR[ 189 ][ 189 ],
   alphaCSR[ 189 ][ 190 ],
   alphaCSR[ 189 ][ 191 ],
   alphaCSR[ 189 ][ 192 ],
   alphaCSR[ 189 ][ 193 ],
   alphaCSR[ 189 ][ 194 ],
   alphaCSR[ 189 ][ 195 ],
   alphaCSR[ 189 ][ 196 ],
   alphaCSR[ 189 ][ 197 ],
   alphaCSR[ 189 ][ 198 ],
   alphaCSR[ 189 ][ 199 ],
   alphaCSR[ 189 ][ 200 ],
   alphaCSR[ 189 ][ 201 ],
   alphaCSR[ 189 ][ 202 ],
   alphaCSR[ 189 ][ 203 ],
   alphaCSR[ 189 ][ 204 ],
   alphaCSR[ 189 ][ 205 ],
   alphaCSR[ 189 ][ 206 ],
   alphaCSR[ 189 ][ 207 ],
   alphaCSR[ 189 ][ 208 ],
   alphaCSR[ 189 ][ 209 ],
   alphaCSR[ 189 ][ 210 ],
   alphaCSR[ 189 ][ 211 ],
   alphaCSR[ 189 ][ 212 ],
   alphaCSR[ 189 ][ 213 ],
   alphaCSR[ 189 ][ 214 ],
   alphaCSR[ 189 ][ 215 ],
   alphaCSR[ 189 ][ 216 ],
   alphaCSR[ 189 ][ 217 ],
   alphaCSR[ 189 ][ 218 ],
   alphaCSR[ 189 ][ 219 ],
   alphaCSR[ 189 ][ 220 ],
   alphaCSR[ 189 ][ 221 ],
   alphaCSR[ 189 ][ 222 ],
   alphaCSR[ 189 ][ 223 ],
   alphaCSR[ 189 ][ 224 ],
   alphaCSR[ 189 ][ 225 ],
   alphaCSR[ 189 ][ 226 ],
   alphaCSR[ 189 ][ 227 ],
   alphaCSR[ 189 ][ 228 ],
   alphaCSR[ 189 ][ 229 ],
   alphaCSR[ 189 ][ 230 ],
   alphaCSR[ 189 ][ 231 ],
   alphaCSR[ 189 ][ 232 ],
   alphaCSR[ 189 ][ 233 ],
   alphaCSR[ 189 ][ 234 ],
   alphaCSR[ 189 ][ 235 ],
   alphaCSR[ 189 ][ 236 ],
   alphaCSR[ 189 ][ 237 ],
   alphaCSR[ 189 ][ 238 ],
   alphaCSR[ 189 ][ 239 ],
   alphaCSR[ 189 ][ 240 ],
   alphaCSR[ 189 ][ 241 ],
   alphaCSR[ 189 ][ 242 ],
   alphaCSR[ 189 ][ 243 ],
   alphaCSR[ 189 ][ 244 ],
   alphaCSR[ 189 ][ 245 ],
   alphaCSR[ 189 ][ 246 ],
   alphaCSR[ 189 ][ 247 ],
   alphaCSR[ 189 ][ 248 ],
   alphaCSR[ 189 ][ 249 ],
   alphaCSR[ 189 ][ 250 ],
   alphaCSR[ 189 ][ 251 ],
   alphaCSR[ 189 ][ 252 ],
   alphaCSR[ 189 ][ 253 ],
   alphaCSR[ 189 ][ 254 ],
   alphaCSR[ 189 ][ 255 ],
   alphaCSR[ 189 ][ 256 ],
   alphaCSR[ 189 ][ 257 ],
   alphaCSR[ 189 ][ 258 ],
   alphaCSR[ 189 ][ 259 ],
   alphaCSR[ 189 ][ 260 ],
   alphaCSR[ 189 ][ 261 ],
   alphaCSR[ 189 ][ 262 ],
   alphaCSR[ 189 ][ 263 ],
   alphaCSR[ 189 ][ 264 ],
   alphaCSR[ 189 ][ 265 ],
   alphaCSR[ 189 ][ 266 ],
   alphaCSR[ 189 ][ 267 ],
   alphaCSR[ 189 ][ 268 ],
   alphaCSR[ 189 ][ 269 ],
   alphaCSR[ 189 ][ 270 ],
   alphaCSR[ 189 ][ 271 ],
   alphaCSR[ 189 ][ 272 ],
   alphaCSR[ 189 ][ 273 ],
   alphaCSR[ 189 ][ 274 ],
   alphaCSR[ 189 ][ 275 ],
   alphaCSR[ 189 ][ 276 ],
   alphaCSR[ 189 ][ 277 ],
   alphaCSR[ 189 ][ 278 ],
   alphaCSR[ 189 ][ 279 ],
   alphaCSR[ 189 ][ 280 ],
   alphaCSR[ 189 ][ 281 ],
   alphaCSR[ 189 ][ 282 ],
   alphaCSR[ 189 ][ 283 ],
   alphaCSR[ 189 ][ 284 ],
   alphaCSR[ 189 ][ 285 ],
   alphaCSR[ 189 ][ 286 ],
   alphaCSR[ 189 ][ 287 ],
   alphaCSR[ 189 ][ 288 ],
   alphaCSR[ 189 ][ 289 ],
   alphaCSR[ 189 ][ 290 ],
   alphaCSR[ 189 ][ 291 ],
   alphaCSR[ 189 ][ 292 ],
   alphaCSR[ 189 ][ 293 ],
   alphaCSR[ 189 ][ 294 ],
   alphaCSR[ 189 ][ 295 ],
   alphaCSR[ 189 ][ 296 ],
   alphaCSR[ 189 ][ 297 ],
   alphaCSR[ 189 ][ 298 ],
   alphaCSR[ 189 ][ 299 ],
   alphaCSR[ 189 ][ 300 ],
   alphaCSR[ 189 ][ 301 ],
   alphaCSR[ 189 ][ 302 ],
   alphaCSR[ 189 ][ 303 ],
   alphaCSR[ 189 ][ 304 ],
   alphaCSR[ 189 ][ 305 ],
   alphaCSR[ 189 ][ 306 ],
   alphaCSR[ 189 ][ 307 ],
   alphaCSR[ 189 ][ 308 ],
   alphaCSR[ 189 ][ 309 ],
   alphaCSR[ 189 ][ 310 ],
   alphaCSR[ 189 ][ 311 ],
   alphaCSR[ 189 ][ 312 ],
   alphaCSR[ 189 ][ 313 ],
   alphaCSR[ 189 ][ 314 ],
   alphaCSR[ 189 ][ 315 ],
   alphaCSR[ 189 ][ 316 ],
   alphaCSR[ 189 ][ 317 ],
   alphaCSR[ 189 ][ 318 ],
   alphaCSR[ 189 ][ 319 ],
   alphaCSR[ 189 ][ 320 ],
   alphaCSR[ 189 ][ 321 ],
   alphaCSR[ 189 ][ 322 ],
   alphaCSR[ 189 ][ 323 ],
   alphaCSR[ 189 ][ 324 ],
   alphaCSR[ 189 ][ 325 ],
   alphaCSR[ 189 ][ 326 ],
   alphaCSR[ 189 ][ 327 ],
   alphaCSR[ 189 ][ 328 ],
   alphaCSR[ 189 ][ 329 ],
   alphaCSR[ 189 ][ 330 ],
   alphaCSR[ 189 ][ 331 ],
   alphaCSR[ 189 ][ 332 ],
   alphaCSR[ 189 ][ 333 ],
   alphaCSR[ 189 ][ 334 ],
   alphaCSR[ 189 ][ 335 ],
   alphaCSR[ 189 ][ 336 ],
   alphaCSR[ 189 ][ 337 ],
   alphaCSR[ 189 ][ 338 ],
   alphaCSR[ 189 ][ 339 ],
   alphaCSR[ 189 ][ 340 ],
   alphaCSR[ 189 ][ 341 ],
   alphaCSR[ 189 ][ 342 ],
   alphaCSR[ 189 ][ 343 ],
   alphaCSR[ 189 ][ 344 ],
   alphaCSR[ 189 ][ 345 ],
   alphaCSR[ 189 ][ 346 ],
   alphaCSR[ 189 ][ 347 ],
   alphaCSR[ 189 ][ 348 ],
   alphaCSR[ 189 ][ 349 ],
   alphaCSR[ 189 ][ 350 ],
   alphaCSR[ 189 ][ 351 ],
   alphaCSR[ 189 ][ 352 ],
   alphaCSR[ 189 ][ 353 ],
   alphaCSR[ 189 ][ 354 ],
   alphaCSR[ 189 ][ 355 ],
   alphaCSR[ 189 ][ 356 ],
   alphaCSR[ 189 ][ 357 ],
   alphaCSR[ 189 ][ 358 ],
   alphaCSR[ 189 ][ 359 ],
   alphaCSR[ 189 ][ 360 ],
   alphaCSR[ 189 ][ 361 ],
   alphaCSR[ 189 ][ 362 ],
   alphaCSR[ 189 ][ 363 ],
   alphaCSR[ 189 ][ 364 ],
   alphaCSR[ 189 ][ 365 ],
   alphaCSR[ 189 ][ 366 ],
   alphaCSR[ 189 ][ 367 ],
   alphaCSR[ 189 ][ 368 ],
   alphaCSR[ 189 ][ 369 ],
   alphaCSR[ 189 ][ 370 ],
   alphaCSR[ 189 ][ 371 ],
   alphaCSR[ 189 ][ 372 ],
   alphaCSR[ 189 ][ 373 ],
   alphaCSR[ 189 ][ 374 ],
   alphaCSR[ 189 ][ 375 ],
   alphaCSR[ 189 ][ 376 ],
   alphaCSR[ 189 ][ 377 ],
   alphaCSR[ 189 ][ 378 ],
   alphaCSR[ 189 ][ 379 ],
   alphaCSR[ 189 ][ 380 ],
   alphaCSR[ 189 ][ 381 ],
   alphaCSR[ 189 ][ 382 ],
   alphaCSR[ 189 ][ 383 ],
   alphaCSR[ 190 ][ 0 ],
   alphaCSR[ 190 ][ 1 ],
   alphaCSR[ 190 ][ 2 ],
   alphaCSR[ 190 ][ 3 ],
   alphaCSR[ 190 ][ 4 ],
   alphaCSR[ 190 ][ 5 ],
   alphaCSR[ 190 ][ 6 ],
   alphaCSR[ 190 ][ 7 ],
   alphaCSR[ 190 ][ 8 ],
   alphaCSR[ 190 ][ 9 ],
   alphaCSR[ 190 ][ 10 ],
   alphaCSR[ 190 ][ 11 ],
   alphaCSR[ 190 ][ 12 ],
   alphaCSR[ 190 ][ 13 ],
   alphaCSR[ 190 ][ 14 ],
   alphaCSR[ 190 ][ 15 ],
   alphaCSR[ 190 ][ 16 ],
   alphaCSR[ 190 ][ 17 ],
   alphaCSR[ 190 ][ 18 ],
   alphaCSR[ 190 ][ 19 ],
   alphaCSR[ 190 ][ 20 ],
   alphaCSR[ 190 ][ 21 ],
   alphaCSR[ 190 ][ 22 ],
   alphaCSR[ 190 ][ 23 ],
   alphaCSR[ 190 ][ 24 ],
   alphaCSR[ 190 ][ 25 ],
   alphaCSR[ 190 ][ 26 ],
   alphaCSR[ 190 ][ 27 ],
   alphaCSR[ 190 ][ 28 ],
   alphaCSR[ 190 ][ 29 ],
   alphaCSR[ 190 ][ 30 ],
   alphaCSR[ 190 ][ 31 ],
   alphaCSR[ 190 ][ 32 ],
   alphaCSR[ 190 ][ 33 ],
   alphaCSR[ 190 ][ 34 ],
   alphaCSR[ 190 ][ 35 ],
   alphaCSR[ 190 ][ 36 ],
   alphaCSR[ 190 ][ 37 ],
   alphaCSR[ 190 ][ 38 ],
   alphaCSR[ 190 ][ 39 ],
   alphaCSR[ 190 ][ 40 ],
   alphaCSR[ 190 ][ 41 ],
   alphaCSR[ 190 ][ 42 ],
   alphaCSR[ 190 ][ 43 ],
   alphaCSR[ 190 ][ 44 ],
   alphaCSR[ 190 ][ 45 ],
   alphaCSR[ 190 ][ 46 ],
   alphaCSR[ 190 ][ 47 ],
   alphaCSR[ 190 ][ 48 ],
   alphaCSR[ 190 ][ 49 ],
   alphaCSR[ 190 ][ 50 ],
   alphaCSR[ 190 ][ 51 ],
   alphaCSR[ 190 ][ 52 ],
   alphaCSR[ 190 ][ 53 ],
   alphaCSR[ 190 ][ 54 ],
   alphaCSR[ 190 ][ 55 ],
   alphaCSR[ 190 ][ 56 ],
   alphaCSR[ 190 ][ 57 ],
   alphaCSR[ 190 ][ 58 ],
   alphaCSR[ 190 ][ 59 ],
   alphaCSR[ 190 ][ 60 ],
   alphaCSR[ 190 ][ 61 ],
   alphaCSR[ 190 ][ 62 ],
   alphaCSR[ 190 ][ 63 ],
   alphaCSR[ 190 ][ 64 ],
   alphaCSR[ 190 ][ 65 ],
   alphaCSR[ 190 ][ 66 ],
   alphaCSR[ 190 ][ 67 ],
   alphaCSR[ 190 ][ 68 ],
   alphaCSR[ 190 ][ 69 ],
   alphaCSR[ 190 ][ 70 ],
   alphaCSR[ 190 ][ 71 ],
   alphaCSR[ 190 ][ 72 ],
   alphaCSR[ 190 ][ 73 ],
   alphaCSR[ 190 ][ 74 ],
   alphaCSR[ 190 ][ 75 ],
   alphaCSR[ 190 ][ 76 ],
   alphaCSR[ 190 ][ 77 ],
   alphaCSR[ 190 ][ 78 ],
   alphaCSR[ 190 ][ 79 ],
   alphaCSR[ 190 ][ 80 ],
   alphaCSR[ 190 ][ 81 ],
   alphaCSR[ 190 ][ 82 ],
   alphaCSR[ 190 ][ 83 ],
   alphaCSR[ 190 ][ 84 ],
   alphaCSR[ 190 ][ 85 ],
   alphaCSR[ 190 ][ 86 ],
   alphaCSR[ 190 ][ 87 ],
   alphaCSR[ 190 ][ 88 ],
   alphaCSR[ 190 ][ 89 ],
   alphaCSR[ 190 ][ 90 ],
   alphaCSR[ 190 ][ 91 ],
   alphaCSR[ 190 ][ 92 ],
   alphaCSR[ 190 ][ 93 ],
   alphaCSR[ 190 ][ 94 ],
   alphaCSR[ 190 ][ 95 ],
   alphaCSR[ 190 ][ 96 ],
   alphaCSR[ 190 ][ 97 ],
   alphaCSR[ 190 ][ 98 ],
   alphaCSR[ 190 ][ 99 ],
   alphaCSR[ 190 ][ 100 ],
   alphaCSR[ 190 ][ 101 ],
   alphaCSR[ 190 ][ 102 ],
   alphaCSR[ 190 ][ 103 ],
   alphaCSR[ 190 ][ 104 ],
   alphaCSR[ 190 ][ 105 ],
   alphaCSR[ 190 ][ 106 ],
   alphaCSR[ 190 ][ 107 ],
   alphaCSR[ 190 ][ 108 ],
   alphaCSR[ 190 ][ 109 ],
   alphaCSR[ 190 ][ 110 ],
   alphaCSR[ 190 ][ 111 ],
   alphaCSR[ 190 ][ 112 ],
   alphaCSR[ 190 ][ 113 ],
   alphaCSR[ 190 ][ 114 ],
   alphaCSR[ 190 ][ 115 ],
   alphaCSR[ 190 ][ 116 ],
   alphaCSR[ 190 ][ 117 ],
   alphaCSR[ 190 ][ 118 ],
   alphaCSR[ 190 ][ 119 ],
   alphaCSR[ 190 ][ 120 ],
   alphaCSR[ 190 ][ 121 ],
   alphaCSR[ 190 ][ 122 ],
   alphaCSR[ 190 ][ 123 ],
   alphaCSR[ 190 ][ 124 ],
   alphaCSR[ 190 ][ 125 ],
   alphaCSR[ 190 ][ 126 ],
   alphaCSR[ 190 ][ 127 ],
   alphaCSR[ 190 ][ 128 ],
   alphaCSR[ 190 ][ 129 ],
   alphaCSR[ 190 ][ 130 ],
   alphaCSR[ 190 ][ 131 ],
   alphaCSR[ 190 ][ 132 ],
   alphaCSR[ 190 ][ 133 ],
   alphaCSR[ 190 ][ 134 ],
   alphaCSR[ 190 ][ 135 ],
   alphaCSR[ 190 ][ 136 ],
   alphaCSR[ 190 ][ 137 ],
   alphaCSR[ 190 ][ 138 ],
   alphaCSR[ 190 ][ 139 ],
   alphaCSR[ 190 ][ 140 ],
   alphaCSR[ 190 ][ 141 ],
   alphaCSR[ 190 ][ 142 ],
   alphaCSR[ 190 ][ 143 ],
   alphaCSR[ 190 ][ 144 ],
   alphaCSR[ 190 ][ 145 ],
   alphaCSR[ 190 ][ 146 ],
   alphaCSR[ 190 ][ 147 ],
   alphaCSR[ 190 ][ 148 ],
   alphaCSR[ 190 ][ 149 ],
   alphaCSR[ 190 ][ 150 ],
   alphaCSR[ 190 ][ 151 ],
   alphaCSR[ 190 ][ 152 ],
   alphaCSR[ 190 ][ 153 ],
   alphaCSR[ 190 ][ 154 ],
   alphaCSR[ 190 ][ 155 ],
   alphaCSR[ 190 ][ 156 ],
   alphaCSR[ 190 ][ 157 ],
   alphaCSR[ 190 ][ 158 ],
   alphaCSR[ 190 ][ 159 ],
   alphaCSR[ 190 ][ 160 ],
   alphaCSR[ 190 ][ 161 ],
   alphaCSR[ 190 ][ 162 ],
   alphaCSR[ 190 ][ 163 ],
   alphaCSR[ 190 ][ 164 ],
   alphaCSR[ 190 ][ 165 ],
   alphaCSR[ 190 ][ 166 ],
   alphaCSR[ 190 ][ 167 ],
   alphaCSR[ 190 ][ 168 ],
   alphaCSR[ 190 ][ 169 ],
   alphaCSR[ 190 ][ 170 ],
   alphaCSR[ 190 ][ 171 ],
   alphaCSR[ 190 ][ 172 ],
   alphaCSR[ 190 ][ 173 ],
   alphaCSR[ 190 ][ 174 ],
   alphaCSR[ 190 ][ 175 ],
   alphaCSR[ 190 ][ 176 ],
   alphaCSR[ 190 ][ 177 ],
   alphaCSR[ 190 ][ 178 ],
   alphaCSR[ 190 ][ 179 ],
   alphaCSR[ 190 ][ 180 ],
   alphaCSR[ 190 ][ 181 ],
   alphaCSR[ 190 ][ 182 ],
   alphaCSR[ 190 ][ 183 ],
   alphaCSR[ 190 ][ 184 ],
   alphaCSR[ 190 ][ 185 ],
   alphaCSR[ 190 ][ 186 ],
   alphaCSR[ 190 ][ 187 ],
   alphaCSR[ 190 ][ 188 ],
   alphaCSR[ 190 ][ 189 ],
   alphaCSR[ 190 ][ 190 ],
   alphaCSR[ 190 ][ 191 ],
   alphaCSR[ 190 ][ 192 ],
   alphaCSR[ 190 ][ 193 ],
   alphaCSR[ 190 ][ 194 ],
   alphaCSR[ 190 ][ 195 ],
   alphaCSR[ 190 ][ 196 ],
   alphaCSR[ 190 ][ 197 ],
   alphaCSR[ 190 ][ 198 ],
   alphaCSR[ 190 ][ 199 ],
   alphaCSR[ 190 ][ 200 ],
   alphaCSR[ 190 ][ 201 ],
   alphaCSR[ 190 ][ 202 ],
   alphaCSR[ 190 ][ 203 ],
   alphaCSR[ 190 ][ 204 ],
   alphaCSR[ 190 ][ 205 ],
   alphaCSR[ 190 ][ 206 ],
   alphaCSR[ 190 ][ 207 ],
   alphaCSR[ 190 ][ 208 ],
   alphaCSR[ 190 ][ 209 ],
   alphaCSR[ 190 ][ 210 ],
   alphaCSR[ 190 ][ 211 ],
   alphaCSR[ 190 ][ 212 ],
   alphaCSR[ 190 ][ 213 ],
   alphaCSR[ 190 ][ 214 ],
   alphaCSR[ 190 ][ 215 ],
   alphaCSR[ 190 ][ 216 ],
   alphaCSR[ 190 ][ 217 ],
   alphaCSR[ 190 ][ 218 ],
   alphaCSR[ 190 ][ 219 ],
   alphaCSR[ 190 ][ 220 ],
   alphaCSR[ 190 ][ 221 ],
   alphaCSR[ 190 ][ 222 ],
   alphaCSR[ 190 ][ 223 ],
   alphaCSR[ 190 ][ 224 ],
   alphaCSR[ 190 ][ 225 ],
   alphaCSR[ 190 ][ 226 ],
   alphaCSR[ 190 ][ 227 ],
   alphaCSR[ 190 ][ 228 ],
   alphaCSR[ 190 ][ 229 ],
   alphaCSR[ 190 ][ 230 ],
   alphaCSR[ 190 ][ 231 ],
   alphaCSR[ 190 ][ 232 ],
   alphaCSR[ 190 ][ 233 ],
   alphaCSR[ 190 ][ 234 ],
   alphaCSR[ 190 ][ 235 ],
   alphaCSR[ 190 ][ 236 ],
   alphaCSR[ 190 ][ 237 ],
   alphaCSR[ 190 ][ 238 ],
   alphaCSR[ 190 ][ 239 ],
   alphaCSR[ 190 ][ 240 ],
   alphaCSR[ 190 ][ 241 ],
   alphaCSR[ 190 ][ 242 ],
   alphaCSR[ 190 ][ 243 ],
   alphaCSR[ 190 ][ 244 ],
   alphaCSR[ 190 ][ 245 ],
   alphaCSR[ 190 ][ 246 ],
   alphaCSR[ 190 ][ 247 ],
   alphaCSR[ 190 ][ 248 ],
   alphaCSR[ 190 ][ 249 ],
   alphaCSR[ 190 ][ 250 ],
   alphaCSR[ 190 ][ 251 ],
   alphaCSR[ 190 ][ 252 ],
   alphaCSR[ 190 ][ 253 ],
   alphaCSR[ 190 ][ 254 ],
   alphaCSR[ 190 ][ 255 ],
   alphaCSR[ 190 ][ 256 ],
   alphaCSR[ 190 ][ 257 ],
   alphaCSR[ 190 ][ 258 ],
   alphaCSR[ 190 ][ 259 ],
   alphaCSR[ 190 ][ 260 ],
   alphaCSR[ 190 ][ 261 ],
   alphaCSR[ 190 ][ 262 ],
   alphaCSR[ 190 ][ 263 ],
   alphaCSR[ 190 ][ 264 ],
   alphaCSR[ 190 ][ 265 ],
   alphaCSR[ 190 ][ 266 ],
   alphaCSR[ 190 ][ 267 ],
   alphaCSR[ 190 ][ 268 ],
   alphaCSR[ 190 ][ 269 ],
   alphaCSR[ 190 ][ 270 ],
   alphaCSR[ 190 ][ 271 ],
   alphaCSR[ 190 ][ 272 ],
   alphaCSR[ 190 ][ 273 ],
   alphaCSR[ 190 ][ 274 ],
   alphaCSR[ 190 ][ 275 ],
   alphaCSR[ 190 ][ 276 ],
   alphaCSR[ 190 ][ 277 ],
   alphaCSR[ 190 ][ 278 ],
   alphaCSR[ 190 ][ 279 ],
   alphaCSR[ 190 ][ 280 ],
   alphaCSR[ 190 ][ 281 ],
   alphaCSR[ 190 ][ 282 ],
   alphaCSR[ 190 ][ 283 ],
   alphaCSR[ 190 ][ 284 ],
   alphaCSR[ 190 ][ 285 ],
   alphaCSR[ 190 ][ 286 ],
   alphaCSR[ 190 ][ 287 ],
   alphaCSR[ 190 ][ 288 ],
   alphaCSR[ 190 ][ 289 ],
   alphaCSR[ 190 ][ 290 ],
   alphaCSR[ 190 ][ 291 ],
   alphaCSR[ 190 ][ 292 ],
   alphaCSR[ 190 ][ 293 ],
   alphaCSR[ 190 ][ 294 ],
   alphaCSR[ 190 ][ 295 ],
   alphaCSR[ 190 ][ 296 ],
   alphaCSR[ 190 ][ 297 ],
   alphaCSR[ 190 ][ 298 ],
   alphaCSR[ 190 ][ 299 ],
   alphaCSR[ 190 ][ 300 ],
   alphaCSR[ 190 ][ 301 ],
   alphaCSR[ 190 ][ 302 ],
   alphaCSR[ 190 ][ 303 ],
   alphaCSR[ 190 ][ 304 ],
   alphaCSR[ 190 ][ 305 ],
   alphaCSR[ 190 ][ 306 ],
   alphaCSR[ 190 ][ 307 ],
   alphaCSR[ 190 ][ 308 ],
   alphaCSR[ 190 ][ 309 ],
   alphaCSR[ 190 ][ 310 ],
   alphaCSR[ 190 ][ 311 ],
   alphaCSR[ 190 ][ 312 ],
   alphaCSR[ 190 ][ 313 ],
   alphaCSR[ 190 ][ 314 ],
   alphaCSR[ 190 ][ 315 ],
   alphaCSR[ 190 ][ 316 ],
   alphaCSR[ 190 ][ 317 ],
   alphaCSR[ 190 ][ 318 ],
   alphaCSR[ 190 ][ 319 ],
   alphaCSR[ 190 ][ 320 ],
   alphaCSR[ 190 ][ 321 ],
   alphaCSR[ 190 ][ 322 ],
   alphaCSR[ 190 ][ 323 ],
   alphaCSR[ 190 ][ 324 ],
   alphaCSR[ 190 ][ 325 ],
   alphaCSR[ 190 ][ 326 ],
   alphaCSR[ 190 ][ 327 ],
   alphaCSR[ 190 ][ 328 ],
   alphaCSR[ 190 ][ 329 ],
   alphaCSR[ 190 ][ 330 ],
   alphaCSR[ 190 ][ 331 ],
   alphaCSR[ 190 ][ 332 ],
   alphaCSR[ 190 ][ 333 ],
   alphaCSR[ 190 ][ 334 ],
   alphaCSR[ 190 ][ 335 ],
   alphaCSR[ 190 ][ 336 ],
   alphaCSR[ 190 ][ 337 ],
   alphaCSR[ 190 ][ 338 ],
   alphaCSR[ 190 ][ 339 ],
   alphaCSR[ 190 ][ 340 ],
   alphaCSR[ 190 ][ 341 ],
   alphaCSR[ 190 ][ 342 ],
   alphaCSR[ 190 ][ 343 ],
   alphaCSR[ 190 ][ 344 ],
   alphaCSR[ 190 ][ 345 ],
   alphaCSR[ 190 ][ 346 ],
   alphaCSR[ 190 ][ 347 ],
   alphaCSR[ 190 ][ 348 ],
   alphaCSR[ 190 ][ 349 ],
   alphaCSR[ 190 ][ 350 ],
   alphaCSR[ 190 ][ 351 ],
   alphaCSR[ 190 ][ 352 ],
   alphaCSR[ 190 ][ 353 ],
   alphaCSR[ 190 ][ 354 ],
   alphaCSR[ 190 ][ 355 ],
   alphaCSR[ 190 ][ 356 ],
   alphaCSR[ 190 ][ 357 ],
   alphaCSR[ 190 ][ 358 ],
   alphaCSR[ 190 ][ 359 ],
   alphaCSR[ 190 ][ 360 ],
   alphaCSR[ 190 ][ 361 ],
   alphaCSR[ 190 ][ 362 ],
   alphaCSR[ 190 ][ 363 ],
   alphaCSR[ 190 ][ 364 ],
   alphaCSR[ 190 ][ 365 ],
   alphaCSR[ 190 ][ 366 ],
   alphaCSR[ 190 ][ 367 ],
   alphaCSR[ 190 ][ 368 ],
   alphaCSR[ 190 ][ 369 ],
   alphaCSR[ 190 ][ 370 ],
   alphaCSR[ 190 ][ 371 ],
   alphaCSR[ 190 ][ 372 ],
   alphaCSR[ 190 ][ 373 ],
   alphaCSR[ 190 ][ 374 ],
   alphaCSR[ 190 ][ 375 ],
   alphaCSR[ 190 ][ 376 ],
   alphaCSR[ 190 ][ 377 ],
   alphaCSR[ 190 ][ 378 ],
   alphaCSR[ 190 ][ 379 ],
   alphaCSR[ 190 ][ 380 ],
   alphaCSR[ 190 ][ 381 ],
   alphaCSR[ 190 ][ 382 ],
   alphaCSR[ 190 ][ 383 ],
   alphaCSR[ 191 ][ 0 ],
   alphaCSR[ 191 ][ 1 ],
   alphaCSR[ 191 ][ 2 ],
   alphaCSR[ 191 ][ 3 ],
   alphaCSR[ 191 ][ 4 ],
   alphaCSR[ 191 ][ 5 ],
   alphaCSR[ 191 ][ 6 ],
   alphaCSR[ 191 ][ 7 ],
   alphaCSR[ 191 ][ 8 ],
   alphaCSR[ 191 ][ 9 ],
   alphaCSR[ 191 ][ 10 ],
   alphaCSR[ 191 ][ 11 ],
   alphaCSR[ 191 ][ 12 ],
   alphaCSR[ 191 ][ 13 ],
   alphaCSR[ 191 ][ 14 ],
   alphaCSR[ 191 ][ 15 ],
   alphaCSR[ 191 ][ 16 ],
   alphaCSR[ 191 ][ 17 ],
   alphaCSR[ 191 ][ 18 ],
   alphaCSR[ 191 ][ 19 ],
   alphaCSR[ 191 ][ 20 ],
   alphaCSR[ 191 ][ 21 ],
   alphaCSR[ 191 ][ 22 ],
   alphaCSR[ 191 ][ 23 ],
   alphaCSR[ 191 ][ 24 ],
   alphaCSR[ 191 ][ 25 ],
   alphaCSR[ 191 ][ 26 ],
   alphaCSR[ 191 ][ 27 ],
   alphaCSR[ 191 ][ 28 ],
   alphaCSR[ 191 ][ 29 ],
   alphaCSR[ 191 ][ 30 ],
   alphaCSR[ 191 ][ 31 ],
   alphaCSR[ 191 ][ 32 ],
   alphaCSR[ 191 ][ 33 ],
   alphaCSR[ 191 ][ 34 ],
   alphaCSR[ 191 ][ 35 ],
   alphaCSR[ 191 ][ 36 ],
   alphaCSR[ 191 ][ 37 ],
   alphaCSR[ 191 ][ 38 ],
   alphaCSR[ 191 ][ 39 ],
   alphaCSR[ 191 ][ 40 ],
   alphaCSR[ 191 ][ 41 ],
   alphaCSR[ 191 ][ 42 ],
   alphaCSR[ 191 ][ 43 ],
   alphaCSR[ 191 ][ 44 ],
   alphaCSR[ 191 ][ 45 ],
   alphaCSR[ 191 ][ 46 ],
   alphaCSR[ 191 ][ 47 ],
   alphaCSR[ 191 ][ 48 ],
   alphaCSR[ 191 ][ 49 ],
   alphaCSR[ 191 ][ 50 ],
   alphaCSR[ 191 ][ 51 ],
   alphaCSR[ 191 ][ 52 ],
   alphaCSR[ 191 ][ 53 ],
   alphaCSR[ 191 ][ 54 ],
   alphaCSR[ 191 ][ 55 ],
   alphaCSR[ 191 ][ 56 ],
   alphaCSR[ 191 ][ 57 ],
   alphaCSR[ 191 ][ 58 ],
   alphaCSR[ 191 ][ 59 ],
   alphaCSR[ 191 ][ 60 ],
   alphaCSR[ 191 ][ 61 ],
   alphaCSR[ 191 ][ 62 ],
   alphaCSR[ 191 ][ 63 ],
   alphaCSR[ 191 ][ 64 ],
   alphaCSR[ 191 ][ 65 ],
   alphaCSR[ 191 ][ 66 ],
   alphaCSR[ 191 ][ 67 ],
   alphaCSR[ 191 ][ 68 ],
   alphaCSR[ 191 ][ 69 ],
   alphaCSR[ 191 ][ 70 ],
   alphaCSR[ 191 ][ 71 ],
   alphaCSR[ 191 ][ 72 ],
   alphaCSR[ 191 ][ 73 ],
   alphaCSR[ 191 ][ 74 ],
   alphaCSR[ 191 ][ 75 ],
   alphaCSR[ 191 ][ 76 ],
   alphaCSR[ 191 ][ 77 ],
   alphaCSR[ 191 ][ 78 ],
   alphaCSR[ 191 ][ 79 ],
   alphaCSR[ 191 ][ 80 ],
   alphaCSR[ 191 ][ 81 ],
   alphaCSR[ 191 ][ 82 ],
   alphaCSR[ 191 ][ 83 ],
   alphaCSR[ 191 ][ 84 ],
   alphaCSR[ 191 ][ 85 ],
   alphaCSR[ 191 ][ 86 ],
   alphaCSR[ 191 ][ 87 ],
   alphaCSR[ 191 ][ 88 ],
   alphaCSR[ 191 ][ 89 ],
   alphaCSR[ 191 ][ 90 ],
   alphaCSR[ 191 ][ 91 ],
   alphaCSR[ 191 ][ 92 ],
   alphaCSR[ 191 ][ 93 ],
   alphaCSR[ 191 ][ 94 ],
   alphaCSR[ 191 ][ 95 ],
   alphaCSR[ 191 ][ 96 ],
   alphaCSR[ 191 ][ 97 ],
   alphaCSR[ 191 ][ 98 ],
   alphaCSR[ 191 ][ 99 ],
   alphaCSR[ 191 ][ 100 ],
   alphaCSR[ 191 ][ 101 ],
   alphaCSR[ 191 ][ 102 ],
   alphaCSR[ 191 ][ 103 ],
   alphaCSR[ 191 ][ 104 ],
   alphaCSR[ 191 ][ 105 ],
   alphaCSR[ 191 ][ 106 ],
   alphaCSR[ 191 ][ 107 ],
   alphaCSR[ 191 ][ 108 ],
   alphaCSR[ 191 ][ 109 ],
   alphaCSR[ 191 ][ 110 ],
   alphaCSR[ 191 ][ 111 ],
   alphaCSR[ 191 ][ 112 ],
   alphaCSR[ 191 ][ 113 ],
   alphaCSR[ 191 ][ 114 ],
   alphaCSR[ 191 ][ 115 ],
   alphaCSR[ 191 ][ 116 ],
   alphaCSR[ 191 ][ 117 ],
   alphaCSR[ 191 ][ 118 ],
   alphaCSR[ 191 ][ 119 ],
   alphaCSR[ 191 ][ 120 ],
   alphaCSR[ 191 ][ 121 ],
   alphaCSR[ 191 ][ 122 ],
   alphaCSR[ 191 ][ 123 ],
   alphaCSR[ 191 ][ 124 ],
   alphaCSR[ 191 ][ 125 ],
   alphaCSR[ 191 ][ 126 ],
   alphaCSR[ 191 ][ 127 ],
   alphaCSR[ 191 ][ 128 ],
   alphaCSR[ 191 ][ 129 ],
   alphaCSR[ 191 ][ 130 ],
   alphaCSR[ 191 ][ 131 ],
   alphaCSR[ 191 ][ 132 ],
   alphaCSR[ 191 ][ 133 ],
   alphaCSR[ 191 ][ 134 ],
   alphaCSR[ 191 ][ 135 ],
   alphaCSR[ 191 ][ 136 ],
   alphaCSR[ 191 ][ 137 ],
   alphaCSR[ 191 ][ 138 ],
   alphaCSR[ 191 ][ 139 ],
   alphaCSR[ 191 ][ 140 ],
   alphaCSR[ 191 ][ 141 ],
   alphaCSR[ 191 ][ 142 ],
   alphaCSR[ 191 ][ 143 ],
   alphaCSR[ 191 ][ 144 ],
   alphaCSR[ 191 ][ 145 ],
   alphaCSR[ 191 ][ 146 ],
   alphaCSR[ 191 ][ 147 ],
   alphaCSR[ 191 ][ 148 ],
   alphaCSR[ 191 ][ 149 ],
   alphaCSR[ 191 ][ 150 ],
   alphaCSR[ 191 ][ 151 ],
   alphaCSR[ 191 ][ 152 ],
   alphaCSR[ 191 ][ 153 ],
   alphaCSR[ 191 ][ 154 ],
   alphaCSR[ 191 ][ 155 ],
   alphaCSR[ 191 ][ 156 ],
   alphaCSR[ 191 ][ 157 ],
   alphaCSR[ 191 ][ 158 ],
   alphaCSR[ 191 ][ 159 ],
   alphaCSR[ 191 ][ 160 ],
   alphaCSR[ 191 ][ 161 ],
   alphaCSR[ 191 ][ 162 ],
   alphaCSR[ 191 ][ 163 ],
   alphaCSR[ 191 ][ 164 ],
   alphaCSR[ 191 ][ 165 ],
   alphaCSR[ 191 ][ 166 ],
   alphaCSR[ 191 ][ 167 ],
   alphaCSR[ 191 ][ 168 ],
   alphaCSR[ 191 ][ 169 ],
   alphaCSR[ 191 ][ 170 ],
   alphaCSR[ 191 ][ 171 ],
   alphaCSR[ 191 ][ 172 ],
   alphaCSR[ 191 ][ 173 ],
   alphaCSR[ 191 ][ 174 ],
   alphaCSR[ 191 ][ 175 ],
   alphaCSR[ 191 ][ 176 ],
   alphaCSR[ 191 ][ 177 ],
   alphaCSR[ 191 ][ 178 ],
   alphaCSR[ 191 ][ 179 ],
   alphaCSR[ 191 ][ 180 ],
   alphaCSR[ 191 ][ 181 ],
   alphaCSR[ 191 ][ 182 ],
   alphaCSR[ 191 ][ 183 ],
   alphaCSR[ 191 ][ 184 ],
   alphaCSR[ 191 ][ 185 ],
   alphaCSR[ 191 ][ 186 ],
   alphaCSR[ 191 ][ 187 ],
   alphaCSR[ 191 ][ 188 ],
   alphaCSR[ 191 ][ 189 ],
   alphaCSR[ 191 ][ 190 ],
   alphaCSR[ 191 ][ 191 ],
   alphaCSR[ 191 ][ 192 ],
   alphaCSR[ 191 ][ 193 ],
   alphaCSR[ 191 ][ 194 ],
   alphaCSR[ 191 ][ 195 ],
   alphaCSR[ 191 ][ 196 ],
   alphaCSR[ 191 ][ 197 ],
   alphaCSR[ 191 ][ 198 ],
   alphaCSR[ 191 ][ 199 ],
   alphaCSR[ 191 ][ 200 ],
   alphaCSR[ 191 ][ 201 ],
   alphaCSR[ 191 ][ 202 ],
   alphaCSR[ 191 ][ 203 ],
   alphaCSR[ 191 ][ 204 ],
   alphaCSR[ 191 ][ 205 ],
   alphaCSR[ 191 ][ 206 ],
   alphaCSR[ 191 ][ 207 ],
   alphaCSR[ 191 ][ 208 ],
   alphaCSR[ 191 ][ 209 ],
   alphaCSR[ 191 ][ 210 ],
   alphaCSR[ 191 ][ 211 ],
   alphaCSR[ 191 ][ 212 ],
   alphaCSR[ 191 ][ 213 ],
   alphaCSR[ 191 ][ 214 ],
   alphaCSR[ 191 ][ 215 ],
   alphaCSR[ 191 ][ 216 ],
   alphaCSR[ 191 ][ 217 ],
   alphaCSR[ 191 ][ 218 ],
   alphaCSR[ 191 ][ 219 ],
   alphaCSR[ 191 ][ 220 ],
   alphaCSR[ 191 ][ 221 ],
   alphaCSR[ 191 ][ 222 ],
   alphaCSR[ 191 ][ 223 ],
   alphaCSR[ 191 ][ 224 ],
   alphaCSR[ 191 ][ 225 ],
   alphaCSR[ 191 ][ 226 ],
   alphaCSR[ 191 ][ 227 ],
   alphaCSR[ 191 ][ 228 ],
   alphaCSR[ 191 ][ 229 ],
   alphaCSR[ 191 ][ 230 ],
   alphaCSR[ 191 ][ 231 ],
   alphaCSR[ 191 ][ 232 ],
   alphaCSR[ 191 ][ 233 ],
   alphaCSR[ 191 ][ 234 ],
   alphaCSR[ 191 ][ 235 ],
   alphaCSR[ 191 ][ 236 ],
   alphaCSR[ 191 ][ 237 ],
   alphaCSR[ 191 ][ 238 ],
   alphaCSR[ 191 ][ 239 ],
   alphaCSR[ 191 ][ 240 ],
   alphaCSR[ 191 ][ 241 ],
   alphaCSR[ 191 ][ 242 ],
   alphaCSR[ 191 ][ 243 ],
   alphaCSR[ 191 ][ 244 ],
   alphaCSR[ 191 ][ 245 ],
   alphaCSR[ 191 ][ 246 ],
   alphaCSR[ 191 ][ 247 ],
   alphaCSR[ 191 ][ 248 ],
   alphaCSR[ 191 ][ 249 ],
   alphaCSR[ 191 ][ 250 ],
   alphaCSR[ 191 ][ 251 ],
   alphaCSR[ 191 ][ 252 ],
   alphaCSR[ 191 ][ 253 ],
   alphaCSR[ 191 ][ 254 ],
   alphaCSR[ 191 ][ 255 ],
   alphaCSR[ 191 ][ 256 ],
   alphaCSR[ 191 ][ 257 ],
   alphaCSR[ 191 ][ 258 ],
   alphaCSR[ 191 ][ 259 ],
   alphaCSR[ 191 ][ 260 ],
   alphaCSR[ 191 ][ 261 ],
   alphaCSR[ 191 ][ 262 ],
   alphaCSR[ 191 ][ 263 ],
   alphaCSR[ 191 ][ 264 ],
   alphaCSR[ 191 ][ 265 ],
   alphaCSR[ 191 ][ 266 ],
   alphaCSR[ 191 ][ 267 ],
   alphaCSR[ 191 ][ 268 ],
   alphaCSR[ 191 ][ 269 ],
   alphaCSR[ 191 ][ 270 ],
   alphaCSR[ 191 ][ 271 ],
   alphaCSR[ 191 ][ 272 ],
   alphaCSR[ 191 ][ 273 ],
   alphaCSR[ 191 ][ 274 ],
   alphaCSR[ 191 ][ 275 ],
   alphaCSR[ 191 ][ 276 ],
   alphaCSR[ 191 ][ 277 ],
   alphaCSR[ 191 ][ 278 ],
   alphaCSR[ 191 ][ 279 ],
   alphaCSR[ 191 ][ 280 ],
   alphaCSR[ 191 ][ 281 ],
   alphaCSR[ 191 ][ 282 ],
   alphaCSR[ 191 ][ 283 ],
   alphaCSR[ 191 ][ 284 ],
   alphaCSR[ 191 ][ 285 ],
   alphaCSR[ 191 ][ 286 ],
   alphaCSR[ 191 ][ 287 ],
   alphaCSR[ 191 ][ 288 ],
   alphaCSR[ 191 ][ 289 ],
   alphaCSR[ 191 ][ 290 ],
   alphaCSR[ 191 ][ 291 ],
   alphaCSR[ 191 ][ 292 ],
   alphaCSR[ 191 ][ 293 ],
   alphaCSR[ 191 ][ 294 ],
   alphaCSR[ 191 ][ 295 ],
   alphaCSR[ 191 ][ 296 ],
   alphaCSR[ 191 ][ 297 ],
   alphaCSR[ 191 ][ 298 ],
   alphaCSR[ 191 ][ 299 ],
   alphaCSR[ 191 ][ 300 ],
   alphaCSR[ 191 ][ 301 ],
   alphaCSR[ 191 ][ 302 ],
   alphaCSR[ 191 ][ 303 ],
   alphaCSR[ 191 ][ 304 ],
   alphaCSR[ 191 ][ 305 ],
   alphaCSR[ 191 ][ 306 ],
   alphaCSR[ 191 ][ 307 ],
   alphaCSR[ 191 ][ 308 ],
   alphaCSR[ 191 ][ 309 ],
   alphaCSR[ 191 ][ 310 ],
   alphaCSR[ 191 ][ 311 ],
   alphaCSR[ 191 ][ 312 ],
   alphaCSR[ 191 ][ 313 ],
   alphaCSR[ 191 ][ 314 ],
   alphaCSR[ 191 ][ 315 ],
   alphaCSR[ 191 ][ 316 ],
   alphaCSR[ 191 ][ 317 ],
   alphaCSR[ 191 ][ 318 ],
   alphaCSR[ 191 ][ 319 ],
   alphaCSR[ 191 ][ 320 ],
   alphaCSR[ 191 ][ 321 ],
   alphaCSR[ 191 ][ 322 ],
   alphaCSR[ 191 ][ 323 ],
   alphaCSR[ 191 ][ 324 ],
   alphaCSR[ 191 ][ 325 ],
   alphaCSR[ 191 ][ 326 ],
   alphaCSR[ 191 ][ 327 ],
   alphaCSR[ 191 ][ 328 ],
   alphaCSR[ 191 ][ 329 ],
   alphaCSR[ 191 ][ 330 ],
   alphaCSR[ 191 ][ 331 ],
   alphaCSR[ 191 ][ 332 ],
   alphaCSR[ 191 ][ 333 ],
   alphaCSR[ 191 ][ 334 ],
   alphaCSR[ 191 ][ 335 ],
   alphaCSR[ 191 ][ 336 ],
   alphaCSR[ 191 ][ 337 ],
   alphaCSR[ 191 ][ 338 ],
   alphaCSR[ 191 ][ 339 ],
   alphaCSR[ 191 ][ 340 ],
   alphaCSR[ 191 ][ 341 ],
   alphaCSR[ 191 ][ 342 ],
   alphaCSR[ 191 ][ 343 ],
   alphaCSR[ 191 ][ 344 ],
   alphaCSR[ 191 ][ 345 ],
   alphaCSR[ 191 ][ 346 ],
   alphaCSR[ 191 ][ 347 ],
   alphaCSR[ 191 ][ 348 ],
   alphaCSR[ 191 ][ 349 ],
   alphaCSR[ 191 ][ 350 ],
   alphaCSR[ 191 ][ 351 ],
   alphaCSR[ 191 ][ 352 ],
   alphaCSR[ 191 ][ 353 ],
   alphaCSR[ 191 ][ 354 ],
   alphaCSR[ 191 ][ 355 ],
   alphaCSR[ 191 ][ 356 ],
   alphaCSR[ 191 ][ 357 ],
   alphaCSR[ 191 ][ 358 ],
   alphaCSR[ 191 ][ 359 ],
   alphaCSR[ 191 ][ 360 ],
   alphaCSR[ 191 ][ 361 ],
   alphaCSR[ 191 ][ 362 ],
   alphaCSR[ 191 ][ 363 ],
   alphaCSR[ 191 ][ 364 ],
   alphaCSR[ 191 ][ 365 ],
   alphaCSR[ 191 ][ 366 ],
   alphaCSR[ 191 ][ 367 ],
   alphaCSR[ 191 ][ 368 ],
   alphaCSR[ 191 ][ 369 ],
   alphaCSR[ 191 ][ 370 ],
   alphaCSR[ 191 ][ 371 ],
   alphaCSR[ 191 ][ 372 ],
   alphaCSR[ 191 ][ 373 ],
   alphaCSR[ 191 ][ 374 ],
   alphaCSR[ 191 ][ 375 ],
   alphaCSR[ 191 ][ 376 ],
   alphaCSR[ 191 ][ 377 ],
   alphaCSR[ 191 ][ 378 ],
   alphaCSR[ 191 ][ 379 ],
   alphaCSR[ 191 ][ 380 ],
   alphaCSR[ 191 ][ 381 ],
   alphaCSR[ 191 ][ 382 ],
   alphaCSR[ 191 ][ 383 ],
   alphaCSR[ 192 ][ 0 ],
   alphaCSR[ 192 ][ 1 ],
   alphaCSR[ 192 ][ 2 ],
   alphaCSR[ 192 ][ 3 ],
   alphaCSR[ 192 ][ 4 ],
   alphaCSR[ 192 ][ 5 ],
   alphaCSR[ 192 ][ 6 ],
   alphaCSR[ 192 ][ 7 ],
   alphaCSR[ 192 ][ 8 ],
   alphaCSR[ 192 ][ 9 ],
   alphaCSR[ 192 ][ 10 ],
   alphaCSR[ 192 ][ 11 ],
   alphaCSR[ 192 ][ 12 ],
   alphaCSR[ 192 ][ 13 ],
   alphaCSR[ 192 ][ 14 ],
   alphaCSR[ 192 ][ 15 ],
   alphaCSR[ 192 ][ 16 ],
   alphaCSR[ 192 ][ 17 ],
   alphaCSR[ 192 ][ 18 ],
   alphaCSR[ 192 ][ 19 ],
   alphaCSR[ 192 ][ 20 ],
   alphaCSR[ 192 ][ 21 ],
   alphaCSR[ 192 ][ 22 ],
   alphaCSR[ 192 ][ 23 ],
   alphaCSR[ 192 ][ 24 ],
   alphaCSR[ 192 ][ 25 ],
   alphaCSR[ 192 ][ 26 ],
   alphaCSR[ 192 ][ 27 ],
   alphaCSR[ 192 ][ 28 ],
   alphaCSR[ 192 ][ 29 ],
   alphaCSR[ 192 ][ 30 ],
   alphaCSR[ 192 ][ 31 ],
   alphaCSR[ 192 ][ 32 ],
   alphaCSR[ 192 ][ 33 ],
   alphaCSR[ 192 ][ 34 ],
   alphaCSR[ 192 ][ 35 ],
   alphaCSR[ 192 ][ 36 ],
   alphaCSR[ 192 ][ 37 ],
   alphaCSR[ 192 ][ 38 ],
   alphaCSR[ 192 ][ 39 ],
   alphaCSR[ 192 ][ 40 ],
   alphaCSR[ 192 ][ 41 ],
   alphaCSR[ 192 ][ 42 ],
   alphaCSR[ 192 ][ 43 ],
   alphaCSR[ 192 ][ 44 ],
   alphaCSR[ 192 ][ 45 ],
   alphaCSR[ 192 ][ 46 ],
   alphaCSR[ 192 ][ 47 ],
   alphaCSR[ 192 ][ 48 ],
   alphaCSR[ 192 ][ 49 ],
   alphaCSR[ 192 ][ 50 ],
   alphaCSR[ 192 ][ 51 ],
   alphaCSR[ 192 ][ 52 ],
   alphaCSR[ 192 ][ 53 ],
   alphaCSR[ 192 ][ 54 ],
   alphaCSR[ 192 ][ 55 ],
   alphaCSR[ 192 ][ 56 ],
   alphaCSR[ 192 ][ 57 ],
   alphaCSR[ 192 ][ 58 ],
   alphaCSR[ 192 ][ 59 ],
   alphaCSR[ 192 ][ 60 ],
   alphaCSR[ 192 ][ 61 ],
   alphaCSR[ 192 ][ 62 ],
   alphaCSR[ 192 ][ 63 ],
   alphaCSR[ 192 ][ 64 ],
   alphaCSR[ 192 ][ 65 ],
   alphaCSR[ 192 ][ 66 ],
   alphaCSR[ 192 ][ 67 ],
   alphaCSR[ 192 ][ 68 ],
   alphaCSR[ 192 ][ 69 ],
   alphaCSR[ 192 ][ 70 ],
   alphaCSR[ 192 ][ 71 ],
   alphaCSR[ 192 ][ 72 ],
   alphaCSR[ 192 ][ 73 ],
   alphaCSR[ 192 ][ 74 ],
   alphaCSR[ 192 ][ 75 ],
   alphaCSR[ 192 ][ 76 ],
   alphaCSR[ 192 ][ 77 ],
   alphaCSR[ 192 ][ 78 ],
   alphaCSR[ 192 ][ 79 ],
   alphaCSR[ 192 ][ 80 ],
   alphaCSR[ 192 ][ 81 ],
   alphaCSR[ 192 ][ 82 ],
   alphaCSR[ 192 ][ 83 ],
   alphaCSR[ 192 ][ 84 ],
   alphaCSR[ 192 ][ 85 ],
   alphaCSR[ 192 ][ 86 ],
   alphaCSR[ 192 ][ 87 ],
   alphaCSR[ 192 ][ 88 ],
   alphaCSR[ 192 ][ 89 ],
   alphaCSR[ 192 ][ 90 ],
   alphaCSR[ 192 ][ 91 ],
   alphaCSR[ 192 ][ 92 ],
   alphaCSR[ 192 ][ 93 ],
   alphaCSR[ 192 ][ 94 ],
   alphaCSR[ 192 ][ 95 ],
   alphaCSR[ 192 ][ 96 ],
   alphaCSR[ 192 ][ 97 ],
   alphaCSR[ 192 ][ 98 ],
   alphaCSR[ 192 ][ 99 ],
   alphaCSR[ 192 ][ 100 ],
   alphaCSR[ 192 ][ 101 ],
   alphaCSR[ 192 ][ 102 ],
   alphaCSR[ 192 ][ 103 ],
   alphaCSR[ 192 ][ 104 ],
   alphaCSR[ 192 ][ 105 ],
   alphaCSR[ 192 ][ 106 ],
   alphaCSR[ 192 ][ 107 ],
   alphaCSR[ 192 ][ 108 ],
   alphaCSR[ 192 ][ 109 ],
   alphaCSR[ 192 ][ 110 ],
   alphaCSR[ 192 ][ 111 ],
   alphaCSR[ 192 ][ 112 ],
   alphaCSR[ 192 ][ 113 ],
   alphaCSR[ 192 ][ 114 ],
   alphaCSR[ 192 ][ 115 ],
   alphaCSR[ 192 ][ 116 ],
   alphaCSR[ 192 ][ 117 ],
   alphaCSR[ 192 ][ 118 ],
   alphaCSR[ 192 ][ 119 ],
   alphaCSR[ 192 ][ 120 ],
   alphaCSR[ 192 ][ 121 ],
   alphaCSR[ 192 ][ 122 ],
   alphaCSR[ 192 ][ 123 ],
   alphaCSR[ 192 ][ 124 ],
   alphaCSR[ 192 ][ 125 ],
   alphaCSR[ 192 ][ 126 ],
   alphaCSR[ 192 ][ 127 ],
   alphaCSR[ 192 ][ 128 ],
   alphaCSR[ 192 ][ 129 ],
   alphaCSR[ 192 ][ 130 ],
   alphaCSR[ 192 ][ 131 ],
   alphaCSR[ 192 ][ 132 ],
   alphaCSR[ 192 ][ 133 ],
   alphaCSR[ 192 ][ 134 ],
   alphaCSR[ 192 ][ 135 ],
   alphaCSR[ 192 ][ 136 ],
   alphaCSR[ 192 ][ 137 ],
   alphaCSR[ 192 ][ 138 ],
   alphaCSR[ 192 ][ 139 ],
   alphaCSR[ 192 ][ 140 ],
   alphaCSR[ 192 ][ 141 ],
   alphaCSR[ 192 ][ 142 ],
   alphaCSR[ 192 ][ 143 ],
   alphaCSR[ 192 ][ 144 ],
   alphaCSR[ 192 ][ 145 ],
   alphaCSR[ 192 ][ 146 ],
   alphaCSR[ 192 ][ 147 ],
   alphaCSR[ 192 ][ 148 ],
   alphaCSR[ 192 ][ 149 ],
   alphaCSR[ 192 ][ 150 ],
   alphaCSR[ 192 ][ 151 ],
   alphaCSR[ 192 ][ 152 ],
   alphaCSR[ 192 ][ 153 ],
   alphaCSR[ 192 ][ 154 ],
   alphaCSR[ 192 ][ 155 ],
   alphaCSR[ 192 ][ 156 ],
   alphaCSR[ 192 ][ 157 ],
   alphaCSR[ 192 ][ 158 ],
   alphaCSR[ 192 ][ 159 ],
   alphaCSR[ 192 ][ 160 ],
   alphaCSR[ 192 ][ 161 ],
   alphaCSR[ 192 ][ 162 ],
   alphaCSR[ 192 ][ 163 ],
   alphaCSR[ 192 ][ 164 ],
   alphaCSR[ 192 ][ 165 ],
   alphaCSR[ 192 ][ 166 ],
   alphaCSR[ 192 ][ 167 ],
   alphaCSR[ 192 ][ 168 ],
   alphaCSR[ 192 ][ 169 ],
   alphaCSR[ 192 ][ 170 ],
   alphaCSR[ 192 ][ 171 ],
   alphaCSR[ 192 ][ 172 ],
   alphaCSR[ 192 ][ 173 ],
   alphaCSR[ 192 ][ 174 ],
   alphaCSR[ 192 ][ 175 ],
   alphaCSR[ 192 ][ 176 ],
   alphaCSR[ 192 ][ 177 ],
   alphaCSR[ 192 ][ 178 ],
   alphaCSR[ 192 ][ 179 ],
   alphaCSR[ 192 ][ 180 ],
   alphaCSR[ 192 ][ 181 ],
   alphaCSR[ 192 ][ 182 ],
   alphaCSR[ 192 ][ 183 ],
   alphaCSR[ 192 ][ 184 ],
   alphaCSR[ 192 ][ 185 ],
   alphaCSR[ 192 ][ 186 ],
   alphaCSR[ 192 ][ 187 ],
   alphaCSR[ 192 ][ 188 ],
   alphaCSR[ 192 ][ 189 ],
   alphaCSR[ 192 ][ 190 ],
   alphaCSR[ 192 ][ 191 ],
   alphaCSR[ 192 ][ 192 ],
   alphaCSR[ 192 ][ 193 ],
   alphaCSR[ 192 ][ 194 ],
   alphaCSR[ 192 ][ 195 ],
   alphaCSR[ 192 ][ 196 ],
   alphaCSR[ 192 ][ 197 ],
   alphaCSR[ 192 ][ 198 ],
   alphaCSR[ 192 ][ 199 ],
   alphaCSR[ 192 ][ 200 ],
   alphaCSR[ 192 ][ 201 ],
   alphaCSR[ 192 ][ 202 ],
   alphaCSR[ 192 ][ 203 ],
   alphaCSR[ 192 ][ 204 ],
   alphaCSR[ 192 ][ 205 ],
   alphaCSR[ 192 ][ 206 ],
   alphaCSR[ 192 ][ 207 ],
   alphaCSR[ 192 ][ 208 ],
   alphaCSR[ 192 ][ 209 ],
   alphaCSR[ 192 ][ 210 ],
   alphaCSR[ 192 ][ 211 ],
   alphaCSR[ 192 ][ 212 ],
   alphaCSR[ 192 ][ 213 ],
   alphaCSR[ 192 ][ 214 ],
   alphaCSR[ 192 ][ 215 ],
   alphaCSR[ 192 ][ 216 ],
   alphaCSR[ 192 ][ 217 ],
   alphaCSR[ 192 ][ 218 ],
   alphaCSR[ 192 ][ 219 ],
   alphaCSR[ 192 ][ 220 ],
   alphaCSR[ 192 ][ 221 ],
   alphaCSR[ 192 ][ 222 ],
   alphaCSR[ 192 ][ 223 ],
   alphaCSR[ 192 ][ 224 ],
   alphaCSR[ 192 ][ 225 ],
   alphaCSR[ 192 ][ 226 ],
   alphaCSR[ 192 ][ 227 ],
   alphaCSR[ 192 ][ 228 ],
   alphaCSR[ 192 ][ 229 ],
   alphaCSR[ 192 ][ 230 ],
   alphaCSR[ 192 ][ 231 ],
   alphaCSR[ 192 ][ 232 ],
   alphaCSR[ 192 ][ 233 ],
   alphaCSR[ 192 ][ 234 ],
   alphaCSR[ 192 ][ 235 ],
   alphaCSR[ 192 ][ 236 ],
   alphaCSR[ 192 ][ 237 ],
   alphaCSR[ 192 ][ 238 ],
   alphaCSR[ 192 ][ 239 ],
   alphaCSR[ 192 ][ 240 ],
   alphaCSR[ 192 ][ 241 ],
   alphaCSR[ 192 ][ 242 ],
   alphaCSR[ 192 ][ 243 ],
   alphaCSR[ 192 ][ 244 ],
   alphaCSR[ 192 ][ 245 ],
   alphaCSR[ 192 ][ 246 ],
   alphaCSR[ 192 ][ 247 ],
   alphaCSR[ 192 ][ 248 ],
   alphaCSR[ 192 ][ 249 ],
   alphaCSR[ 192 ][ 250 ],
   alphaCSR[ 192 ][ 251 ],
   alphaCSR[ 192 ][ 252 ],
   alphaCSR[ 192 ][ 253 ],
   alphaCSR[ 192 ][ 254 ],
   alphaCSR[ 192 ][ 255 ],
   alphaCSR[ 192 ][ 256 ],
   alphaCSR[ 192 ][ 257 ],
   alphaCSR[ 192 ][ 258 ],
   alphaCSR[ 192 ][ 259 ],
   alphaCSR[ 192 ][ 260 ],
   alphaCSR[ 192 ][ 261 ],
   alphaCSR[ 192 ][ 262 ],
   alphaCSR[ 192 ][ 263 ],
   alphaCSR[ 192 ][ 264 ],
   alphaCSR[ 192 ][ 265 ],
   alphaCSR[ 192 ][ 266 ],
   alphaCSR[ 192 ][ 267 ],
   alphaCSR[ 192 ][ 268 ],
   alphaCSR[ 192 ][ 269 ],
   alphaCSR[ 192 ][ 270 ],
   alphaCSR[ 192 ][ 271 ],
   alphaCSR[ 192 ][ 272 ],
   alphaCSR[ 192 ][ 273 ],
   alphaCSR[ 192 ][ 274 ],
   alphaCSR[ 192 ][ 275 ],
   alphaCSR[ 192 ][ 276 ],
   alphaCSR[ 192 ][ 277 ],
   alphaCSR[ 192 ][ 278 ],
   alphaCSR[ 192 ][ 279 ],
   alphaCSR[ 192 ][ 280 ],
   alphaCSR[ 192 ][ 281 ],
   alphaCSR[ 192 ][ 282 ],
   alphaCSR[ 192 ][ 283 ],
   alphaCSR[ 192 ][ 284 ],
   alphaCSR[ 192 ][ 285 ],
   alphaCSR[ 192 ][ 286 ],
   alphaCSR[ 192 ][ 287 ],
   alphaCSR[ 192 ][ 288 ],
   alphaCSR[ 192 ][ 289 ],
   alphaCSR[ 192 ][ 290 ],
   alphaCSR[ 192 ][ 291 ],
   alphaCSR[ 192 ][ 292 ],
   alphaCSR[ 192 ][ 293 ],
   alphaCSR[ 192 ][ 294 ],
   alphaCSR[ 192 ][ 295 ],
   alphaCSR[ 192 ][ 296 ],
   alphaCSR[ 192 ][ 297 ],
   alphaCSR[ 192 ][ 298 ],
   alphaCSR[ 192 ][ 299 ],
   alphaCSR[ 192 ][ 300 ],
   alphaCSR[ 192 ][ 301 ],
   alphaCSR[ 192 ][ 302 ],
   alphaCSR[ 192 ][ 303 ],
   alphaCSR[ 192 ][ 304 ],
   alphaCSR[ 192 ][ 305 ],
   alphaCSR[ 192 ][ 306 ],
   alphaCSR[ 192 ][ 307 ],
   alphaCSR[ 192 ][ 308 ],
   alphaCSR[ 192 ][ 309 ],
   alphaCSR[ 192 ][ 310 ],
   alphaCSR[ 192 ][ 311 ],
   alphaCSR[ 192 ][ 312 ],
   alphaCSR[ 192 ][ 313 ],
   alphaCSR[ 192 ][ 314 ],
   alphaCSR[ 192 ][ 315 ],
   alphaCSR[ 192 ][ 316 ],
   alphaCSR[ 192 ][ 317 ],
   alphaCSR[ 192 ][ 318 ],
   alphaCSR[ 192 ][ 319 ],
   alphaCSR[ 192 ][ 320 ],
   alphaCSR[ 192 ][ 321 ],
   alphaCSR[ 192 ][ 322 ],
   alphaCSR[ 192 ][ 323 ],
   alphaCSR[ 192 ][ 324 ],
   alphaCSR[ 192 ][ 325 ],
   alphaCSR[ 192 ][ 326 ],
   alphaCSR[ 192 ][ 327 ],
   alphaCSR[ 192 ][ 328 ],
   alphaCSR[ 192 ][ 329 ],
   alphaCSR[ 192 ][ 330 ],
   alphaCSR[ 192 ][ 331 ],
   alphaCSR[ 192 ][ 332 ],
   alphaCSR[ 192 ][ 333 ],
   alphaCSR[ 192 ][ 334 ],
   alphaCSR[ 192 ][ 335 ],
   alphaCSR[ 192 ][ 336 ],
   alphaCSR[ 192 ][ 337 ],
   alphaCSR[ 192 ][ 338 ],
   alphaCSR[ 192 ][ 339 ],
   alphaCSR[ 192 ][ 340 ],
   alphaCSR[ 192 ][ 341 ],
   alphaCSR[ 192 ][ 342 ],
   alphaCSR[ 192 ][ 343 ],
   alphaCSR[ 192 ][ 344 ],
   alphaCSR[ 192 ][ 345 ],
   alphaCSR[ 192 ][ 346 ],
   alphaCSR[ 192 ][ 347 ],
   alphaCSR[ 192 ][ 348 ],
   alphaCSR[ 192 ][ 349 ],
   alphaCSR[ 192 ][ 350 ],
   alphaCSR[ 192 ][ 351 ],
   alphaCSR[ 192 ][ 352 ],
   alphaCSR[ 192 ][ 353 ],
   alphaCSR[ 192 ][ 354 ],
   alphaCSR[ 192 ][ 355 ],
   alphaCSR[ 192 ][ 356 ],
   alphaCSR[ 192 ][ 357 ],
   alphaCSR[ 192 ][ 358 ],
   alphaCSR[ 192 ][ 359 ],
   alphaCSR[ 192 ][ 360 ],
   alphaCSR[ 192 ][ 361 ],
   alphaCSR[ 192 ][ 362 ],
   alphaCSR[ 192 ][ 363 ],
   alphaCSR[ 192 ][ 364 ],
   alphaCSR[ 192 ][ 365 ],
   alphaCSR[ 192 ][ 366 ],
   alphaCSR[ 192 ][ 367 ],
   alphaCSR[ 192 ][ 368 ],
   alphaCSR[ 192 ][ 369 ],
   alphaCSR[ 192 ][ 370 ],
   alphaCSR[ 192 ][ 371 ],
   alphaCSR[ 192 ][ 372 ],
   alphaCSR[ 192 ][ 373 ],
   alphaCSR[ 192 ][ 374 ],
   alphaCSR[ 192 ][ 375 ],
   alphaCSR[ 192 ][ 376 ],
   alphaCSR[ 192 ][ 377 ],
   alphaCSR[ 192 ][ 378 ],
   alphaCSR[ 192 ][ 379 ],
   alphaCSR[ 192 ][ 380 ],
   alphaCSR[ 192 ][ 381 ],
   alphaCSR[ 192 ][ 382 ],
   alphaCSR[ 192 ][ 383 ],
   alphaCSR[ 193 ][ 0 ],
   alphaCSR[ 193 ][ 1 ],
   alphaCSR[ 193 ][ 2 ],
   alphaCSR[ 193 ][ 3 ],
   alphaCSR[ 193 ][ 4 ],
   alphaCSR[ 193 ][ 5 ],
   alphaCSR[ 193 ][ 6 ],
   alphaCSR[ 193 ][ 7 ],
   alphaCSR[ 193 ][ 8 ],
   alphaCSR[ 193 ][ 9 ],
   alphaCSR[ 193 ][ 10 ],
   alphaCSR[ 193 ][ 11 ],
   alphaCSR[ 193 ][ 12 ],
   alphaCSR[ 193 ][ 13 ],
   alphaCSR[ 193 ][ 14 ],
   alphaCSR[ 193 ][ 15 ],
   alphaCSR[ 193 ][ 16 ],
   alphaCSR[ 193 ][ 17 ],
   alphaCSR[ 193 ][ 18 ],
   alphaCSR[ 193 ][ 19 ],
   alphaCSR[ 193 ][ 20 ],
   alphaCSR[ 193 ][ 21 ],
   alphaCSR[ 193 ][ 22 ],
   alphaCSR[ 193 ][ 23 ],
   alphaCSR[ 193 ][ 24 ],
   alphaCSR[ 193 ][ 25 ],
   alphaCSR[ 193 ][ 26 ],
   alphaCSR[ 193 ][ 27 ],
   alphaCSR[ 193 ][ 28 ],
   alphaCSR[ 193 ][ 29 ],
   alphaCSR[ 193 ][ 30 ],
   alphaCSR[ 193 ][ 31 ],
   alphaCSR[ 193 ][ 32 ],
   alphaCSR[ 193 ][ 33 ],
   alphaCSR[ 193 ][ 34 ],
   alphaCSR[ 193 ][ 35 ],
   alphaCSR[ 193 ][ 36 ],
   alphaCSR[ 193 ][ 37 ],
   alphaCSR[ 193 ][ 38 ],
   alphaCSR[ 193 ][ 39 ],
   alphaCSR[ 193 ][ 40 ],
   alphaCSR[ 193 ][ 41 ],
   alphaCSR[ 193 ][ 42 ],
   alphaCSR[ 193 ][ 43 ],
   alphaCSR[ 193 ][ 44 ],
   alphaCSR[ 193 ][ 45 ],
   alphaCSR[ 193 ][ 46 ],
   alphaCSR[ 193 ][ 47 ],
   alphaCSR[ 193 ][ 48 ],
   alphaCSR[ 193 ][ 49 ],
   alphaCSR[ 193 ][ 50 ],
   alphaCSR[ 193 ][ 51 ],
   alphaCSR[ 193 ][ 52 ],
   alphaCSR[ 193 ][ 53 ],
   alphaCSR[ 193 ][ 54 ],
   alphaCSR[ 193 ][ 55 ],
   alphaCSR[ 193 ][ 56 ],
   alphaCSR[ 193 ][ 57 ],
   alphaCSR[ 193 ][ 58 ],
   alphaCSR[ 193 ][ 59 ],
   alphaCSR[ 193 ][ 60 ],
   alphaCSR[ 193 ][ 61 ],
   alphaCSR[ 193 ][ 62 ],
   alphaCSR[ 193 ][ 63 ],
   alphaCSR[ 193 ][ 64 ],
   alphaCSR[ 193 ][ 65 ],
   alphaCSR[ 193 ][ 66 ],
   alphaCSR[ 193 ][ 67 ],
   alphaCSR[ 193 ][ 68 ],
   alphaCSR[ 193 ][ 69 ],
   alphaCSR[ 193 ][ 70 ],
   alphaCSR[ 193 ][ 71 ],
   alphaCSR[ 193 ][ 72 ],
   alphaCSR[ 193 ][ 73 ],
   alphaCSR[ 193 ][ 74 ],
   alphaCSR[ 193 ][ 75 ],
   alphaCSR[ 193 ][ 76 ],
   alphaCSR[ 193 ][ 77 ],
   alphaCSR[ 193 ][ 78 ],
   alphaCSR[ 193 ][ 79 ],
   alphaCSR[ 193 ][ 80 ],
   alphaCSR[ 193 ][ 81 ],
   alphaCSR[ 193 ][ 82 ],
   alphaCSR[ 193 ][ 83 ],
   alphaCSR[ 193 ][ 84 ],
   alphaCSR[ 193 ][ 85 ],
   alphaCSR[ 193 ][ 86 ],
   alphaCSR[ 193 ][ 87 ],
   alphaCSR[ 193 ][ 88 ],
   alphaCSR[ 193 ][ 89 ],
   alphaCSR[ 193 ][ 90 ],
   alphaCSR[ 193 ][ 91 ],
   alphaCSR[ 193 ][ 92 ],
   alphaCSR[ 193 ][ 93 ],
   alphaCSR[ 193 ][ 94 ],
   alphaCSR[ 193 ][ 95 ],
   alphaCSR[ 193 ][ 96 ],
   alphaCSR[ 193 ][ 97 ],
   alphaCSR[ 193 ][ 98 ],
   alphaCSR[ 193 ][ 99 ],
   alphaCSR[ 193 ][ 100 ],
   alphaCSR[ 193 ][ 101 ],
   alphaCSR[ 193 ][ 102 ],
   alphaCSR[ 193 ][ 103 ],
   alphaCSR[ 193 ][ 104 ],
   alphaCSR[ 193 ][ 105 ],
   alphaCSR[ 193 ][ 106 ],
   alphaCSR[ 193 ][ 107 ],
   alphaCSR[ 193 ][ 108 ],
   alphaCSR[ 193 ][ 109 ],
   alphaCSR[ 193 ][ 110 ],
   alphaCSR[ 193 ][ 111 ],
   alphaCSR[ 193 ][ 112 ],
   alphaCSR[ 193 ][ 113 ],
   alphaCSR[ 193 ][ 114 ],
   alphaCSR[ 193 ][ 115 ],
   alphaCSR[ 193 ][ 116 ],
   alphaCSR[ 193 ][ 117 ],
   alphaCSR[ 193 ][ 118 ],
   alphaCSR[ 193 ][ 119 ],
   alphaCSR[ 193 ][ 120 ],
   alphaCSR[ 193 ][ 121 ],
   alphaCSR[ 193 ][ 122 ],
   alphaCSR[ 193 ][ 123 ],
   alphaCSR[ 193 ][ 124 ],
   alphaCSR[ 193 ][ 125 ],
   alphaCSR[ 193 ][ 126 ],
   alphaCSR[ 193 ][ 127 ],
   alphaCSR[ 193 ][ 128 ],
   alphaCSR[ 193 ][ 129 ],
   alphaCSR[ 193 ][ 130 ],
   alphaCSR[ 193 ][ 131 ],
   alphaCSR[ 193 ][ 132 ],
   alphaCSR[ 193 ][ 133 ],
   alphaCSR[ 193 ][ 134 ],
   alphaCSR[ 193 ][ 135 ],
   alphaCSR[ 193 ][ 136 ],
   alphaCSR[ 193 ][ 137 ],
   alphaCSR[ 193 ][ 138 ],
   alphaCSR[ 193 ][ 139 ],
   alphaCSR[ 193 ][ 140 ],
   alphaCSR[ 193 ][ 141 ],
   alphaCSR[ 193 ][ 142 ],
   alphaCSR[ 193 ][ 143 ],
   alphaCSR[ 193 ][ 144 ],
   alphaCSR[ 193 ][ 145 ],
   alphaCSR[ 193 ][ 146 ],
   alphaCSR[ 193 ][ 147 ],
   alphaCSR[ 193 ][ 148 ],
   alphaCSR[ 193 ][ 149 ],
   alphaCSR[ 193 ][ 150 ],
   alphaCSR[ 193 ][ 151 ],
   alphaCSR[ 193 ][ 152 ],
   alphaCSR[ 193 ][ 153 ],
   alphaCSR[ 193 ][ 154 ],
   alphaCSR[ 193 ][ 155 ],
   alphaCSR[ 193 ][ 156 ],
   alphaCSR[ 193 ][ 157 ],
   alphaCSR[ 193 ][ 158 ],
   alphaCSR[ 193 ][ 159 ],
   alphaCSR[ 193 ][ 160 ],
   alphaCSR[ 193 ][ 161 ],
   alphaCSR[ 193 ][ 162 ],
   alphaCSR[ 193 ][ 163 ],
   alphaCSR[ 193 ][ 164 ],
   alphaCSR[ 193 ][ 165 ],
   alphaCSR[ 193 ][ 166 ],
   alphaCSR[ 193 ][ 167 ],
   alphaCSR[ 193 ][ 168 ],
   alphaCSR[ 193 ][ 169 ],
   alphaCSR[ 193 ][ 170 ],
   alphaCSR[ 193 ][ 171 ],
   alphaCSR[ 193 ][ 172 ],
   alphaCSR[ 193 ][ 173 ],
   alphaCSR[ 193 ][ 174 ],
   alphaCSR[ 193 ][ 175 ],
   alphaCSR[ 193 ][ 176 ],
   alphaCSR[ 193 ][ 177 ],
   alphaCSR[ 193 ][ 178 ],
   alphaCSR[ 193 ][ 179 ],
   alphaCSR[ 193 ][ 180 ],
   alphaCSR[ 193 ][ 181 ],
   alphaCSR[ 193 ][ 182 ],
   alphaCSR[ 193 ][ 183 ],
   alphaCSR[ 193 ][ 184 ],
   alphaCSR[ 193 ][ 185 ],
   alphaCSR[ 193 ][ 186 ],
   alphaCSR[ 193 ][ 187 ],
   alphaCSR[ 193 ][ 188 ],
   alphaCSR[ 193 ][ 189 ],
   alphaCSR[ 193 ][ 190 ],
   alphaCSR[ 193 ][ 191 ],
   alphaCSR[ 193 ][ 192 ],
   alphaCSR[ 193 ][ 193 ],
   alphaCSR[ 193 ][ 194 ],
   alphaCSR[ 193 ][ 195 ],
   alphaCSR[ 193 ][ 196 ],
   alphaCSR[ 193 ][ 197 ],
   alphaCSR[ 193 ][ 198 ],
   alphaCSR[ 193 ][ 199 ],
   alphaCSR[ 193 ][ 200 ],
   alphaCSR[ 193 ][ 201 ],
   alphaCSR[ 193 ][ 202 ],
   alphaCSR[ 193 ][ 203 ],
   alphaCSR[ 193 ][ 204 ],
   alphaCSR[ 193 ][ 205 ],
   alphaCSR[ 193 ][ 206 ],
   alphaCSR[ 193 ][ 207 ],
   alphaCSR[ 193 ][ 208 ],
   alphaCSR[ 193 ][ 209 ],
   alphaCSR[ 193 ][ 210 ],
   alphaCSR[ 193 ][ 211 ],
   alphaCSR[ 193 ][ 212 ],
   alphaCSR[ 193 ][ 213 ],
   alphaCSR[ 193 ][ 214 ],
   alphaCSR[ 193 ][ 215 ],
   alphaCSR[ 193 ][ 216 ],
   alphaCSR[ 193 ][ 217 ],
   alphaCSR[ 193 ][ 218 ],
   alphaCSR[ 193 ][ 219 ],
   alphaCSR[ 193 ][ 220 ],
   alphaCSR[ 193 ][ 221 ],
   alphaCSR[ 193 ][ 222 ],
   alphaCSR[ 193 ][ 223 ],
   alphaCSR[ 193 ][ 224 ],
   alphaCSR[ 193 ][ 225 ],
   alphaCSR[ 193 ][ 226 ],
   alphaCSR[ 193 ][ 227 ],
   alphaCSR[ 193 ][ 228 ],
   alphaCSR[ 193 ][ 229 ],
   alphaCSR[ 193 ][ 230 ],
   alphaCSR[ 193 ][ 231 ],
   alphaCSR[ 193 ][ 232 ],
   alphaCSR[ 193 ][ 233 ],
   alphaCSR[ 193 ][ 234 ],
   alphaCSR[ 193 ][ 235 ],
   alphaCSR[ 193 ][ 236 ],
   alphaCSR[ 193 ][ 237 ],
   alphaCSR[ 193 ][ 238 ],
   alphaCSR[ 193 ][ 239 ],
   alphaCSR[ 193 ][ 240 ],
   alphaCSR[ 193 ][ 241 ],
   alphaCSR[ 193 ][ 242 ],
   alphaCSR[ 193 ][ 243 ],
   alphaCSR[ 193 ][ 244 ],
   alphaCSR[ 193 ][ 245 ],
   alphaCSR[ 193 ][ 246 ],
   alphaCSR[ 193 ][ 247 ],
   alphaCSR[ 193 ][ 248 ],
   alphaCSR[ 193 ][ 249 ],
   alphaCSR[ 193 ][ 250 ],
   alphaCSR[ 193 ][ 251 ],
   alphaCSR[ 193 ][ 252 ],
   alphaCSR[ 193 ][ 253 ],
   alphaCSR[ 193 ][ 254 ],
   alphaCSR[ 193 ][ 255 ],
   alphaCSR[ 193 ][ 256 ],
   alphaCSR[ 193 ][ 257 ],
   alphaCSR[ 193 ][ 258 ],
   alphaCSR[ 193 ][ 259 ],
   alphaCSR[ 193 ][ 260 ],
   alphaCSR[ 193 ][ 261 ],
   alphaCSR[ 193 ][ 262 ],
   alphaCSR[ 193 ][ 263 ],
   alphaCSR[ 193 ][ 264 ],
   alphaCSR[ 193 ][ 265 ],
   alphaCSR[ 193 ][ 266 ],
   alphaCSR[ 193 ][ 267 ],
   alphaCSR[ 193 ][ 268 ],
   alphaCSR[ 193 ][ 269 ],
   alphaCSR[ 193 ][ 270 ],
   alphaCSR[ 193 ][ 271 ],
   alphaCSR[ 193 ][ 272 ],
   alphaCSR[ 193 ][ 273 ],
   alphaCSR[ 193 ][ 274 ],
   alphaCSR[ 193 ][ 275 ],
   alphaCSR[ 193 ][ 276 ],
   alphaCSR[ 193 ][ 277 ],
   alphaCSR[ 193 ][ 278 ],
   alphaCSR[ 193 ][ 279 ],
   alphaCSR[ 193 ][ 280 ],
   alphaCSR[ 193 ][ 281 ],
   alphaCSR[ 193 ][ 282 ],
   alphaCSR[ 193 ][ 283 ],
   alphaCSR[ 193 ][ 284 ],
   alphaCSR[ 193 ][ 285 ],
   alphaCSR[ 193 ][ 286 ],
   alphaCSR[ 193 ][ 287 ],
   alphaCSR[ 193 ][ 288 ],
   alphaCSR[ 193 ][ 289 ],
   alphaCSR[ 193 ][ 290 ],
   alphaCSR[ 193 ][ 291 ],
   alphaCSR[ 193 ][ 292 ],
   alphaCSR[ 193 ][ 293 ],
   alphaCSR[ 193 ][ 294 ],
   alphaCSR[ 193 ][ 295 ],
   alphaCSR[ 193 ][ 296 ],
   alphaCSR[ 193 ][ 297 ],
   alphaCSR[ 193 ][ 298 ],
   alphaCSR[ 193 ][ 299 ],
   alphaCSR[ 193 ][ 300 ],
   alphaCSR[ 193 ][ 301 ],
   alphaCSR[ 193 ][ 302 ],
   alphaCSR[ 193 ][ 303 ],
   alphaCSR[ 193 ][ 304 ],
   alphaCSR[ 193 ][ 305 ],
   alphaCSR[ 193 ][ 306 ],
   alphaCSR[ 193 ][ 307 ],
   alphaCSR[ 193 ][ 308 ],
   alphaCSR[ 193 ][ 309 ],
   alphaCSR[ 193 ][ 310 ],
   alphaCSR[ 193 ][ 311 ],
   alphaCSR[ 193 ][ 312 ],
   alphaCSR[ 193 ][ 313 ],
   alphaCSR[ 193 ][ 314 ],
   alphaCSR[ 193 ][ 315 ],
   alphaCSR[ 193 ][ 316 ],
   alphaCSR[ 193 ][ 317 ],
   alphaCSR[ 193 ][ 318 ],
   alphaCSR[ 193 ][ 319 ],
   alphaCSR[ 193 ][ 320 ],
   alphaCSR[ 193 ][ 321 ],
   alphaCSR[ 193 ][ 322 ],
   alphaCSR[ 193 ][ 323 ],
   alphaCSR[ 193 ][ 324 ],
   alphaCSR[ 193 ][ 325 ],
   alphaCSR[ 193 ][ 326 ],
   alphaCSR[ 193 ][ 327 ],
   alphaCSR[ 193 ][ 328 ],
   alphaCSR[ 193 ][ 329 ],
   alphaCSR[ 193 ][ 330 ],
   alphaCSR[ 193 ][ 331 ],
   alphaCSR[ 193 ][ 332 ],
   alphaCSR[ 193 ][ 333 ],
   alphaCSR[ 193 ][ 334 ],
   alphaCSR[ 193 ][ 335 ],
   alphaCSR[ 193 ][ 336 ],
   alphaCSR[ 193 ][ 337 ],
   alphaCSR[ 193 ][ 338 ],
   alphaCSR[ 193 ][ 339 ],
   alphaCSR[ 193 ][ 340 ],
   alphaCSR[ 193 ][ 341 ],
   alphaCSR[ 193 ][ 342 ],
   alphaCSR[ 193 ][ 343 ],
   alphaCSR[ 193 ][ 344 ],
   alphaCSR[ 193 ][ 345 ],
   alphaCSR[ 193 ][ 346 ],
   alphaCSR[ 193 ][ 347 ],
   alphaCSR[ 193 ][ 348 ],
   alphaCSR[ 193 ][ 349 ],
   alphaCSR[ 193 ][ 350 ],
   alphaCSR[ 193 ][ 351 ],
   alphaCSR[ 193 ][ 352 ],
   alphaCSR[ 193 ][ 353 ],
   alphaCSR[ 193 ][ 354 ],
   alphaCSR[ 193 ][ 355 ],
   alphaCSR[ 193 ][ 356 ],
   alphaCSR[ 193 ][ 357 ],
   alphaCSR[ 193 ][ 358 ],
   alphaCSR[ 193 ][ 359 ],
   alphaCSR[ 193 ][ 360 ],
   alphaCSR[ 193 ][ 361 ],
   alphaCSR[ 193 ][ 362 ],
   alphaCSR[ 193 ][ 363 ],
   alphaCSR[ 193 ][ 364 ],
   alphaCSR[ 193 ][ 365 ],
   alphaCSR[ 193 ][ 366 ],
   alphaCSR[ 193 ][ 367 ],
   alphaCSR[ 193 ][ 368 ],
   alphaCSR[ 193 ][ 369 ],
   alphaCSR[ 193 ][ 370 ],
   alphaCSR[ 193 ][ 371 ],
   alphaCSR[ 193 ][ 372 ],
   alphaCSR[ 193 ][ 373 ],
   alphaCSR[ 193 ][ 374 ],
   alphaCSR[ 193 ][ 375 ],
   alphaCSR[ 193 ][ 376 ],
   alphaCSR[ 193 ][ 377 ],
   alphaCSR[ 193 ][ 378 ],
   alphaCSR[ 193 ][ 379 ],
   alphaCSR[ 193 ][ 380 ],
   alphaCSR[ 193 ][ 381 ],
   alphaCSR[ 193 ][ 382 ],
   alphaCSR[ 193 ][ 383 ],
   alphaCSR[ 194 ][ 0 ],
   alphaCSR[ 194 ][ 1 ],
   alphaCSR[ 194 ][ 2 ],
   alphaCSR[ 194 ][ 3 ],
   alphaCSR[ 194 ][ 4 ],
   alphaCSR[ 194 ][ 5 ],
   alphaCSR[ 194 ][ 6 ],
   alphaCSR[ 194 ][ 7 ],
   alphaCSR[ 194 ][ 8 ],
   alphaCSR[ 194 ][ 9 ],
   alphaCSR[ 194 ][ 10 ],
   alphaCSR[ 194 ][ 11 ],
   alphaCSR[ 194 ][ 12 ],
   alphaCSR[ 194 ][ 13 ],
   alphaCSR[ 194 ][ 14 ],
   alphaCSR[ 194 ][ 15 ],
   alphaCSR[ 194 ][ 16 ],
   alphaCSR[ 194 ][ 17 ],
   alphaCSR[ 194 ][ 18 ],
   alphaCSR[ 194 ][ 19 ],
   alphaCSR[ 194 ][ 20 ],
   alphaCSR[ 194 ][ 21 ],
   alphaCSR[ 194 ][ 22 ],
   alphaCSR[ 194 ][ 23 ],
   alphaCSR[ 194 ][ 24 ],
   alphaCSR[ 194 ][ 25 ],
   alphaCSR[ 194 ][ 26 ],
   alphaCSR[ 194 ][ 27 ],
   alphaCSR[ 194 ][ 28 ],
   alphaCSR[ 194 ][ 29 ],
   alphaCSR[ 194 ][ 30 ],
   alphaCSR[ 194 ][ 31 ],
   alphaCSR[ 194 ][ 32 ],
   alphaCSR[ 194 ][ 33 ],
   alphaCSR[ 194 ][ 34 ],
   alphaCSR[ 194 ][ 35 ],
   alphaCSR[ 194 ][ 36 ],
   alphaCSR[ 194 ][ 37 ],
   alphaCSR[ 194 ][ 38 ],
   alphaCSR[ 194 ][ 39 ],
   alphaCSR[ 194 ][ 40 ],
   alphaCSR[ 194 ][ 41 ],
   alphaCSR[ 194 ][ 42 ],
   alphaCSR[ 194 ][ 43 ],
   alphaCSR[ 194 ][ 44 ],
   alphaCSR[ 194 ][ 45 ],
   alphaCSR[ 194 ][ 46 ],
   alphaCSR[ 194 ][ 47 ],
   alphaCSR[ 194 ][ 48 ],
   alphaCSR[ 194 ][ 49 ],
   alphaCSR[ 194 ][ 50 ],
   alphaCSR[ 194 ][ 51 ],
   alphaCSR[ 194 ][ 52 ],
   alphaCSR[ 194 ][ 53 ],
   alphaCSR[ 194 ][ 54 ],
   alphaCSR[ 194 ][ 55 ],
   alphaCSR[ 194 ][ 56 ],
   alphaCSR[ 194 ][ 57 ],
   alphaCSR[ 194 ][ 58 ],
   alphaCSR[ 194 ][ 59 ],
   alphaCSR[ 194 ][ 60 ],
   alphaCSR[ 194 ][ 61 ],
   alphaCSR[ 194 ][ 62 ],
   alphaCSR[ 194 ][ 63 ],
   alphaCSR[ 194 ][ 64 ],
   alphaCSR[ 194 ][ 65 ],
   alphaCSR[ 194 ][ 66 ],
   alphaCSR[ 194 ][ 67 ],
   alphaCSR[ 194 ][ 68 ],
   alphaCSR[ 194 ][ 69 ],
   alphaCSR[ 194 ][ 70 ],
   alphaCSR[ 194 ][ 71 ],
   alphaCSR[ 194 ][ 72 ],
   alphaCSR[ 194 ][ 73 ],
   alphaCSR[ 194 ][ 74 ],
   alphaCSR[ 194 ][ 75 ],
   alphaCSR[ 194 ][ 76 ],
   alphaCSR[ 194 ][ 77 ],
   alphaCSR[ 194 ][ 78 ],
   alphaCSR[ 194 ][ 79 ],
   alphaCSR[ 194 ][ 80 ],
   alphaCSR[ 194 ][ 81 ],
   alphaCSR[ 194 ][ 82 ],
   alphaCSR[ 194 ][ 83 ],
   alphaCSR[ 194 ][ 84 ],
   alphaCSR[ 194 ][ 85 ],
   alphaCSR[ 194 ][ 86 ],
   alphaCSR[ 194 ][ 87 ],
   alphaCSR[ 194 ][ 88 ],
   alphaCSR[ 194 ][ 89 ],
   alphaCSR[ 194 ][ 90 ],
   alphaCSR[ 194 ][ 91 ],
   alphaCSR[ 194 ][ 92 ],
   alphaCSR[ 194 ][ 93 ],
   alphaCSR[ 194 ][ 94 ],
   alphaCSR[ 194 ][ 95 ],
   alphaCSR[ 194 ][ 96 ],
   alphaCSR[ 194 ][ 97 ],
   alphaCSR[ 194 ][ 98 ],
   alphaCSR[ 194 ][ 99 ],
   alphaCSR[ 194 ][ 100 ],
   alphaCSR[ 194 ][ 101 ],
   alphaCSR[ 194 ][ 102 ],
   alphaCSR[ 194 ][ 103 ],
   alphaCSR[ 194 ][ 104 ],
   alphaCSR[ 194 ][ 105 ],
   alphaCSR[ 194 ][ 106 ],
   alphaCSR[ 194 ][ 107 ],
   alphaCSR[ 194 ][ 108 ],
   alphaCSR[ 194 ][ 109 ],
   alphaCSR[ 194 ][ 110 ],
   alphaCSR[ 194 ][ 111 ],
   alphaCSR[ 194 ][ 112 ],
   alphaCSR[ 194 ][ 113 ],
   alphaCSR[ 194 ][ 114 ],
   alphaCSR[ 194 ][ 115 ],
   alphaCSR[ 194 ][ 116 ],
   alphaCSR[ 194 ][ 117 ],
   alphaCSR[ 194 ][ 118 ],
   alphaCSR[ 194 ][ 119 ],
   alphaCSR[ 194 ][ 120 ],
   alphaCSR[ 194 ][ 121 ],
   alphaCSR[ 194 ][ 122 ],
   alphaCSR[ 194 ][ 123 ],
   alphaCSR[ 194 ][ 124 ],
   alphaCSR[ 194 ][ 125 ],
   alphaCSR[ 194 ][ 126 ],
   alphaCSR[ 194 ][ 127 ],
   alphaCSR[ 194 ][ 128 ],
   alphaCSR[ 194 ][ 129 ],
   alphaCSR[ 194 ][ 130 ],
   alphaCSR[ 194 ][ 131 ],
   alphaCSR[ 194 ][ 132 ],
   alphaCSR[ 194 ][ 133 ],
   alphaCSR[ 194 ][ 134 ],
   alphaCSR[ 194 ][ 135 ],
   alphaCSR[ 194 ][ 136 ],
   alphaCSR[ 194 ][ 137 ],
   alphaCSR[ 194 ][ 138 ],
   alphaCSR[ 194 ][ 139 ],
   alphaCSR[ 194 ][ 140 ],
   alphaCSR[ 194 ][ 141 ],
   alphaCSR[ 194 ][ 142 ],
   alphaCSR[ 194 ][ 143 ],
   alphaCSR[ 194 ][ 144 ],
   alphaCSR[ 194 ][ 145 ],
   alphaCSR[ 194 ][ 146 ],
   alphaCSR[ 194 ][ 147 ],
   alphaCSR[ 194 ][ 148 ],
   alphaCSR[ 194 ][ 149 ],
   alphaCSR[ 194 ][ 150 ],
   alphaCSR[ 194 ][ 151 ],
   alphaCSR[ 194 ][ 152 ],
   alphaCSR[ 194 ][ 153 ],
   alphaCSR[ 194 ][ 154 ],
   alphaCSR[ 194 ][ 155 ],
   alphaCSR[ 194 ][ 156 ],
   alphaCSR[ 194 ][ 157 ],
   alphaCSR[ 194 ][ 158 ],
   alphaCSR[ 194 ][ 159 ],
   alphaCSR[ 194 ][ 160 ],
   alphaCSR[ 194 ][ 161 ],
   alphaCSR[ 194 ][ 162 ],
   alphaCSR[ 194 ][ 163 ],
   alphaCSR[ 194 ][ 164 ],
   alphaCSR[ 194 ][ 165 ],
   alphaCSR[ 194 ][ 166 ],
   alphaCSR[ 194 ][ 167 ],
   alphaCSR[ 194 ][ 168 ],
   alphaCSR[ 194 ][ 169 ],
   alphaCSR[ 194 ][ 170 ],
   alphaCSR[ 194 ][ 171 ],
   alphaCSR[ 194 ][ 172 ],
   alphaCSR[ 194 ][ 173 ],
   alphaCSR[ 194 ][ 174 ],
   alphaCSR[ 194 ][ 175 ],
   alphaCSR[ 194 ][ 176 ],
   alphaCSR[ 194 ][ 177 ],
   alphaCSR[ 194 ][ 178 ],
   alphaCSR[ 194 ][ 179 ],
   alphaCSR[ 194 ][ 180 ],
   alphaCSR[ 194 ][ 181 ],
   alphaCSR[ 194 ][ 182 ],
   alphaCSR[ 194 ][ 183 ],
   alphaCSR[ 194 ][ 184 ],
   alphaCSR[ 194 ][ 185 ],
   alphaCSR[ 194 ][ 186 ],
   alphaCSR[ 194 ][ 187 ],
   alphaCSR[ 194 ][ 188 ],
   alphaCSR[ 194 ][ 189 ],
   alphaCSR[ 194 ][ 190 ],
   alphaCSR[ 194 ][ 191 ],
   alphaCSR[ 194 ][ 192 ],
   alphaCSR[ 194 ][ 193 ],
   alphaCSR[ 194 ][ 194 ],
   alphaCSR[ 194 ][ 195 ],
   alphaCSR[ 194 ][ 196 ],
   alphaCSR[ 194 ][ 197 ],
   alphaCSR[ 194 ][ 198 ],
   alphaCSR[ 194 ][ 199 ],
   alphaCSR[ 194 ][ 200 ],
   alphaCSR[ 194 ][ 201 ],
   alphaCSR[ 194 ][ 202 ],
   alphaCSR[ 194 ][ 203 ],
   alphaCSR[ 194 ][ 204 ],
   alphaCSR[ 194 ][ 205 ],
   alphaCSR[ 194 ][ 206 ],
   alphaCSR[ 194 ][ 207 ],
   alphaCSR[ 194 ][ 208 ],
   alphaCSR[ 194 ][ 209 ],
   alphaCSR[ 194 ][ 210 ],
   alphaCSR[ 194 ][ 211 ],
   alphaCSR[ 194 ][ 212 ],
   alphaCSR[ 194 ][ 213 ],
   alphaCSR[ 194 ][ 214 ],
   alphaCSR[ 194 ][ 215 ],
   alphaCSR[ 194 ][ 216 ],
   alphaCSR[ 194 ][ 217 ],
   alphaCSR[ 194 ][ 218 ],
   alphaCSR[ 194 ][ 219 ],
   alphaCSR[ 194 ][ 220 ],
   alphaCSR[ 194 ][ 221 ],
   alphaCSR[ 194 ][ 222 ],
   alphaCSR[ 194 ][ 223 ],
   alphaCSR[ 194 ][ 224 ],
   alphaCSR[ 194 ][ 225 ],
   alphaCSR[ 194 ][ 226 ],
   alphaCSR[ 194 ][ 227 ],
   alphaCSR[ 194 ][ 228 ],
   alphaCSR[ 194 ][ 229 ],
   alphaCSR[ 194 ][ 230 ],
   alphaCSR[ 194 ][ 231 ],
   alphaCSR[ 194 ][ 232 ],
   alphaCSR[ 194 ][ 233 ],
   alphaCSR[ 194 ][ 234 ],
   alphaCSR[ 194 ][ 235 ],
   alphaCSR[ 194 ][ 236 ],
   alphaCSR[ 194 ][ 237 ],
   alphaCSR[ 194 ][ 238 ],
   alphaCSR[ 194 ][ 239 ],
   alphaCSR[ 194 ][ 240 ],
   alphaCSR[ 194 ][ 241 ],
   alphaCSR[ 194 ][ 242 ],
   alphaCSR[ 194 ][ 243 ],
   alphaCSR[ 194 ][ 244 ],
   alphaCSR[ 194 ][ 245 ],
   alphaCSR[ 194 ][ 246 ],
   alphaCSR[ 194 ][ 247 ],
   alphaCSR[ 194 ][ 248 ],
   alphaCSR[ 194 ][ 249 ],
   alphaCSR[ 194 ][ 250 ],
   alphaCSR[ 194 ][ 251 ],
   alphaCSR[ 194 ][ 252 ],
   alphaCSR[ 194 ][ 253 ],
   alphaCSR[ 194 ][ 254 ],
   alphaCSR[ 194 ][ 255 ],
   alphaCSR[ 194 ][ 256 ],
   alphaCSR[ 194 ][ 257 ],
   alphaCSR[ 194 ][ 258 ],
   alphaCSR[ 194 ][ 259 ],
   alphaCSR[ 194 ][ 260 ],
   alphaCSR[ 194 ][ 261 ],
   alphaCSR[ 194 ][ 262 ],
   alphaCSR[ 194 ][ 263 ],
   alphaCSR[ 194 ][ 264 ],
   alphaCSR[ 194 ][ 265 ],
   alphaCSR[ 194 ][ 266 ],
   alphaCSR[ 194 ][ 267 ],
   alphaCSR[ 194 ][ 268 ],
   alphaCSR[ 194 ][ 269 ],
   alphaCSR[ 194 ][ 270 ],
   alphaCSR[ 194 ][ 271 ],
   alphaCSR[ 194 ][ 272 ],
   alphaCSR[ 194 ][ 273 ],
   alphaCSR[ 194 ][ 274 ],
   alphaCSR[ 194 ][ 275 ],
   alphaCSR[ 194 ][ 276 ],
   alphaCSR[ 194 ][ 277 ],
   alphaCSR[ 194 ][ 278 ],
   alphaCSR[ 194 ][ 279 ],
   alphaCSR[ 194 ][ 280 ],
   alphaCSR[ 194 ][ 281 ],
   alphaCSR[ 194 ][ 282 ],
   alphaCSR[ 194 ][ 283 ],
   alphaCSR[ 194 ][ 284 ],
   alphaCSR[ 194 ][ 285 ],
   alphaCSR[ 194 ][ 286 ],
   alphaCSR[ 194 ][ 287 ],
   alphaCSR[ 194 ][ 288 ],
   alphaCSR[ 194 ][ 289 ],
   alphaCSR[ 194 ][ 290 ],
   alphaCSR[ 194 ][ 291 ],
   alphaCSR[ 194 ][ 292 ],
   alphaCSR[ 194 ][ 293 ],
   alphaCSR[ 194 ][ 294 ],
   alphaCSR[ 194 ][ 295 ],
   alphaCSR[ 194 ][ 296 ],
   alphaCSR[ 194 ][ 297 ],
   alphaCSR[ 194 ][ 298 ],
   alphaCSR[ 194 ][ 299 ],
   alphaCSR[ 194 ][ 300 ],
   alphaCSR[ 194 ][ 301 ],
   alphaCSR[ 194 ][ 302 ],
   alphaCSR[ 194 ][ 303 ],
   alphaCSR[ 194 ][ 304 ],
   alphaCSR[ 194 ][ 305 ],
   alphaCSR[ 194 ][ 306 ],
   alphaCSR[ 194 ][ 307 ],
   alphaCSR[ 194 ][ 308 ],
   alphaCSR[ 194 ][ 309 ],
   alphaCSR[ 194 ][ 310 ],
   alphaCSR[ 194 ][ 311 ],
   alphaCSR[ 194 ][ 312 ],
   alphaCSR[ 194 ][ 313 ],
   alphaCSR[ 194 ][ 314 ],
   alphaCSR[ 194 ][ 315 ],
   alphaCSR[ 194 ][ 316 ],
   alphaCSR[ 194 ][ 317 ],
   alphaCSR[ 194 ][ 318 ],
   alphaCSR[ 194 ][ 319 ],
   alphaCSR[ 194 ][ 320 ],
   alphaCSR[ 194 ][ 321 ],
   alphaCSR[ 194 ][ 322 ],
   alphaCSR[ 194 ][ 323 ],
   alphaCSR[ 194 ][ 324 ],
   alphaCSR[ 194 ][ 325 ],
   alphaCSR[ 194 ][ 326 ],
   alphaCSR[ 194 ][ 327 ],
   alphaCSR[ 194 ][ 328 ],
   alphaCSR[ 194 ][ 329 ],
   alphaCSR[ 194 ][ 330 ],
   alphaCSR[ 194 ][ 331 ],
   alphaCSR[ 194 ][ 332 ],
   alphaCSR[ 194 ][ 333 ],
   alphaCSR[ 194 ][ 334 ],
   alphaCSR[ 194 ][ 335 ],
   alphaCSR[ 194 ][ 336 ],
   alphaCSR[ 194 ][ 337 ],
   alphaCSR[ 194 ][ 338 ],
   alphaCSR[ 194 ][ 339 ],
   alphaCSR[ 194 ][ 340 ],
   alphaCSR[ 194 ][ 341 ],
   alphaCSR[ 194 ][ 342 ],
   alphaCSR[ 194 ][ 343 ],
   alphaCSR[ 194 ][ 344 ],
   alphaCSR[ 194 ][ 345 ],
   alphaCSR[ 194 ][ 346 ],
   alphaCSR[ 194 ][ 347 ],
   alphaCSR[ 194 ][ 348 ],
   alphaCSR[ 194 ][ 349 ],
   alphaCSR[ 194 ][ 350 ],
   alphaCSR[ 194 ][ 351 ],
   alphaCSR[ 194 ][ 352 ],
   alphaCSR[ 194 ][ 353 ],
   alphaCSR[ 194 ][ 354 ],
   alphaCSR[ 194 ][ 355 ],
   alphaCSR[ 194 ][ 356 ],
   alphaCSR[ 194 ][ 357 ],
   alphaCSR[ 194 ][ 358 ],
   alphaCSR[ 194 ][ 359 ],
   alphaCSR[ 194 ][ 360 ],
   alphaCSR[ 194 ][ 361 ],
   alphaCSR[ 194 ][ 362 ],
   alphaCSR[ 194 ][ 363 ],
   alphaCSR[ 194 ][ 364 ],
   alphaCSR[ 194 ][ 365 ],
   alphaCSR[ 194 ][ 366 ],
   alphaCSR[ 194 ][ 367 ],
   alphaCSR[ 194 ][ 368 ],
   alphaCSR[ 194 ][ 369 ],
   alphaCSR[ 194 ][ 370 ],
   alphaCSR[ 194 ][ 371 ],
   alphaCSR[ 194 ][ 372 ],
   alphaCSR[ 194 ][ 373 ],
   alphaCSR[ 194 ][ 374 ],
   alphaCSR[ 194 ][ 375 ],
   alphaCSR[ 194 ][ 376 ],
   alphaCSR[ 194 ][ 377 ],
   alphaCSR[ 194 ][ 378 ],
   alphaCSR[ 194 ][ 379 ],
   alphaCSR[ 194 ][ 380 ],
   alphaCSR[ 194 ][ 381 ],
   alphaCSR[ 194 ][ 382 ],
   alphaCSR[ 194 ][ 383 ],
   alphaCSR[ 195 ][ 0 ],
   alphaCSR[ 195 ][ 1 ],
   alphaCSR[ 195 ][ 2 ],
   alphaCSR[ 195 ][ 3 ],
   alphaCSR[ 195 ][ 4 ],
   alphaCSR[ 195 ][ 5 ],
   alphaCSR[ 195 ][ 6 ],
   alphaCSR[ 195 ][ 7 ],
   alphaCSR[ 195 ][ 8 ],
   alphaCSR[ 195 ][ 9 ],
   alphaCSR[ 195 ][ 10 ],
   alphaCSR[ 195 ][ 11 ],
   alphaCSR[ 195 ][ 12 ],
   alphaCSR[ 195 ][ 13 ],
   alphaCSR[ 195 ][ 14 ],
   alphaCSR[ 195 ][ 15 ],
   alphaCSR[ 195 ][ 16 ],
   alphaCSR[ 195 ][ 17 ],
   alphaCSR[ 195 ][ 18 ],
   alphaCSR[ 195 ][ 19 ],
   alphaCSR[ 195 ][ 20 ],
   alphaCSR[ 195 ][ 21 ],
   alphaCSR[ 195 ][ 22 ],
   alphaCSR[ 195 ][ 23 ],
   alphaCSR[ 195 ][ 24 ],
   alphaCSR[ 195 ][ 25 ],
   alphaCSR[ 195 ][ 26 ],
   alphaCSR[ 195 ][ 27 ],
   alphaCSR[ 195 ][ 28 ],
   alphaCSR[ 195 ][ 29 ],
   alphaCSR[ 195 ][ 30 ],
   alphaCSR[ 195 ][ 31 ],
   alphaCSR[ 195 ][ 32 ],
   alphaCSR[ 195 ][ 33 ],
   alphaCSR[ 195 ][ 34 ],
   alphaCSR[ 195 ][ 35 ],
   alphaCSR[ 195 ][ 36 ],
   alphaCSR[ 195 ][ 37 ],
   alphaCSR[ 195 ][ 38 ],
   alphaCSR[ 195 ][ 39 ],
   alphaCSR[ 195 ][ 40 ],
   alphaCSR[ 195 ][ 41 ],
   alphaCSR[ 195 ][ 42 ],
   alphaCSR[ 195 ][ 43 ],
   alphaCSR[ 195 ][ 44 ],
   alphaCSR[ 195 ][ 45 ],
   alphaCSR[ 195 ][ 46 ],
   alphaCSR[ 195 ][ 47 ],
   alphaCSR[ 195 ][ 48 ],
   alphaCSR[ 195 ][ 49 ],
   alphaCSR[ 195 ][ 50 ],
   alphaCSR[ 195 ][ 51 ],
   alphaCSR[ 195 ][ 52 ],
   alphaCSR[ 195 ][ 53 ],
   alphaCSR[ 195 ][ 54 ],
   alphaCSR[ 195 ][ 55 ],
   alphaCSR[ 195 ][ 56 ],
   alphaCSR[ 195 ][ 57 ],
   alphaCSR[ 195 ][ 58 ],
   alphaCSR[ 195 ][ 59 ],
   alphaCSR[ 195 ][ 60 ],
   alphaCSR[ 195 ][ 61 ],
   alphaCSR[ 195 ][ 62 ],
   alphaCSR[ 195 ][ 63 ],
   alphaCSR[ 195 ][ 64 ],
   alphaCSR[ 195 ][ 65 ],
   alphaCSR[ 195 ][ 66 ],
   alphaCSR[ 195 ][ 67 ],
   alphaCSR[ 195 ][ 68 ],
   alphaCSR[ 195 ][ 69 ],
   alphaCSR[ 195 ][ 70 ],
   alphaCSR[ 195 ][ 71 ],
   alphaCSR[ 195 ][ 72 ],
   alphaCSR[ 195 ][ 73 ],
   alphaCSR[ 195 ][ 74 ],
   alphaCSR[ 195 ][ 75 ],
   alphaCSR[ 195 ][ 76 ],
   alphaCSR[ 195 ][ 77 ],
   alphaCSR[ 195 ][ 78 ],
   alphaCSR[ 195 ][ 79 ],
   alphaCSR[ 195 ][ 80 ],
   alphaCSR[ 195 ][ 81 ],
   alphaCSR[ 195 ][ 82 ],
   alphaCSR[ 195 ][ 83 ],
   alphaCSR[ 195 ][ 84 ],
   alphaCSR[ 195 ][ 85 ],
   alphaCSR[ 195 ][ 86 ],
   alphaCSR[ 195 ][ 87 ],
   alphaCSR[ 195 ][ 88 ],
   alphaCSR[ 195 ][ 89 ],
   alphaCSR[ 195 ][ 90 ],
   alphaCSR[ 195 ][ 91 ],
   alphaCSR[ 195 ][ 92 ],
   alphaCSR[ 195 ][ 93 ],
   alphaCSR[ 195 ][ 94 ],
   alphaCSR[ 195 ][ 95 ],
   alphaCSR[ 195 ][ 96 ],
   alphaCSR[ 195 ][ 97 ],
   alphaCSR[ 195 ][ 98 ],
   alphaCSR[ 195 ][ 99 ],
   alphaCSR[ 195 ][ 100 ],
   alphaCSR[ 195 ][ 101 ],
   alphaCSR[ 195 ][ 102 ],
   alphaCSR[ 195 ][ 103 ],
   alphaCSR[ 195 ][ 104 ],
   alphaCSR[ 195 ][ 105 ],
   alphaCSR[ 195 ][ 106 ],
   alphaCSR[ 195 ][ 107 ],
   alphaCSR[ 195 ][ 108 ],
   alphaCSR[ 195 ][ 109 ],
   alphaCSR[ 195 ][ 110 ],
   alphaCSR[ 195 ][ 111 ],
   alphaCSR[ 195 ][ 112 ],
   alphaCSR[ 195 ][ 113 ],
   alphaCSR[ 195 ][ 114 ],
   alphaCSR[ 195 ][ 115 ],
   alphaCSR[ 195 ][ 116 ],
   alphaCSR[ 195 ][ 117 ],
   alphaCSR[ 195 ][ 118 ],
   alphaCSR[ 195 ][ 119 ],
   alphaCSR[ 195 ][ 120 ],
   alphaCSR[ 195 ][ 121 ],
   alphaCSR[ 195 ][ 122 ],
   alphaCSR[ 195 ][ 123 ],
   alphaCSR[ 195 ][ 124 ],
   alphaCSR[ 195 ][ 125 ],
   alphaCSR[ 195 ][ 126 ],
   alphaCSR[ 195 ][ 127 ],
   alphaCSR[ 195 ][ 128 ],
   alphaCSR[ 195 ][ 129 ],
   alphaCSR[ 195 ][ 130 ],
   alphaCSR[ 195 ][ 131 ],
   alphaCSR[ 195 ][ 132 ],
   alphaCSR[ 195 ][ 133 ],
   alphaCSR[ 195 ][ 134 ],
   alphaCSR[ 195 ][ 135 ],
   alphaCSR[ 195 ][ 136 ],
   alphaCSR[ 195 ][ 137 ],
   alphaCSR[ 195 ][ 138 ],
   alphaCSR[ 195 ][ 139 ],
   alphaCSR[ 195 ][ 140 ],
   alphaCSR[ 195 ][ 141 ],
   alphaCSR[ 195 ][ 142 ],
   alphaCSR[ 195 ][ 143 ],
   alphaCSR[ 195 ][ 144 ],
   alphaCSR[ 195 ][ 145 ],
   alphaCSR[ 195 ][ 146 ],
   alphaCSR[ 195 ][ 147 ],
   alphaCSR[ 195 ][ 148 ],
   alphaCSR[ 195 ][ 149 ],
   alphaCSR[ 195 ][ 150 ],
   alphaCSR[ 195 ][ 151 ],
   alphaCSR[ 195 ][ 152 ],
   alphaCSR[ 195 ][ 153 ],
   alphaCSR[ 195 ][ 154 ],
   alphaCSR[ 195 ][ 155 ],
   alphaCSR[ 195 ][ 156 ],
   alphaCSR[ 195 ][ 157 ],
   alphaCSR[ 195 ][ 158 ],
   alphaCSR[ 195 ][ 159 ],
   alphaCSR[ 195 ][ 160 ],
   alphaCSR[ 195 ][ 161 ],
   alphaCSR[ 195 ][ 162 ],
   alphaCSR[ 195 ][ 163 ],
   alphaCSR[ 195 ][ 164 ],
   alphaCSR[ 195 ][ 165 ],
   alphaCSR[ 195 ][ 166 ],
   alphaCSR[ 195 ][ 167 ],
   alphaCSR[ 195 ][ 168 ],
   alphaCSR[ 195 ][ 169 ],
   alphaCSR[ 195 ][ 170 ],
   alphaCSR[ 195 ][ 171 ],
   alphaCSR[ 195 ][ 172 ],
   alphaCSR[ 195 ][ 173 ],
   alphaCSR[ 195 ][ 174 ],
   alphaCSR[ 195 ][ 175 ],
   alphaCSR[ 195 ][ 176 ],
   alphaCSR[ 195 ][ 177 ],
   alphaCSR[ 195 ][ 178 ],
   alphaCSR[ 195 ][ 179 ],
   alphaCSR[ 195 ][ 180 ],
   alphaCSR[ 195 ][ 181 ],
   alphaCSR[ 195 ][ 182 ],
   alphaCSR[ 195 ][ 183 ],
   alphaCSR[ 195 ][ 184 ],
   alphaCSR[ 195 ][ 185 ],
   alphaCSR[ 195 ][ 186 ],
   alphaCSR[ 195 ][ 187 ],
   alphaCSR[ 195 ][ 188 ],
   alphaCSR[ 195 ][ 189 ],
   alphaCSR[ 195 ][ 190 ],
   alphaCSR[ 195 ][ 191 ],
   alphaCSR[ 195 ][ 192 ],
   alphaCSR[ 195 ][ 193 ],
   alphaCSR[ 195 ][ 194 ],
   alphaCSR[ 195 ][ 195 ],
   alphaCSR[ 195 ][ 196 ],
   alphaCSR[ 195 ][ 197 ],
   alphaCSR[ 195 ][ 198 ],
   alphaCSR[ 195 ][ 199 ],
   alphaCSR[ 195 ][ 200 ],
   alphaCSR[ 195 ][ 201 ],
   alphaCSR[ 195 ][ 202 ],
   alphaCSR[ 195 ][ 203 ],
   alphaCSR[ 195 ][ 204 ],
   alphaCSR[ 195 ][ 205 ],
   alphaCSR[ 195 ][ 206 ],
   alphaCSR[ 195 ][ 207 ],
   alphaCSR[ 195 ][ 208 ],
   alphaCSR[ 195 ][ 209 ],
   alphaCSR[ 195 ][ 210 ],
   alphaCSR[ 195 ][ 211 ],
   alphaCSR[ 195 ][ 212 ],
   alphaCSR[ 195 ][ 213 ],
   alphaCSR[ 195 ][ 214 ],
   alphaCSR[ 195 ][ 215 ],
   alphaCSR[ 195 ][ 216 ],
   alphaCSR[ 195 ][ 217 ],
   alphaCSR[ 195 ][ 218 ],
   alphaCSR[ 195 ][ 219 ],
   alphaCSR[ 195 ][ 220 ],
   alphaCSR[ 195 ][ 221 ],
   alphaCSR[ 195 ][ 222 ],
   alphaCSR[ 195 ][ 223 ],
   alphaCSR[ 195 ][ 224 ],
   alphaCSR[ 195 ][ 225 ],
   alphaCSR[ 195 ][ 226 ],
   alphaCSR[ 195 ][ 227 ],
   alphaCSR[ 195 ][ 228 ],
   alphaCSR[ 195 ][ 229 ],
   alphaCSR[ 195 ][ 230 ],
   alphaCSR[ 195 ][ 231 ],
   alphaCSR[ 195 ][ 232 ],
   alphaCSR[ 195 ][ 233 ],
   alphaCSR[ 195 ][ 234 ],
   alphaCSR[ 195 ][ 235 ],
   alphaCSR[ 195 ][ 236 ],
   alphaCSR[ 195 ][ 237 ],
   alphaCSR[ 195 ][ 238 ],
   alphaCSR[ 195 ][ 239 ],
   alphaCSR[ 195 ][ 240 ],
   alphaCSR[ 195 ][ 241 ],
   alphaCSR[ 195 ][ 242 ],
   alphaCSR[ 195 ][ 243 ],
   alphaCSR[ 195 ][ 244 ],
   alphaCSR[ 195 ][ 245 ],
   alphaCSR[ 195 ][ 246 ],
   alphaCSR[ 195 ][ 247 ],
   alphaCSR[ 195 ][ 248 ],
   alphaCSR[ 195 ][ 249 ],
   alphaCSR[ 195 ][ 250 ],
   alphaCSR[ 195 ][ 251 ],
   alphaCSR[ 195 ][ 252 ],
   alphaCSR[ 195 ][ 253 ],
   alphaCSR[ 195 ][ 254 ],
   alphaCSR[ 195 ][ 255 ],
   alphaCSR[ 195 ][ 256 ],
   alphaCSR[ 195 ][ 257 ],
   alphaCSR[ 195 ][ 258 ],
   alphaCSR[ 195 ][ 259 ],
   alphaCSR[ 195 ][ 260 ],
   alphaCSR[ 195 ][ 261 ],
   alphaCSR[ 195 ][ 262 ],
   alphaCSR[ 195 ][ 263 ],
   alphaCSR[ 195 ][ 264 ],
   alphaCSR[ 195 ][ 265 ],
   alphaCSR[ 195 ][ 266 ],
   alphaCSR[ 195 ][ 267 ],
   alphaCSR[ 195 ][ 268 ],
   alphaCSR[ 195 ][ 269 ],
   alphaCSR[ 195 ][ 270 ],
   alphaCSR[ 195 ][ 271 ],
   alphaCSR[ 195 ][ 272 ],
   alphaCSR[ 195 ][ 273 ],
   alphaCSR[ 195 ][ 274 ],
   alphaCSR[ 195 ][ 275 ],
   alphaCSR[ 195 ][ 276 ],
   alphaCSR[ 195 ][ 277 ],
   alphaCSR[ 195 ][ 278 ],
   alphaCSR[ 195 ][ 279 ],
   alphaCSR[ 195 ][ 280 ],
   alphaCSR[ 195 ][ 281 ],
   alphaCSR[ 195 ][ 282 ],
   alphaCSR[ 195 ][ 283 ],
   alphaCSR[ 195 ][ 284 ],
   alphaCSR[ 195 ][ 285 ],
   alphaCSR[ 195 ][ 286 ],
   alphaCSR[ 195 ][ 287 ],
   alphaCSR[ 195 ][ 288 ],
   alphaCSR[ 195 ][ 289 ],
   alphaCSR[ 195 ][ 290 ],
   alphaCSR[ 195 ][ 291 ],
   alphaCSR[ 195 ][ 292 ],
   alphaCSR[ 195 ][ 293 ],
   alphaCSR[ 195 ][ 294 ],
   alphaCSR[ 195 ][ 295 ],
   alphaCSR[ 195 ][ 296 ],
   alphaCSR[ 195 ][ 297 ],
   alphaCSR[ 195 ][ 298 ],
   alphaCSR[ 195 ][ 299 ],
   alphaCSR[ 195 ][ 300 ],
   alphaCSR[ 195 ][ 301 ],
   alphaCSR[ 195 ][ 302 ],
   alphaCSR[ 195 ][ 303 ],
   alphaCSR[ 195 ][ 304 ],
   alphaCSR[ 195 ][ 305 ],
   alphaCSR[ 195 ][ 306 ],
   alphaCSR[ 195 ][ 307 ],
   alphaCSR[ 195 ][ 308 ],
   alphaCSR[ 195 ][ 309 ],
   alphaCSR[ 195 ][ 310 ],
   alphaCSR[ 195 ][ 311 ],
   alphaCSR[ 195 ][ 312 ],
   alphaCSR[ 195 ][ 313 ],
   alphaCSR[ 195 ][ 314 ],
   alphaCSR[ 195 ][ 315 ],
   alphaCSR[ 195 ][ 316 ],
   alphaCSR[ 195 ][ 317 ],
   alphaCSR[ 195 ][ 318 ],
   alphaCSR[ 195 ][ 319 ],
   alphaCSR[ 195 ][ 320 ],
   alphaCSR[ 195 ][ 321 ],
   alphaCSR[ 195 ][ 322 ],
   alphaCSR[ 195 ][ 323 ],
   alphaCSR[ 195 ][ 324 ],
   alphaCSR[ 195 ][ 325 ],
   alphaCSR[ 195 ][ 326 ],
   alphaCSR[ 195 ][ 327 ],
   alphaCSR[ 195 ][ 328 ],
   alphaCSR[ 195 ][ 329 ],
   alphaCSR[ 195 ][ 330 ],
   alphaCSR[ 195 ][ 331 ],
   alphaCSR[ 195 ][ 332 ],
   alphaCSR[ 195 ][ 333 ],
   alphaCSR[ 195 ][ 334 ],
   alphaCSR[ 195 ][ 335 ],
   alphaCSR[ 195 ][ 336 ],
   alphaCSR[ 195 ][ 337 ],
   alphaCSR[ 195 ][ 338 ],
   alphaCSR[ 195 ][ 339 ],
   alphaCSR[ 195 ][ 340 ],
   alphaCSR[ 195 ][ 341 ],
   alphaCSR[ 195 ][ 342 ],
   alphaCSR[ 195 ][ 343 ],
   alphaCSR[ 195 ][ 344 ],
   alphaCSR[ 195 ][ 345 ],
   alphaCSR[ 195 ][ 346 ],
   alphaCSR[ 195 ][ 347 ],
   alphaCSR[ 195 ][ 348 ],
   alphaCSR[ 195 ][ 349 ],
   alphaCSR[ 195 ][ 350 ],
   alphaCSR[ 195 ][ 351 ],
   alphaCSR[ 195 ][ 352 ],
   alphaCSR[ 195 ][ 353 ],
   alphaCSR[ 195 ][ 354 ],
   alphaCSR[ 195 ][ 355 ],
   alphaCSR[ 195 ][ 356 ],
   alphaCSR[ 195 ][ 357 ],
   alphaCSR[ 195 ][ 358 ],
   alphaCSR[ 195 ][ 359 ],
   alphaCSR[ 195 ][ 360 ],
   alphaCSR[ 195 ][ 361 ],
   alphaCSR[ 195 ][ 362 ],
   alphaCSR[ 195 ][ 363 ],
   alphaCSR[ 195 ][ 364 ],
   alphaCSR[ 195 ][ 365 ],
   alphaCSR[ 195 ][ 366 ],
   alphaCSR[ 195 ][ 367 ],
   alphaCSR[ 195 ][ 368 ],
   alphaCSR[ 195 ][ 369 ],
   alphaCSR[ 195 ][ 370 ],
   alphaCSR[ 195 ][ 371 ],
   alphaCSR[ 195 ][ 372 ],
   alphaCSR[ 195 ][ 373 ],
   alphaCSR[ 195 ][ 374 ],
   alphaCSR[ 195 ][ 375 ],
   alphaCSR[ 195 ][ 376 ],
   alphaCSR[ 195 ][ 377 ],
   alphaCSR[ 195 ][ 378 ],
   alphaCSR[ 195 ][ 379 ],
   alphaCSR[ 195 ][ 380 ],
   alphaCSR[ 195 ][ 381 ],
   alphaCSR[ 195 ][ 382 ],
   alphaCSR[ 195 ][ 383 ],
   alphaCSR[ 196 ][ 0 ],
   alphaCSR[ 196 ][ 1 ],
   alphaCSR[ 196 ][ 2 ],
   alphaCSR[ 196 ][ 3 ],
   alphaCSR[ 196 ][ 4 ],
   alphaCSR[ 196 ][ 5 ],
   alphaCSR[ 196 ][ 6 ],
   alphaCSR[ 196 ][ 7 ],
   alphaCSR[ 196 ][ 8 ],
   alphaCSR[ 196 ][ 9 ],
   alphaCSR[ 196 ][ 10 ],
   alphaCSR[ 196 ][ 11 ],
   alphaCSR[ 196 ][ 12 ],
   alphaCSR[ 196 ][ 13 ],
   alphaCSR[ 196 ][ 14 ],
   alphaCSR[ 196 ][ 15 ],
   alphaCSR[ 196 ][ 16 ],
   alphaCSR[ 196 ][ 17 ],
   alphaCSR[ 196 ][ 18 ],
   alphaCSR[ 196 ][ 19 ],
   alphaCSR[ 196 ][ 20 ],
   alphaCSR[ 196 ][ 21 ],
   alphaCSR[ 196 ][ 22 ],
   alphaCSR[ 196 ][ 23 ],
   alphaCSR[ 196 ][ 24 ],
   alphaCSR[ 196 ][ 25 ],
   alphaCSR[ 196 ][ 26 ],
   alphaCSR[ 196 ][ 27 ],
   alphaCSR[ 196 ][ 28 ],
   alphaCSR[ 196 ][ 29 ],
   alphaCSR[ 196 ][ 30 ],
   alphaCSR[ 196 ][ 31 ],
   alphaCSR[ 196 ][ 32 ],
   alphaCSR[ 196 ][ 33 ],
   alphaCSR[ 196 ][ 34 ],
   alphaCSR[ 196 ][ 35 ],
   alphaCSR[ 196 ][ 36 ],
   alphaCSR[ 196 ][ 37 ],
   alphaCSR[ 196 ][ 38 ],
   alphaCSR[ 196 ][ 39 ],
   alphaCSR[ 196 ][ 40 ],
   alphaCSR[ 196 ][ 41 ],
   alphaCSR[ 196 ][ 42 ],
   alphaCSR[ 196 ][ 43 ],
   alphaCSR[ 196 ][ 44 ],
   alphaCSR[ 196 ][ 45 ],
   alphaCSR[ 196 ][ 46 ],
   alphaCSR[ 196 ][ 47 ],
   alphaCSR[ 196 ][ 48 ],
   alphaCSR[ 196 ][ 49 ],
   alphaCSR[ 196 ][ 50 ],
   alphaCSR[ 196 ][ 51 ],
   alphaCSR[ 196 ][ 52 ],
   alphaCSR[ 196 ][ 53 ],
   alphaCSR[ 196 ][ 54 ],
   alphaCSR[ 196 ][ 55 ],
   alphaCSR[ 196 ][ 56 ],
   alphaCSR[ 196 ][ 57 ],
   alphaCSR[ 196 ][ 58 ],
   alphaCSR[ 196 ][ 59 ],
   alphaCSR[ 196 ][ 60 ],
   alphaCSR[ 196 ][ 61 ],
   alphaCSR[ 196 ][ 62 ],
   alphaCSR[ 196 ][ 63 ],
   alphaCSR[ 196 ][ 64 ],
   alphaCSR[ 196 ][ 65 ],
   alphaCSR[ 196 ][ 66 ],
   alphaCSR[ 196 ][ 67 ],
   alphaCSR[ 196 ][ 68 ],
   alphaCSR[ 196 ][ 69 ],
   alphaCSR[ 196 ][ 70 ],
   alphaCSR[ 196 ][ 71 ],
   alphaCSR[ 196 ][ 72 ],
   alphaCSR[ 196 ][ 73 ],
   alphaCSR[ 196 ][ 74 ],
   alphaCSR[ 196 ][ 75 ],
   alphaCSR[ 196 ][ 76 ],
   alphaCSR[ 196 ][ 77 ],
   alphaCSR[ 196 ][ 78 ],
   alphaCSR[ 196 ][ 79 ],
   alphaCSR[ 196 ][ 80 ],
   alphaCSR[ 196 ][ 81 ],
   alphaCSR[ 196 ][ 82 ],
   alphaCSR[ 196 ][ 83 ],
   alphaCSR[ 196 ][ 84 ],
   alphaCSR[ 196 ][ 85 ],
   alphaCSR[ 196 ][ 86 ],
   alphaCSR[ 196 ][ 87 ],
   alphaCSR[ 196 ][ 88 ],
   alphaCSR[ 196 ][ 89 ],
   alphaCSR[ 196 ][ 90 ],
   alphaCSR[ 196 ][ 91 ],
   alphaCSR[ 196 ][ 92 ],
   alphaCSR[ 196 ][ 93 ],
   alphaCSR[ 196 ][ 94 ],
   alphaCSR[ 196 ][ 95 ],
   alphaCSR[ 196 ][ 96 ],
   alphaCSR[ 196 ][ 97 ],
   alphaCSR[ 196 ][ 98 ],
   alphaCSR[ 196 ][ 99 ],
   alphaCSR[ 196 ][ 100 ],
   alphaCSR[ 196 ][ 101 ],
   alphaCSR[ 196 ][ 102 ],
   alphaCSR[ 196 ][ 103 ],
   alphaCSR[ 196 ][ 104 ],
   alphaCSR[ 196 ][ 105 ],
   alphaCSR[ 196 ][ 106 ],
   alphaCSR[ 196 ][ 107 ],
   alphaCSR[ 196 ][ 108 ],
   alphaCSR[ 196 ][ 109 ],
   alphaCSR[ 196 ][ 110 ],
   alphaCSR[ 196 ][ 111 ],
   alphaCSR[ 196 ][ 112 ],
   alphaCSR[ 196 ][ 113 ],
   alphaCSR[ 196 ][ 114 ],
   alphaCSR[ 196 ][ 115 ],
   alphaCSR[ 196 ][ 116 ],
   alphaCSR[ 196 ][ 117 ],
   alphaCSR[ 196 ][ 118 ],
   alphaCSR[ 196 ][ 119 ],
   alphaCSR[ 196 ][ 120 ],
   alphaCSR[ 196 ][ 121 ],
   alphaCSR[ 196 ][ 122 ],
   alphaCSR[ 196 ][ 123 ],
   alphaCSR[ 196 ][ 124 ],
   alphaCSR[ 196 ][ 125 ],
   alphaCSR[ 196 ][ 126 ],
   alphaCSR[ 196 ][ 127 ],
   alphaCSR[ 196 ][ 128 ],
   alphaCSR[ 196 ][ 129 ],
   alphaCSR[ 196 ][ 130 ],
   alphaCSR[ 196 ][ 131 ],
   alphaCSR[ 196 ][ 132 ],
   alphaCSR[ 196 ][ 133 ],
   alphaCSR[ 196 ][ 134 ],
   alphaCSR[ 196 ][ 135 ],
   alphaCSR[ 196 ][ 136 ],
   alphaCSR[ 196 ][ 137 ],
   alphaCSR[ 196 ][ 138 ],
   alphaCSR[ 196 ][ 139 ],
   alphaCSR[ 196 ][ 140 ],
   alphaCSR[ 196 ][ 141 ],
   alphaCSR[ 196 ][ 142 ],
   alphaCSR[ 196 ][ 143 ],
   alphaCSR[ 196 ][ 144 ],
   alphaCSR[ 196 ][ 145 ],
   alphaCSR[ 196 ][ 146 ],
   alphaCSR[ 196 ][ 147 ],
   alphaCSR[ 196 ][ 148 ],
   alphaCSR[ 196 ][ 149 ],
   alphaCSR[ 196 ][ 150 ],
   alphaCSR[ 196 ][ 151 ],
   alphaCSR[ 196 ][ 152 ],
   alphaCSR[ 196 ][ 153 ],
   alphaCSR[ 196 ][ 154 ],
   alphaCSR[ 196 ][ 155 ],
   alphaCSR[ 196 ][ 156 ],
   alphaCSR[ 196 ][ 157 ],
   alphaCSR[ 196 ][ 158 ],
   alphaCSR[ 196 ][ 159 ],
   alphaCSR[ 196 ][ 160 ],
   alphaCSR[ 196 ][ 161 ],
   alphaCSR[ 196 ][ 162 ],
   alphaCSR[ 196 ][ 163 ],
   alphaCSR[ 196 ][ 164 ],
   alphaCSR[ 196 ][ 165 ],
   alphaCSR[ 196 ][ 166 ],
   alphaCSR[ 196 ][ 167 ],
   alphaCSR[ 196 ][ 168 ],
   alphaCSR[ 196 ][ 169 ],
   alphaCSR[ 196 ][ 170 ],
   alphaCSR[ 196 ][ 171 ],
   alphaCSR[ 196 ][ 172 ],
   alphaCSR[ 196 ][ 173 ],
   alphaCSR[ 196 ][ 174 ],
   alphaCSR[ 196 ][ 175 ],
   alphaCSR[ 196 ][ 176 ],
   alphaCSR[ 196 ][ 177 ],
   alphaCSR[ 196 ][ 178 ],
   alphaCSR[ 196 ][ 179 ],
   alphaCSR[ 196 ][ 180 ],
   alphaCSR[ 196 ][ 181 ],
   alphaCSR[ 196 ][ 182 ],
   alphaCSR[ 196 ][ 183 ],
   alphaCSR[ 196 ][ 184 ],
   alphaCSR[ 196 ][ 185 ],
   alphaCSR[ 196 ][ 186 ],
   alphaCSR[ 196 ][ 187 ],
   alphaCSR[ 196 ][ 188 ],
   alphaCSR[ 196 ][ 189 ],
   alphaCSR[ 196 ][ 190 ],
   alphaCSR[ 196 ][ 191 ],
   alphaCSR[ 196 ][ 192 ],
   alphaCSR[ 196 ][ 193 ],
   alphaCSR[ 196 ][ 194 ],
   alphaCSR[ 196 ][ 195 ],
   alphaCSR[ 196 ][ 196 ],
   alphaCSR[ 196 ][ 197 ],
   alphaCSR[ 196 ][ 198 ],
   alphaCSR[ 196 ][ 199 ],
   alphaCSR[ 196 ][ 200 ],
   alphaCSR[ 196 ][ 201 ],
   alphaCSR[ 196 ][ 202 ],
   alphaCSR[ 196 ][ 203 ],
   alphaCSR[ 196 ][ 204 ],
   alphaCSR[ 196 ][ 205 ],
   alphaCSR[ 196 ][ 206 ],
   alphaCSR[ 196 ][ 207 ],
   alphaCSR[ 196 ][ 208 ],
   alphaCSR[ 196 ][ 209 ],
   alphaCSR[ 196 ][ 210 ],
   alphaCSR[ 196 ][ 211 ],
   alphaCSR[ 196 ][ 212 ],
   alphaCSR[ 196 ][ 213 ],
   alphaCSR[ 196 ][ 214 ],
   alphaCSR[ 196 ][ 215 ],
   alphaCSR[ 196 ][ 216 ],
   alphaCSR[ 196 ][ 217 ],
   alphaCSR[ 196 ][ 218 ],
   alphaCSR[ 196 ][ 219 ],
   alphaCSR[ 196 ][ 220 ],
   alphaCSR[ 196 ][ 221 ],
   alphaCSR[ 196 ][ 222 ],
   alphaCSR[ 196 ][ 223 ],
   alphaCSR[ 196 ][ 224 ],
   alphaCSR[ 196 ][ 225 ],
   alphaCSR[ 196 ][ 226 ],
   alphaCSR[ 196 ][ 227 ],
   alphaCSR[ 196 ][ 228 ],
   alphaCSR[ 196 ][ 229 ],
   alphaCSR[ 196 ][ 230 ],
   alphaCSR[ 196 ][ 231 ],
   alphaCSR[ 196 ][ 232 ],
   alphaCSR[ 196 ][ 233 ],
   alphaCSR[ 196 ][ 234 ],
   alphaCSR[ 196 ][ 235 ],
   alphaCSR[ 196 ][ 236 ],
   alphaCSR[ 196 ][ 237 ],
   alphaCSR[ 196 ][ 238 ],
   alphaCSR[ 196 ][ 239 ],
   alphaCSR[ 196 ][ 240 ],
   alphaCSR[ 196 ][ 241 ],
   alphaCSR[ 196 ][ 242 ],
   alphaCSR[ 196 ][ 243 ],
   alphaCSR[ 196 ][ 244 ],
   alphaCSR[ 196 ][ 245 ],
   alphaCSR[ 196 ][ 246 ],
   alphaCSR[ 196 ][ 247 ],
   alphaCSR[ 196 ][ 248 ],
   alphaCSR[ 196 ][ 249 ],
   alphaCSR[ 196 ][ 250 ],
   alphaCSR[ 196 ][ 251 ],
   alphaCSR[ 196 ][ 252 ],
   alphaCSR[ 196 ][ 253 ],
   alphaCSR[ 196 ][ 254 ],
   alphaCSR[ 196 ][ 255 ],
   alphaCSR[ 196 ][ 256 ],
   alphaCSR[ 196 ][ 257 ],
   alphaCSR[ 196 ][ 258 ],
   alphaCSR[ 196 ][ 259 ],
   alphaCSR[ 196 ][ 260 ],
   alphaCSR[ 196 ][ 261 ],
   alphaCSR[ 196 ][ 262 ],
   alphaCSR[ 196 ][ 263 ],
   alphaCSR[ 196 ][ 264 ],
   alphaCSR[ 196 ][ 265 ],
   alphaCSR[ 196 ][ 266 ],
   alphaCSR[ 196 ][ 267 ],
   alphaCSR[ 196 ][ 268 ],
   alphaCSR[ 196 ][ 269 ],
   alphaCSR[ 196 ][ 270 ],
   alphaCSR[ 196 ][ 271 ],
   alphaCSR[ 196 ][ 272 ],
   alphaCSR[ 196 ][ 273 ],
   alphaCSR[ 196 ][ 274 ],
   alphaCSR[ 196 ][ 275 ],
   alphaCSR[ 196 ][ 276 ],
   alphaCSR[ 196 ][ 277 ],
   alphaCSR[ 196 ][ 278 ],
   alphaCSR[ 196 ][ 279 ],
   alphaCSR[ 196 ][ 280 ],
   alphaCSR[ 196 ][ 281 ],
   alphaCSR[ 196 ][ 282 ],
   alphaCSR[ 196 ][ 283 ],
   alphaCSR[ 196 ][ 284 ],
   alphaCSR[ 196 ][ 285 ],
   alphaCSR[ 196 ][ 286 ],
   alphaCSR[ 196 ][ 287 ],
   alphaCSR[ 196 ][ 288 ],
   alphaCSR[ 196 ][ 289 ],
   alphaCSR[ 196 ][ 290 ],
   alphaCSR[ 196 ][ 291 ],
   alphaCSR[ 196 ][ 292 ],
   alphaCSR[ 196 ][ 293 ],
   alphaCSR[ 196 ][ 294 ],
   alphaCSR[ 196 ][ 295 ],
   alphaCSR[ 196 ][ 296 ],
   alphaCSR[ 196 ][ 297 ],
   alphaCSR[ 196 ][ 298 ],
   alphaCSR[ 196 ][ 299 ],
   alphaCSR[ 196 ][ 300 ],
   alphaCSR[ 196 ][ 301 ],
   alphaCSR[ 196 ][ 302 ],
   alphaCSR[ 196 ][ 303 ],
   alphaCSR[ 196 ][ 304 ],
   alphaCSR[ 196 ][ 305 ],
   alphaCSR[ 196 ][ 306 ],
   alphaCSR[ 196 ][ 307 ],
   alphaCSR[ 196 ][ 308 ],
   alphaCSR[ 196 ][ 309 ],
   alphaCSR[ 196 ][ 310 ],
   alphaCSR[ 196 ][ 311 ],
   alphaCSR[ 196 ][ 312 ],
   alphaCSR[ 196 ][ 313 ],
   alphaCSR[ 196 ][ 314 ],
   alphaCSR[ 196 ][ 315 ],
   alphaCSR[ 196 ][ 316 ],
   alphaCSR[ 196 ][ 317 ],
   alphaCSR[ 196 ][ 318 ],
   alphaCSR[ 196 ][ 319 ],
   alphaCSR[ 196 ][ 320 ],
   alphaCSR[ 196 ][ 321 ],
   alphaCSR[ 196 ][ 322 ],
   alphaCSR[ 196 ][ 323 ],
   alphaCSR[ 196 ][ 324 ],
   alphaCSR[ 196 ][ 325 ],
   alphaCSR[ 196 ][ 326 ],
   alphaCSR[ 196 ][ 327 ],
   alphaCSR[ 196 ][ 328 ],
   alphaCSR[ 196 ][ 329 ],
   alphaCSR[ 196 ][ 330 ],
   alphaCSR[ 196 ][ 331 ],
   alphaCSR[ 196 ][ 332 ],
   alphaCSR[ 196 ][ 333 ],
   alphaCSR[ 196 ][ 334 ],
   alphaCSR[ 196 ][ 335 ],
   alphaCSR[ 196 ][ 336 ],
   alphaCSR[ 196 ][ 337 ],
   alphaCSR[ 196 ][ 338 ],
   alphaCSR[ 196 ][ 339 ],
   alphaCSR[ 196 ][ 340 ],
   alphaCSR[ 196 ][ 341 ],
   alphaCSR[ 196 ][ 342 ],
   alphaCSR[ 196 ][ 343 ],
   alphaCSR[ 196 ][ 344 ],
   alphaCSR[ 196 ][ 345 ],
   alphaCSR[ 196 ][ 346 ],
   alphaCSR[ 196 ][ 347 ],
   alphaCSR[ 196 ][ 348 ],
   alphaCSR[ 196 ][ 349 ],
   alphaCSR[ 196 ][ 350 ],
   alphaCSR[ 196 ][ 351 ],
   alphaCSR[ 196 ][ 352 ],
   alphaCSR[ 196 ][ 353 ],
   alphaCSR[ 196 ][ 354 ],
   alphaCSR[ 196 ][ 355 ],
   alphaCSR[ 196 ][ 356 ],
   alphaCSR[ 196 ][ 357 ],
   alphaCSR[ 196 ][ 358 ],
   alphaCSR[ 196 ][ 359 ],
   alphaCSR[ 196 ][ 360 ],
   alphaCSR[ 196 ][ 361 ],
   alphaCSR[ 196 ][ 362 ],
   alphaCSR[ 196 ][ 363 ],
   alphaCSR[ 196 ][ 364 ],
   alphaCSR[ 196 ][ 365 ],
   alphaCSR[ 196 ][ 366 ],
   alphaCSR[ 196 ][ 367 ],
   alphaCSR[ 196 ][ 368 ],
   alphaCSR[ 196 ][ 369 ],
   alphaCSR[ 196 ][ 370 ],
   alphaCSR[ 196 ][ 371 ],
   alphaCSR[ 196 ][ 372 ],
   alphaCSR[ 196 ][ 373 ],
   alphaCSR[ 196 ][ 374 ],
   alphaCSR[ 196 ][ 375 ],
   alphaCSR[ 196 ][ 376 ],
   alphaCSR[ 196 ][ 377 ],
   alphaCSR[ 196 ][ 378 ],
   alphaCSR[ 196 ][ 379 ],
   alphaCSR[ 196 ][ 380 ],
   alphaCSR[ 196 ][ 381 ],
   alphaCSR[ 196 ][ 382 ],
   alphaCSR[ 196 ][ 383 ],
   alphaCSR[ 197 ][ 0 ],
   alphaCSR[ 197 ][ 1 ],
   alphaCSR[ 197 ][ 2 ],
   alphaCSR[ 197 ][ 3 ],
   alphaCSR[ 197 ][ 4 ],
   alphaCSR[ 197 ][ 5 ],
   alphaCSR[ 197 ][ 6 ],
   alphaCSR[ 197 ][ 7 ],
   alphaCSR[ 197 ][ 8 ],
   alphaCSR[ 197 ][ 9 ],
   alphaCSR[ 197 ][ 10 ],
   alphaCSR[ 197 ][ 11 ],
   alphaCSR[ 197 ][ 12 ],
   alphaCSR[ 197 ][ 13 ],
   alphaCSR[ 197 ][ 14 ],
   alphaCSR[ 197 ][ 15 ],
   alphaCSR[ 197 ][ 16 ],
   alphaCSR[ 197 ][ 17 ],
   alphaCSR[ 197 ][ 18 ],
   alphaCSR[ 197 ][ 19 ],
   alphaCSR[ 197 ][ 20 ],
   alphaCSR[ 197 ][ 21 ],
   alphaCSR[ 197 ][ 22 ],
   alphaCSR[ 197 ][ 23 ],
   alphaCSR[ 197 ][ 24 ],
   alphaCSR[ 197 ][ 25 ],
   alphaCSR[ 197 ][ 26 ],
   alphaCSR[ 197 ][ 27 ],
   alphaCSR[ 197 ][ 28 ],
   alphaCSR[ 197 ][ 29 ],
   alphaCSR[ 197 ][ 30 ],
   alphaCSR[ 197 ][ 31 ],
   alphaCSR[ 197 ][ 32 ],
   alphaCSR[ 197 ][ 33 ],
   alphaCSR[ 197 ][ 34 ],
   alphaCSR[ 197 ][ 35 ],
   alphaCSR[ 197 ][ 36 ],
   alphaCSR[ 197 ][ 37 ],
   alphaCSR[ 197 ][ 38 ],
   alphaCSR[ 197 ][ 39 ],
   alphaCSR[ 197 ][ 40 ],
   alphaCSR[ 197 ][ 41 ],
   alphaCSR[ 197 ][ 42 ],
   alphaCSR[ 197 ][ 43 ],
   alphaCSR[ 197 ][ 44 ],
   alphaCSR[ 197 ][ 45 ],
   alphaCSR[ 197 ][ 46 ],
   alphaCSR[ 197 ][ 47 ],
   alphaCSR[ 197 ][ 48 ],
   alphaCSR[ 197 ][ 49 ],
   alphaCSR[ 197 ][ 50 ],
   alphaCSR[ 197 ][ 51 ],
   alphaCSR[ 197 ][ 52 ],
   alphaCSR[ 197 ][ 53 ],
   alphaCSR[ 197 ][ 54 ],
   alphaCSR[ 197 ][ 55 ],
   alphaCSR[ 197 ][ 56 ],
   alphaCSR[ 197 ][ 57 ],
   alphaCSR[ 197 ][ 58 ],
   alphaCSR[ 197 ][ 59 ],
   alphaCSR[ 197 ][ 60 ],
   alphaCSR[ 197 ][ 61 ],
   alphaCSR[ 197 ][ 62 ],
   alphaCSR[ 197 ][ 63 ],
   alphaCSR[ 197 ][ 64 ],
   alphaCSR[ 197 ][ 65 ],
   alphaCSR[ 197 ][ 66 ],
   alphaCSR[ 197 ][ 67 ],
   alphaCSR[ 197 ][ 68 ],
   alphaCSR[ 197 ][ 69 ],
   alphaCSR[ 197 ][ 70 ],
   alphaCSR[ 197 ][ 71 ],
   alphaCSR[ 197 ][ 72 ],
   alphaCSR[ 197 ][ 73 ],
   alphaCSR[ 197 ][ 74 ],
   alphaCSR[ 197 ][ 75 ],
   alphaCSR[ 197 ][ 76 ],
   alphaCSR[ 197 ][ 77 ],
   alphaCSR[ 197 ][ 78 ],
   alphaCSR[ 197 ][ 79 ],
   alphaCSR[ 197 ][ 80 ],
   alphaCSR[ 197 ][ 81 ],
   alphaCSR[ 197 ][ 82 ],
   alphaCSR[ 197 ][ 83 ],
   alphaCSR[ 197 ][ 84 ],
   alphaCSR[ 197 ][ 85 ],
   alphaCSR[ 197 ][ 86 ],
   alphaCSR[ 197 ][ 87 ],
   alphaCSR[ 197 ][ 88 ],
   alphaCSR[ 197 ][ 89 ],
   alphaCSR[ 197 ][ 90 ],
   alphaCSR[ 197 ][ 91 ],
   alphaCSR[ 197 ][ 92 ],
   alphaCSR[ 197 ][ 93 ],
   alphaCSR[ 197 ][ 94 ],
   alphaCSR[ 197 ][ 95 ],
   alphaCSR[ 197 ][ 96 ],
   alphaCSR[ 197 ][ 97 ],
   alphaCSR[ 197 ][ 98 ],
   alphaCSR[ 197 ][ 99 ],
   alphaCSR[ 197 ][ 100 ],
   alphaCSR[ 197 ][ 101 ],
   alphaCSR[ 197 ][ 102 ],
   alphaCSR[ 197 ][ 103 ],
   alphaCSR[ 197 ][ 104 ],
   alphaCSR[ 197 ][ 105 ],
   alphaCSR[ 197 ][ 106 ],
   alphaCSR[ 197 ][ 107 ],
   alphaCSR[ 197 ][ 108 ],
   alphaCSR[ 197 ][ 109 ],
   alphaCSR[ 197 ][ 110 ],
   alphaCSR[ 197 ][ 111 ],
   alphaCSR[ 197 ][ 112 ],
   alphaCSR[ 197 ][ 113 ],
   alphaCSR[ 197 ][ 114 ],
   alphaCSR[ 197 ][ 115 ],
   alphaCSR[ 197 ][ 116 ],
   alphaCSR[ 197 ][ 117 ],
   alphaCSR[ 197 ][ 118 ],
   alphaCSR[ 197 ][ 119 ],
   alphaCSR[ 197 ][ 120 ],
   alphaCSR[ 197 ][ 121 ],
   alphaCSR[ 197 ][ 122 ],
   alphaCSR[ 197 ][ 123 ],
   alphaCSR[ 197 ][ 124 ],
   alphaCSR[ 197 ][ 125 ],
   alphaCSR[ 197 ][ 126 ],
   alphaCSR[ 197 ][ 127 ],
   alphaCSR[ 197 ][ 128 ],
   alphaCSR[ 197 ][ 129 ],
   alphaCSR[ 197 ][ 130 ],
   alphaCSR[ 197 ][ 131 ],
   alphaCSR[ 197 ][ 132 ],
   alphaCSR[ 197 ][ 133 ],
   alphaCSR[ 197 ][ 134 ],
   alphaCSR[ 197 ][ 135 ],
   alphaCSR[ 197 ][ 136 ],
   alphaCSR[ 197 ][ 137 ],
   alphaCSR[ 197 ][ 138 ],
   alphaCSR[ 197 ][ 139 ],
   alphaCSR[ 197 ][ 140 ],
   alphaCSR[ 197 ][ 141 ],
   alphaCSR[ 197 ][ 142 ],
   alphaCSR[ 197 ][ 143 ],
   alphaCSR[ 197 ][ 144 ],
   alphaCSR[ 197 ][ 145 ],
   alphaCSR[ 197 ][ 146 ],
   alphaCSR[ 197 ][ 147 ],
   alphaCSR[ 197 ][ 148 ],
   alphaCSR[ 197 ][ 149 ],
   alphaCSR[ 197 ][ 150 ],
   alphaCSR[ 197 ][ 151 ],
   alphaCSR[ 197 ][ 152 ],
   alphaCSR[ 197 ][ 153 ],
   alphaCSR[ 197 ][ 154 ],
   alphaCSR[ 197 ][ 155 ],
   alphaCSR[ 197 ][ 156 ],
   alphaCSR[ 197 ][ 157 ],
   alphaCSR[ 197 ][ 158 ],
   alphaCSR[ 197 ][ 159 ],
   alphaCSR[ 197 ][ 160 ],
   alphaCSR[ 197 ][ 161 ],
   alphaCSR[ 197 ][ 162 ],
   alphaCSR[ 197 ][ 163 ],
   alphaCSR[ 197 ][ 164 ],
   alphaCSR[ 197 ][ 165 ],
   alphaCSR[ 197 ][ 166 ],
   alphaCSR[ 197 ][ 167 ],
   alphaCSR[ 197 ][ 168 ],
   alphaCSR[ 197 ][ 169 ],
   alphaCSR[ 197 ][ 170 ],
   alphaCSR[ 197 ][ 171 ],
   alphaCSR[ 197 ][ 172 ],
   alphaCSR[ 197 ][ 173 ],
   alphaCSR[ 197 ][ 174 ],
   alphaCSR[ 197 ][ 175 ],
   alphaCSR[ 197 ][ 176 ],
   alphaCSR[ 197 ][ 177 ],
   alphaCSR[ 197 ][ 178 ],
   alphaCSR[ 197 ][ 179 ],
   alphaCSR[ 197 ][ 180 ],
   alphaCSR[ 197 ][ 181 ],
   alphaCSR[ 197 ][ 182 ],
   alphaCSR[ 197 ][ 183 ],
   alphaCSR[ 197 ][ 184 ],
   alphaCSR[ 197 ][ 185 ],
   alphaCSR[ 197 ][ 186 ],
   alphaCSR[ 197 ][ 187 ],
   alphaCSR[ 197 ][ 188 ],
   alphaCSR[ 197 ][ 189 ],
   alphaCSR[ 197 ][ 190 ],
   alphaCSR[ 197 ][ 191 ],
   alphaCSR[ 197 ][ 192 ],
   alphaCSR[ 197 ][ 193 ],
   alphaCSR[ 197 ][ 194 ],
   alphaCSR[ 197 ][ 195 ],
   alphaCSR[ 197 ][ 196 ],
   alphaCSR[ 197 ][ 197 ],
   alphaCSR[ 197 ][ 198 ],
   alphaCSR[ 197 ][ 199 ],
   alphaCSR[ 197 ][ 200 ],
   alphaCSR[ 197 ][ 201 ],
   alphaCSR[ 197 ][ 202 ],
   alphaCSR[ 197 ][ 203 ],
   alphaCSR[ 197 ][ 204 ],
   alphaCSR[ 197 ][ 205 ],
   alphaCSR[ 197 ][ 206 ],
   alphaCSR[ 197 ][ 207 ],
   alphaCSR[ 197 ][ 208 ],
   alphaCSR[ 197 ][ 209 ],
   alphaCSR[ 197 ][ 210 ],
   alphaCSR[ 197 ][ 211 ],
   alphaCSR[ 197 ][ 212 ],
   alphaCSR[ 197 ][ 213 ],
   alphaCSR[ 197 ][ 214 ],
   alphaCSR[ 197 ][ 215 ],
   alphaCSR[ 197 ][ 216 ],
   alphaCSR[ 197 ][ 217 ],
   alphaCSR[ 197 ][ 218 ],
   alphaCSR[ 197 ][ 219 ],
   alphaCSR[ 197 ][ 220 ],
   alphaCSR[ 197 ][ 221 ],
   alphaCSR[ 197 ][ 222 ],
   alphaCSR[ 197 ][ 223 ],
   alphaCSR[ 197 ][ 224 ],
   alphaCSR[ 197 ][ 225 ],
   alphaCSR[ 197 ][ 226 ],
   alphaCSR[ 197 ][ 227 ],
   alphaCSR[ 197 ][ 228 ],
   alphaCSR[ 197 ][ 229 ],
   alphaCSR[ 197 ][ 230 ],
   alphaCSR[ 197 ][ 231 ],
   alphaCSR[ 197 ][ 232 ],
   alphaCSR[ 197 ][ 233 ],
   alphaCSR[ 197 ][ 234 ],
   alphaCSR[ 197 ][ 235 ],
   alphaCSR[ 197 ][ 236 ],
   alphaCSR[ 197 ][ 237 ],
   alphaCSR[ 197 ][ 238 ],
   alphaCSR[ 197 ][ 239 ],
   alphaCSR[ 197 ][ 240 ],
   alphaCSR[ 197 ][ 241 ],
   alphaCSR[ 197 ][ 242 ],
   alphaCSR[ 197 ][ 243 ],
   alphaCSR[ 197 ][ 244 ],
   alphaCSR[ 197 ][ 245 ],
   alphaCSR[ 197 ][ 246 ],
   alphaCSR[ 197 ][ 247 ],
   alphaCSR[ 197 ][ 248 ],
   alphaCSR[ 197 ][ 249 ],
   alphaCSR[ 197 ][ 250 ],
   alphaCSR[ 197 ][ 251 ],
   alphaCSR[ 197 ][ 252 ],
   alphaCSR[ 197 ][ 253 ],
   alphaCSR[ 197 ][ 254 ],
   alphaCSR[ 197 ][ 255 ],
   alphaCSR[ 197 ][ 256 ],
   alphaCSR[ 197 ][ 257 ],
   alphaCSR[ 197 ][ 258 ],
   alphaCSR[ 197 ][ 259 ],
   alphaCSR[ 197 ][ 260 ],
   alphaCSR[ 197 ][ 261 ],
   alphaCSR[ 197 ][ 262 ],
   alphaCSR[ 197 ][ 263 ],
   alphaCSR[ 197 ][ 264 ],
   alphaCSR[ 197 ][ 265 ],
   alphaCSR[ 197 ][ 266 ],
   alphaCSR[ 197 ][ 267 ],
   alphaCSR[ 197 ][ 268 ],
   alphaCSR[ 197 ][ 269 ],
   alphaCSR[ 197 ][ 270 ],
   alphaCSR[ 197 ][ 271 ],
   alphaCSR[ 197 ][ 272 ],
   alphaCSR[ 197 ][ 273 ],
   alphaCSR[ 197 ][ 274 ],
   alphaCSR[ 197 ][ 275 ],
   alphaCSR[ 197 ][ 276 ],
   alphaCSR[ 197 ][ 277 ],
   alphaCSR[ 197 ][ 278 ],
   alphaCSR[ 197 ][ 279 ],
   alphaCSR[ 197 ][ 280 ],
   alphaCSR[ 197 ][ 281 ],
   alphaCSR[ 197 ][ 282 ],
   alphaCSR[ 197 ][ 283 ],
   alphaCSR[ 197 ][ 284 ],
   alphaCSR[ 197 ][ 285 ],
   alphaCSR[ 197 ][ 286 ],
   alphaCSR[ 197 ][ 287 ],
   alphaCSR[ 197 ][ 288 ],
   alphaCSR[ 197 ][ 289 ],
   alphaCSR[ 197 ][ 290 ],
   alphaCSR[ 197 ][ 291 ],
   alphaCSR[ 197 ][ 292 ],
   alphaCSR[ 197 ][ 293 ],
   alphaCSR[ 197 ][ 294 ],
   alphaCSR[ 197 ][ 295 ],
   alphaCSR[ 197 ][ 296 ],
   alphaCSR[ 197 ][ 297 ],
   alphaCSR[ 197 ][ 298 ],
   alphaCSR[ 197 ][ 299 ],
   alphaCSR[ 197 ][ 300 ],
   alphaCSR[ 197 ][ 301 ],
   alphaCSR[ 197 ][ 302 ],
   alphaCSR[ 197 ][ 303 ],
   alphaCSR[ 197 ][ 304 ],
   alphaCSR[ 197 ][ 305 ],
   alphaCSR[ 197 ][ 306 ],
   alphaCSR[ 197 ][ 307 ],
   alphaCSR[ 197 ][ 308 ],
   alphaCSR[ 197 ][ 309 ],
   alphaCSR[ 197 ][ 310 ],
   alphaCSR[ 197 ][ 311 ],
   alphaCSR[ 197 ][ 312 ],
   alphaCSR[ 197 ][ 313 ],
   alphaCSR[ 197 ][ 314 ],
   alphaCSR[ 197 ][ 315 ],
   alphaCSR[ 197 ][ 316 ],
   alphaCSR[ 197 ][ 317 ],
   alphaCSR[ 197 ][ 318 ],
   alphaCSR[ 197 ][ 319 ],
   alphaCSR[ 197 ][ 320 ],
   alphaCSR[ 197 ][ 321 ],
   alphaCSR[ 197 ][ 322 ],
   alphaCSR[ 197 ][ 323 ],
   alphaCSR[ 197 ][ 324 ],
   alphaCSR[ 197 ][ 325 ],
   alphaCSR[ 197 ][ 326 ],
   alphaCSR[ 197 ][ 327 ],
   alphaCSR[ 197 ][ 328 ],
   alphaCSR[ 197 ][ 329 ],
   alphaCSR[ 197 ][ 330 ],
   alphaCSR[ 197 ][ 331 ],
   alphaCSR[ 197 ][ 332 ],
   alphaCSR[ 197 ][ 333 ],
   alphaCSR[ 197 ][ 334 ],
   alphaCSR[ 197 ][ 335 ],
   alphaCSR[ 197 ][ 336 ],
   alphaCSR[ 197 ][ 337 ],
   alphaCSR[ 197 ][ 338 ],
   alphaCSR[ 197 ][ 339 ],
   alphaCSR[ 197 ][ 340 ],
   alphaCSR[ 197 ][ 341 ],
   alphaCSR[ 197 ][ 342 ],
   alphaCSR[ 197 ][ 343 ],
   alphaCSR[ 197 ][ 344 ],
   alphaCSR[ 197 ][ 345 ],
   alphaCSR[ 197 ][ 346 ],
   alphaCSR[ 197 ][ 347 ],
   alphaCSR[ 197 ][ 348 ],
   alphaCSR[ 197 ][ 349 ],
   alphaCSR[ 197 ][ 350 ],
   alphaCSR[ 197 ][ 351 ],
   alphaCSR[ 197 ][ 352 ],
   alphaCSR[ 197 ][ 353 ],
   alphaCSR[ 197 ][ 354 ],
   alphaCSR[ 197 ][ 355 ],
   alphaCSR[ 197 ][ 356 ],
   alphaCSR[ 197 ][ 357 ],
   alphaCSR[ 197 ][ 358 ],
   alphaCSR[ 197 ][ 359 ],
   alphaCSR[ 197 ][ 360 ],
   alphaCSR[ 197 ][ 361 ],
   alphaCSR[ 197 ][ 362 ],
   alphaCSR[ 197 ][ 363 ],
   alphaCSR[ 197 ][ 364 ],
   alphaCSR[ 197 ][ 365 ],
   alphaCSR[ 197 ][ 366 ],
   alphaCSR[ 197 ][ 367 ],
   alphaCSR[ 197 ][ 368 ],
   alphaCSR[ 197 ][ 369 ],
   alphaCSR[ 197 ][ 370 ],
   alphaCSR[ 197 ][ 371 ],
   alphaCSR[ 197 ][ 372 ],
   alphaCSR[ 197 ][ 373 ],
   alphaCSR[ 197 ][ 374 ],
   alphaCSR[ 197 ][ 375 ],
   alphaCSR[ 197 ][ 376 ],
   alphaCSR[ 197 ][ 377 ],
   alphaCSR[ 197 ][ 378 ],
   alphaCSR[ 197 ][ 379 ],
   alphaCSR[ 197 ][ 380 ],
   alphaCSR[ 197 ][ 381 ],
   alphaCSR[ 197 ][ 382 ],
   alphaCSR[ 197 ][ 383 ],
   alphaCSR[ 198 ][ 0 ],
   alphaCSR[ 198 ][ 1 ],
   alphaCSR[ 198 ][ 2 ],
   alphaCSR[ 198 ][ 3 ],
   alphaCSR[ 198 ][ 4 ],
   alphaCSR[ 198 ][ 5 ],
   alphaCSR[ 198 ][ 6 ],
   alphaCSR[ 198 ][ 7 ],
   alphaCSR[ 198 ][ 8 ],
   alphaCSR[ 198 ][ 9 ],
   alphaCSR[ 198 ][ 10 ],
   alphaCSR[ 198 ][ 11 ],
   alphaCSR[ 198 ][ 12 ],
   alphaCSR[ 198 ][ 13 ],
   alphaCSR[ 198 ][ 14 ],
   alphaCSR[ 198 ][ 15 ],
   alphaCSR[ 198 ][ 16 ],
   alphaCSR[ 198 ][ 17 ],
   alphaCSR[ 198 ][ 18 ],
   alphaCSR[ 198 ][ 19 ],
   alphaCSR[ 198 ][ 20 ],
   alphaCSR[ 198 ][ 21 ],
   alphaCSR[ 198 ][ 22 ],
   alphaCSR[ 198 ][ 23 ],
   alphaCSR[ 198 ][ 24 ],
   alphaCSR[ 198 ][ 25 ],
   alphaCSR[ 198 ][ 26 ],
   alphaCSR[ 198 ][ 27 ],
   alphaCSR[ 198 ][ 28 ],
   alphaCSR[ 198 ][ 29 ],
   alphaCSR[ 198 ][ 30 ],
   alphaCSR[ 198 ][ 31 ],
   alphaCSR[ 198 ][ 32 ],
   alphaCSR[ 198 ][ 33 ],
   alphaCSR[ 198 ][ 34 ],
   alphaCSR[ 198 ][ 35 ],
   alphaCSR[ 198 ][ 36 ],
   alphaCSR[ 198 ][ 37 ],
   alphaCSR[ 198 ][ 38 ],
   alphaCSR[ 198 ][ 39 ],
   alphaCSR[ 198 ][ 40 ],
   alphaCSR[ 198 ][ 41 ],
   alphaCSR[ 198 ][ 42 ],
   alphaCSR[ 198 ][ 43 ],
   alphaCSR[ 198 ][ 44 ],
   alphaCSR[ 198 ][ 45 ],
   alphaCSR[ 198 ][ 46 ],
   alphaCSR[ 198 ][ 47 ],
   alphaCSR[ 198 ][ 48 ],
   alphaCSR[ 198 ][ 49 ],
   alphaCSR[ 198 ][ 50 ],
   alphaCSR[ 198 ][ 51 ],
   alphaCSR[ 198 ][ 52 ],
   alphaCSR[ 198 ][ 53 ],
   alphaCSR[ 198 ][ 54 ],
   alphaCSR[ 198 ][ 55 ],
   alphaCSR[ 198 ][ 56 ],
   alphaCSR[ 198 ][ 57 ],
   alphaCSR[ 198 ][ 58 ],
   alphaCSR[ 198 ][ 59 ],
   alphaCSR[ 198 ][ 60 ],
   alphaCSR[ 198 ][ 61 ],
   alphaCSR[ 198 ][ 62 ],
   alphaCSR[ 198 ][ 63 ],
   alphaCSR[ 198 ][ 64 ],
   alphaCSR[ 198 ][ 65 ],
   alphaCSR[ 198 ][ 66 ],
   alphaCSR[ 198 ][ 67 ],
   alphaCSR[ 198 ][ 68 ],
   alphaCSR[ 198 ][ 69 ],
   alphaCSR[ 198 ][ 70 ],
   alphaCSR[ 198 ][ 71 ],
   alphaCSR[ 198 ][ 72 ],
   alphaCSR[ 198 ][ 73 ],
   alphaCSR[ 198 ][ 74 ],
   alphaCSR[ 198 ][ 75 ],
   alphaCSR[ 198 ][ 76 ],
   alphaCSR[ 198 ][ 77 ],
   alphaCSR[ 198 ][ 78 ],
   alphaCSR[ 198 ][ 79 ],
   alphaCSR[ 198 ][ 80 ],
   alphaCSR[ 198 ][ 81 ],
   alphaCSR[ 198 ][ 82 ],
   alphaCSR[ 198 ][ 83 ],
   alphaCSR[ 198 ][ 84 ],
   alphaCSR[ 198 ][ 85 ],
   alphaCSR[ 198 ][ 86 ],
   alphaCSR[ 198 ][ 87 ],
   alphaCSR[ 198 ][ 88 ],
   alphaCSR[ 198 ][ 89 ],
   alphaCSR[ 198 ][ 90 ],
   alphaCSR[ 198 ][ 91 ],
   alphaCSR[ 198 ][ 92 ],
   alphaCSR[ 198 ][ 93 ],
   alphaCSR[ 198 ][ 94 ],
   alphaCSR[ 198 ][ 95 ],
   alphaCSR[ 198 ][ 96 ],
   alphaCSR[ 198 ][ 97 ],
   alphaCSR[ 198 ][ 98 ],
   alphaCSR[ 198 ][ 99 ],
   alphaCSR[ 198 ][ 100 ],
   alphaCSR[ 198 ][ 101 ],
   alphaCSR[ 198 ][ 102 ],
   alphaCSR[ 198 ][ 103 ],
   alphaCSR[ 198 ][ 104 ],
   alphaCSR[ 198 ][ 105 ],
   alphaCSR[ 198 ][ 106 ],
   alphaCSR[ 198 ][ 107 ],
   alphaCSR[ 198 ][ 108 ],
   alphaCSR[ 198 ][ 109 ],
   alphaCSR[ 198 ][ 110 ],
   alphaCSR[ 198 ][ 111 ],
   alphaCSR[ 198 ][ 112 ],
   alphaCSR[ 198 ][ 113 ],
   alphaCSR[ 198 ][ 114 ],
   alphaCSR[ 198 ][ 115 ],
   alphaCSR[ 198 ][ 116 ],
   alphaCSR[ 198 ][ 117 ],
   alphaCSR[ 198 ][ 118 ],
   alphaCSR[ 198 ][ 119 ],
   alphaCSR[ 198 ][ 120 ],
   alphaCSR[ 198 ][ 121 ],
   alphaCSR[ 198 ][ 122 ],
   alphaCSR[ 198 ][ 123 ],
   alphaCSR[ 198 ][ 124 ],
   alphaCSR[ 198 ][ 125 ],
   alphaCSR[ 198 ][ 126 ],
   alphaCSR[ 198 ][ 127 ],
   alphaCSR[ 198 ][ 128 ],
   alphaCSR[ 198 ][ 129 ],
   alphaCSR[ 198 ][ 130 ],
   alphaCSR[ 198 ][ 131 ],
   alphaCSR[ 198 ][ 132 ],
   alphaCSR[ 198 ][ 133 ],
   alphaCSR[ 198 ][ 134 ],
   alphaCSR[ 198 ][ 135 ],
   alphaCSR[ 198 ][ 136 ],
   alphaCSR[ 198 ][ 137 ],
   alphaCSR[ 198 ][ 138 ],
   alphaCSR[ 198 ][ 139 ],
   alphaCSR[ 198 ][ 140 ],
   alphaCSR[ 198 ][ 141 ],
   alphaCSR[ 198 ][ 142 ],
   alphaCSR[ 198 ][ 143 ],
   alphaCSR[ 198 ][ 144 ],
   alphaCSR[ 198 ][ 145 ],
   alphaCSR[ 198 ][ 146 ],
   alphaCSR[ 198 ][ 147 ],
   alphaCSR[ 198 ][ 148 ],
   alphaCSR[ 198 ][ 149 ],
   alphaCSR[ 198 ][ 150 ],
   alphaCSR[ 198 ][ 151 ],
   alphaCSR[ 198 ][ 152 ],
   alphaCSR[ 198 ][ 153 ],
   alphaCSR[ 198 ][ 154 ],
   alphaCSR[ 198 ][ 155 ],
   alphaCSR[ 198 ][ 156 ],
   alphaCSR[ 198 ][ 157 ],
   alphaCSR[ 198 ][ 158 ],
   alphaCSR[ 198 ][ 159 ],
   alphaCSR[ 198 ][ 160 ],
   alphaCSR[ 198 ][ 161 ],
   alphaCSR[ 198 ][ 162 ],
   alphaCSR[ 198 ][ 163 ],
   alphaCSR[ 198 ][ 164 ],
   alphaCSR[ 198 ][ 165 ],
   alphaCSR[ 198 ][ 166 ],
   alphaCSR[ 198 ][ 167 ],
   alphaCSR[ 198 ][ 168 ],
   alphaCSR[ 198 ][ 169 ],
   alphaCSR[ 198 ][ 170 ],
   alphaCSR[ 198 ][ 171 ],
   alphaCSR[ 198 ][ 172 ],
   alphaCSR[ 198 ][ 173 ],
   alphaCSR[ 198 ][ 174 ],
   alphaCSR[ 198 ][ 175 ],
   alphaCSR[ 198 ][ 176 ],
   alphaCSR[ 198 ][ 177 ],
   alphaCSR[ 198 ][ 178 ],
   alphaCSR[ 198 ][ 179 ],
   alphaCSR[ 198 ][ 180 ],
   alphaCSR[ 198 ][ 181 ],
   alphaCSR[ 198 ][ 182 ],
   alphaCSR[ 198 ][ 183 ],
   alphaCSR[ 198 ][ 184 ],
   alphaCSR[ 198 ][ 185 ],
   alphaCSR[ 198 ][ 186 ],
   alphaCSR[ 198 ][ 187 ],
   alphaCSR[ 198 ][ 188 ],
   alphaCSR[ 198 ][ 189 ],
   alphaCSR[ 198 ][ 190 ],
   alphaCSR[ 198 ][ 191 ],
   alphaCSR[ 198 ][ 192 ],
   alphaCSR[ 198 ][ 193 ],
   alphaCSR[ 198 ][ 194 ],
   alphaCSR[ 198 ][ 195 ],
   alphaCSR[ 198 ][ 196 ],
   alphaCSR[ 198 ][ 197 ],
   alphaCSR[ 198 ][ 198 ],
   alphaCSR[ 198 ][ 199 ],
   alphaCSR[ 198 ][ 200 ],
   alphaCSR[ 198 ][ 201 ],
   alphaCSR[ 198 ][ 202 ],
   alphaCSR[ 198 ][ 203 ],
   alphaCSR[ 198 ][ 204 ],
   alphaCSR[ 198 ][ 205 ],
   alphaCSR[ 198 ][ 206 ],
   alphaCSR[ 198 ][ 207 ],
   alphaCSR[ 198 ][ 208 ],
   alphaCSR[ 198 ][ 209 ],
   alphaCSR[ 198 ][ 210 ],
   alphaCSR[ 198 ][ 211 ],
   alphaCSR[ 198 ][ 212 ],
   alphaCSR[ 198 ][ 213 ],
   alphaCSR[ 198 ][ 214 ],
   alphaCSR[ 198 ][ 215 ],
   alphaCSR[ 198 ][ 216 ],
   alphaCSR[ 198 ][ 217 ],
   alphaCSR[ 198 ][ 218 ],
   alphaCSR[ 198 ][ 219 ],
   alphaCSR[ 198 ][ 220 ],
   alphaCSR[ 198 ][ 221 ],
   alphaCSR[ 198 ][ 222 ],
   alphaCSR[ 198 ][ 223 ],
   alphaCSR[ 198 ][ 224 ],
   alphaCSR[ 198 ][ 225 ],
   alphaCSR[ 198 ][ 226 ],
   alphaCSR[ 198 ][ 227 ],
   alphaCSR[ 198 ][ 228 ],
   alphaCSR[ 198 ][ 229 ],
   alphaCSR[ 198 ][ 230 ],
   alphaCSR[ 198 ][ 231 ],
   alphaCSR[ 198 ][ 232 ],
   alphaCSR[ 198 ][ 233 ],
   alphaCSR[ 198 ][ 234 ],
   alphaCSR[ 198 ][ 235 ],
   alphaCSR[ 198 ][ 236 ],
   alphaCSR[ 198 ][ 237 ],
   alphaCSR[ 198 ][ 238 ],
   alphaCSR[ 198 ][ 239 ],
   alphaCSR[ 198 ][ 240 ],
   alphaCSR[ 198 ][ 241 ],
   alphaCSR[ 198 ][ 242 ],
   alphaCSR[ 198 ][ 243 ],
   alphaCSR[ 198 ][ 244 ],
   alphaCSR[ 198 ][ 245 ],
   alphaCSR[ 198 ][ 246 ],
   alphaCSR[ 198 ][ 247 ],
   alphaCSR[ 198 ][ 248 ],
   alphaCSR[ 198 ][ 249 ],
   alphaCSR[ 198 ][ 250 ],
   alphaCSR[ 198 ][ 251 ],
   alphaCSR[ 198 ][ 252 ],
   alphaCSR[ 198 ][ 253 ],
   alphaCSR[ 198 ][ 254 ],
   alphaCSR[ 198 ][ 255 ],
   alphaCSR[ 198 ][ 256 ],
   alphaCSR[ 198 ][ 257 ],
   alphaCSR[ 198 ][ 258 ],
   alphaCSR[ 198 ][ 259 ],
   alphaCSR[ 198 ][ 260 ],
   alphaCSR[ 198 ][ 261 ],
   alphaCSR[ 198 ][ 262 ],
   alphaCSR[ 198 ][ 263 ],
   alphaCSR[ 198 ][ 264 ],
   alphaCSR[ 198 ][ 265 ],
   alphaCSR[ 198 ][ 266 ],
   alphaCSR[ 198 ][ 267 ],
   alphaCSR[ 198 ][ 268 ],
   alphaCSR[ 198 ][ 269 ],
   alphaCSR[ 198 ][ 270 ],
   alphaCSR[ 198 ][ 271 ],
   alphaCSR[ 198 ][ 272 ],
   alphaCSR[ 198 ][ 273 ],
   alphaCSR[ 198 ][ 274 ],
   alphaCSR[ 198 ][ 275 ],
   alphaCSR[ 198 ][ 276 ],
   alphaCSR[ 198 ][ 277 ],
   alphaCSR[ 198 ][ 278 ],
   alphaCSR[ 198 ][ 279 ],
   alphaCSR[ 198 ][ 280 ],
   alphaCSR[ 198 ][ 281 ],
   alphaCSR[ 198 ][ 282 ],
   alphaCSR[ 198 ][ 283 ],
   alphaCSR[ 198 ][ 284 ],
   alphaCSR[ 198 ][ 285 ],
   alphaCSR[ 198 ][ 286 ],
   alphaCSR[ 198 ][ 287 ],
   alphaCSR[ 198 ][ 288 ],
   alphaCSR[ 198 ][ 289 ],
   alphaCSR[ 198 ][ 290 ],
   alphaCSR[ 198 ][ 291 ],
   alphaCSR[ 198 ][ 292 ],
   alphaCSR[ 198 ][ 293 ],
   alphaCSR[ 198 ][ 294 ],
   alphaCSR[ 198 ][ 295 ],
   alphaCSR[ 198 ][ 296 ],
   alphaCSR[ 198 ][ 297 ],
   alphaCSR[ 198 ][ 298 ],
   alphaCSR[ 198 ][ 299 ],
   alphaCSR[ 198 ][ 300 ],
   alphaCSR[ 198 ][ 301 ],
   alphaCSR[ 198 ][ 302 ],
   alphaCSR[ 198 ][ 303 ],
   alphaCSR[ 198 ][ 304 ],
   alphaCSR[ 198 ][ 305 ],
   alphaCSR[ 198 ][ 306 ],
   alphaCSR[ 198 ][ 307 ],
   alphaCSR[ 198 ][ 308 ],
   alphaCSR[ 198 ][ 309 ],
   alphaCSR[ 198 ][ 310 ],
   alphaCSR[ 198 ][ 311 ],
   alphaCSR[ 198 ][ 312 ],
   alphaCSR[ 198 ][ 313 ],
   alphaCSR[ 198 ][ 314 ],
   alphaCSR[ 198 ][ 315 ],
   alphaCSR[ 198 ][ 316 ],
   alphaCSR[ 198 ][ 317 ],
   alphaCSR[ 198 ][ 318 ],
   alphaCSR[ 198 ][ 319 ],
   alphaCSR[ 198 ][ 320 ],
   alphaCSR[ 198 ][ 321 ],
   alphaCSR[ 198 ][ 322 ],
   alphaCSR[ 198 ][ 323 ],
   alphaCSR[ 198 ][ 324 ],
   alphaCSR[ 198 ][ 325 ],
   alphaCSR[ 198 ][ 326 ],
   alphaCSR[ 198 ][ 327 ],
   alphaCSR[ 198 ][ 328 ],
   alphaCSR[ 198 ][ 329 ],
   alphaCSR[ 198 ][ 330 ],
   alphaCSR[ 198 ][ 331 ],
   alphaCSR[ 198 ][ 332 ],
   alphaCSR[ 198 ][ 333 ],
   alphaCSR[ 198 ][ 334 ],
   alphaCSR[ 198 ][ 335 ],
   alphaCSR[ 198 ][ 336 ],
   alphaCSR[ 198 ][ 337 ],
   alphaCSR[ 198 ][ 338 ],
   alphaCSR[ 198 ][ 339 ],
   alphaCSR[ 198 ][ 340 ],
   alphaCSR[ 198 ][ 341 ],
   alphaCSR[ 198 ][ 342 ],
   alphaCSR[ 198 ][ 343 ],
   alphaCSR[ 198 ][ 344 ],
   alphaCSR[ 198 ][ 345 ],
   alphaCSR[ 198 ][ 346 ],
   alphaCSR[ 198 ][ 347 ],
   alphaCSR[ 198 ][ 348 ],
   alphaCSR[ 198 ][ 349 ],
   alphaCSR[ 198 ][ 350 ],
   alphaCSR[ 198 ][ 351 ],
   alphaCSR[ 198 ][ 352 ],
   alphaCSR[ 198 ][ 353 ],
   alphaCSR[ 198 ][ 354 ],
   alphaCSR[ 198 ][ 355 ],
   alphaCSR[ 198 ][ 356 ],
   alphaCSR[ 198 ][ 357 ],
   alphaCSR[ 198 ][ 358 ],
   alphaCSR[ 198 ][ 359 ],
   alphaCSR[ 198 ][ 360 ],
   alphaCSR[ 198 ][ 361 ],
   alphaCSR[ 198 ][ 362 ],
   alphaCSR[ 198 ][ 363 ],
   alphaCSR[ 198 ][ 364 ],
   alphaCSR[ 198 ][ 365 ],
   alphaCSR[ 198 ][ 366 ],
   alphaCSR[ 198 ][ 367 ],
   alphaCSR[ 198 ][ 368 ],
   alphaCSR[ 198 ][ 369 ],
   alphaCSR[ 198 ][ 370 ],
   alphaCSR[ 198 ][ 371 ],
   alphaCSR[ 198 ][ 372 ],
   alphaCSR[ 198 ][ 373 ],
   alphaCSR[ 198 ][ 374 ],
   alphaCSR[ 198 ][ 375 ],
   alphaCSR[ 198 ][ 376 ],
   alphaCSR[ 198 ][ 377 ],
   alphaCSR[ 198 ][ 378 ],
   alphaCSR[ 198 ][ 379 ],
   alphaCSR[ 198 ][ 380 ],
   alphaCSR[ 198 ][ 381 ],
   alphaCSR[ 198 ][ 382 ],
   alphaCSR[ 198 ][ 383 ],
   alphaCSR[ 199 ][ 0 ],
   alphaCSR[ 199 ][ 1 ],
   alphaCSR[ 199 ][ 2 ],
   alphaCSR[ 199 ][ 3 ],
   alphaCSR[ 199 ][ 4 ],
   alphaCSR[ 199 ][ 5 ],
   alphaCSR[ 199 ][ 6 ],
   alphaCSR[ 199 ][ 7 ],
   alphaCSR[ 199 ][ 8 ],
   alphaCSR[ 199 ][ 9 ],
   alphaCSR[ 199 ][ 10 ],
   alphaCSR[ 199 ][ 11 ],
   alphaCSR[ 199 ][ 12 ],
   alphaCSR[ 199 ][ 13 ],
   alphaCSR[ 199 ][ 14 ],
   alphaCSR[ 199 ][ 15 ],
   alphaCSR[ 199 ][ 16 ],
   alphaCSR[ 199 ][ 17 ],
   alphaCSR[ 199 ][ 18 ],
   alphaCSR[ 199 ][ 19 ],
   alphaCSR[ 199 ][ 20 ],
   alphaCSR[ 199 ][ 21 ],
   alphaCSR[ 199 ][ 22 ],
   alphaCSR[ 199 ][ 23 ],
   alphaCSR[ 199 ][ 24 ],
   alphaCSR[ 199 ][ 25 ],
   alphaCSR[ 199 ][ 26 ],
   alphaCSR[ 199 ][ 27 ],
   alphaCSR[ 199 ][ 28 ],
   alphaCSR[ 199 ][ 29 ],
   alphaCSR[ 199 ][ 30 ],
   alphaCSR[ 199 ][ 31 ],
   alphaCSR[ 199 ][ 32 ],
   alphaCSR[ 199 ][ 33 ],
   alphaCSR[ 199 ][ 34 ],
   alphaCSR[ 199 ][ 35 ],
   alphaCSR[ 199 ][ 36 ],
   alphaCSR[ 199 ][ 37 ],
   alphaCSR[ 199 ][ 38 ],
   alphaCSR[ 199 ][ 39 ],
   alphaCSR[ 199 ][ 40 ],
   alphaCSR[ 199 ][ 41 ],
   alphaCSR[ 199 ][ 42 ],
   alphaCSR[ 199 ][ 43 ],
   alphaCSR[ 199 ][ 44 ],
   alphaCSR[ 199 ][ 45 ],
   alphaCSR[ 199 ][ 46 ],
   alphaCSR[ 199 ][ 47 ],
   alphaCSR[ 199 ][ 48 ],
   alphaCSR[ 199 ][ 49 ],
   alphaCSR[ 199 ][ 50 ],
   alphaCSR[ 199 ][ 51 ],
   alphaCSR[ 199 ][ 52 ],
   alphaCSR[ 199 ][ 53 ],
   alphaCSR[ 199 ][ 54 ],
   alphaCSR[ 199 ][ 55 ],
   alphaCSR[ 199 ][ 56 ],
   alphaCSR[ 199 ][ 57 ],
   alphaCSR[ 199 ][ 58 ],
   alphaCSR[ 199 ][ 59 ],
   alphaCSR[ 199 ][ 60 ],
   alphaCSR[ 199 ][ 61 ],
   alphaCSR[ 199 ][ 62 ],
   alphaCSR[ 199 ][ 63 ],
   alphaCSR[ 199 ][ 64 ],
   alphaCSR[ 199 ][ 65 ],
   alphaCSR[ 199 ][ 66 ],
   alphaCSR[ 199 ][ 67 ],
   alphaCSR[ 199 ][ 68 ],
   alphaCSR[ 199 ][ 69 ],
   alphaCSR[ 199 ][ 70 ],
   alphaCSR[ 199 ][ 71 ],
   alphaCSR[ 199 ][ 72 ],
   alphaCSR[ 199 ][ 73 ],
   alphaCSR[ 199 ][ 74 ],
   alphaCSR[ 199 ][ 75 ],
   alphaCSR[ 199 ][ 76 ],
   alphaCSR[ 199 ][ 77 ],
   alphaCSR[ 199 ][ 78 ],
   alphaCSR[ 199 ][ 79 ],
   alphaCSR[ 199 ][ 80 ],
   alphaCSR[ 199 ][ 81 ],
   alphaCSR[ 199 ][ 82 ],
   alphaCSR[ 199 ][ 83 ],
   alphaCSR[ 199 ][ 84 ],
   alphaCSR[ 199 ][ 85 ],
   alphaCSR[ 199 ][ 86 ],
   alphaCSR[ 199 ][ 87 ],
   alphaCSR[ 199 ][ 88 ],
   alphaCSR[ 199 ][ 89 ],
   alphaCSR[ 199 ][ 90 ],
   alphaCSR[ 199 ][ 91 ],
   alphaCSR[ 199 ][ 92 ],
   alphaCSR[ 199 ][ 93 ],
   alphaCSR[ 199 ][ 94 ],
   alphaCSR[ 199 ][ 95 ],
   alphaCSR[ 199 ][ 96 ],
   alphaCSR[ 199 ][ 97 ],
   alphaCSR[ 199 ][ 98 ],
   alphaCSR[ 199 ][ 99 ],
   alphaCSR[ 199 ][ 100 ],
   alphaCSR[ 199 ][ 101 ],
   alphaCSR[ 199 ][ 102 ],
   alphaCSR[ 199 ][ 103 ],
   alphaCSR[ 199 ][ 104 ],
   alphaCSR[ 199 ][ 105 ],
   alphaCSR[ 199 ][ 106 ],
   alphaCSR[ 199 ][ 107 ],
   alphaCSR[ 199 ][ 108 ],
   alphaCSR[ 199 ][ 109 ],
   alphaCSR[ 199 ][ 110 ],
   alphaCSR[ 199 ][ 111 ],
   alphaCSR[ 199 ][ 112 ],
   alphaCSR[ 199 ][ 113 ],
   alphaCSR[ 199 ][ 114 ],
   alphaCSR[ 199 ][ 115 ],
   alphaCSR[ 199 ][ 116 ],
   alphaCSR[ 199 ][ 117 ],
   alphaCSR[ 199 ][ 118 ],
   alphaCSR[ 199 ][ 119 ],
   alphaCSR[ 199 ][ 120 ],
   alphaCSR[ 199 ][ 121 ],
   alphaCSR[ 199 ][ 122 ],
   alphaCSR[ 199 ][ 123 ],
   alphaCSR[ 199 ][ 124 ],
   alphaCSR[ 199 ][ 125 ],
   alphaCSR[ 199 ][ 126 ],
   alphaCSR[ 199 ][ 127 ],
   alphaCSR[ 199 ][ 128 ],
   alphaCSR[ 199 ][ 129 ],
   alphaCSR[ 199 ][ 130 ],
   alphaCSR[ 199 ][ 131 ],
   alphaCSR[ 199 ][ 132 ],
   alphaCSR[ 199 ][ 133 ],
   alphaCSR[ 199 ][ 134 ],
   alphaCSR[ 199 ][ 135 ],
   alphaCSR[ 199 ][ 136 ],
   alphaCSR[ 199 ][ 137 ],
   alphaCSR[ 199 ][ 138 ],
   alphaCSR[ 199 ][ 139 ],
   alphaCSR[ 199 ][ 140 ],
   alphaCSR[ 199 ][ 141 ],
   alphaCSR[ 199 ][ 142 ],
   alphaCSR[ 199 ][ 143 ],
   alphaCSR[ 199 ][ 144 ],
   alphaCSR[ 199 ][ 145 ],
   alphaCSR[ 199 ][ 146 ],
   alphaCSR[ 199 ][ 147 ],
   alphaCSR[ 199 ][ 148 ],
   alphaCSR[ 199 ][ 149 ],
   alphaCSR[ 199 ][ 150 ],
   alphaCSR[ 199 ][ 151 ],
   alphaCSR[ 199 ][ 152 ],
   alphaCSR[ 199 ][ 153 ],
   alphaCSR[ 199 ][ 154 ],
   alphaCSR[ 199 ][ 155 ],
   alphaCSR[ 199 ][ 156 ],
   alphaCSR[ 199 ][ 157 ],
   alphaCSR[ 199 ][ 158 ],
   alphaCSR[ 199 ][ 159 ],
   alphaCSR[ 199 ][ 160 ],
   alphaCSR[ 199 ][ 161 ],
   alphaCSR[ 199 ][ 162 ],
   alphaCSR[ 199 ][ 163 ],
   alphaCSR[ 199 ][ 164 ],
   alphaCSR[ 199 ][ 165 ],
   alphaCSR[ 199 ][ 166 ],
   alphaCSR[ 199 ][ 167 ],
   alphaCSR[ 199 ][ 168 ],
   alphaCSR[ 199 ][ 169 ],
   alphaCSR[ 199 ][ 170 ],
   alphaCSR[ 199 ][ 171 ],
   alphaCSR[ 199 ][ 172 ],
   alphaCSR[ 199 ][ 173 ],
   alphaCSR[ 199 ][ 174 ],
   alphaCSR[ 199 ][ 175 ],
   alphaCSR[ 199 ][ 176 ],
   alphaCSR[ 199 ][ 177 ],
   alphaCSR[ 199 ][ 178 ],
   alphaCSR[ 199 ][ 179 ],
   alphaCSR[ 199 ][ 180 ],
   alphaCSR[ 199 ][ 181 ],
   alphaCSR[ 199 ][ 182 ],
   alphaCSR[ 199 ][ 183 ],
   alphaCSR[ 199 ][ 184 ],
   alphaCSR[ 199 ][ 185 ],
   alphaCSR[ 199 ][ 186 ],
   alphaCSR[ 199 ][ 187 ],
   alphaCSR[ 199 ][ 188 ],
   alphaCSR[ 199 ][ 189 ],
   alphaCSR[ 199 ][ 190 ],
   alphaCSR[ 199 ][ 191 ],
   alphaCSR[ 199 ][ 192 ],
   alphaCSR[ 199 ][ 193 ],
   alphaCSR[ 199 ][ 194 ],
   alphaCSR[ 199 ][ 195 ],
   alphaCSR[ 199 ][ 196 ],
   alphaCSR[ 199 ][ 197 ],
   alphaCSR[ 199 ][ 198 ],
   alphaCSR[ 199 ][ 199 ],
   alphaCSR[ 199 ][ 200 ],
   alphaCSR[ 199 ][ 201 ],
   alphaCSR[ 199 ][ 202 ],
   alphaCSR[ 199 ][ 203 ],
   alphaCSR[ 199 ][ 204 ],
   alphaCSR[ 199 ][ 205 ],
   alphaCSR[ 199 ][ 206 ],
   alphaCSR[ 199 ][ 207 ],
   alphaCSR[ 199 ][ 208 ],
   alphaCSR[ 199 ][ 209 ],
   alphaCSR[ 199 ][ 210 ],
   alphaCSR[ 199 ][ 211 ],
   alphaCSR[ 199 ][ 212 ],
   alphaCSR[ 199 ][ 213 ],
   alphaCSR[ 199 ][ 214 ],
   alphaCSR[ 199 ][ 215 ],
   alphaCSR[ 199 ][ 216 ],
   alphaCSR[ 199 ][ 217 ],
   alphaCSR[ 199 ][ 218 ],
   alphaCSR[ 199 ][ 219 ],
   alphaCSR[ 199 ][ 220 ],
   alphaCSR[ 199 ][ 221 ],
   alphaCSR[ 199 ][ 222 ],
   alphaCSR[ 199 ][ 223 ],
   alphaCSR[ 199 ][ 224 ],
   alphaCSR[ 199 ][ 225 ],
   alphaCSR[ 199 ][ 226 ],
   alphaCSR[ 199 ][ 227 ],
   alphaCSR[ 199 ][ 228 ],
   alphaCSR[ 199 ][ 229 ],
   alphaCSR[ 199 ][ 230 ],
   alphaCSR[ 199 ][ 231 ],
   alphaCSR[ 199 ][ 232 ],
   alphaCSR[ 199 ][ 233 ],
   alphaCSR[ 199 ][ 234 ],
   alphaCSR[ 199 ][ 235 ],
   alphaCSR[ 199 ][ 236 ],
   alphaCSR[ 199 ][ 237 ],
   alphaCSR[ 199 ][ 238 ],
   alphaCSR[ 199 ][ 239 ],
   alphaCSR[ 199 ][ 240 ],
   alphaCSR[ 199 ][ 241 ],
   alphaCSR[ 199 ][ 242 ],
   alphaCSR[ 199 ][ 243 ],
   alphaCSR[ 199 ][ 244 ],
   alphaCSR[ 199 ][ 245 ],
   alphaCSR[ 199 ][ 246 ],
   alphaCSR[ 199 ][ 247 ],
   alphaCSR[ 199 ][ 248 ],
   alphaCSR[ 199 ][ 249 ],
   alphaCSR[ 199 ][ 250 ],
   alphaCSR[ 199 ][ 251 ],
   alphaCSR[ 199 ][ 252 ],
   alphaCSR[ 199 ][ 253 ],
   alphaCSR[ 199 ][ 254 ],
   alphaCSR[ 199 ][ 255 ],
   alphaCSR[ 199 ][ 256 ],
   alphaCSR[ 199 ][ 257 ],
   alphaCSR[ 199 ][ 258 ],
   alphaCSR[ 199 ][ 259 ],
   alphaCSR[ 199 ][ 260 ],
   alphaCSR[ 199 ][ 261 ],
   alphaCSR[ 199 ][ 262 ],
   alphaCSR[ 199 ][ 263 ],
   alphaCSR[ 199 ][ 264 ],
   alphaCSR[ 199 ][ 265 ],
   alphaCSR[ 199 ][ 266 ],
   alphaCSR[ 199 ][ 267 ],
   alphaCSR[ 199 ][ 268 ],
   alphaCSR[ 199 ][ 269 ],
   alphaCSR[ 199 ][ 270 ],
   alphaCSR[ 199 ][ 271 ],
   alphaCSR[ 199 ][ 272 ],
   alphaCSR[ 199 ][ 273 ],
   alphaCSR[ 199 ][ 274 ],
   alphaCSR[ 199 ][ 275 ],
   alphaCSR[ 199 ][ 276 ],
   alphaCSR[ 199 ][ 277 ],
   alphaCSR[ 199 ][ 278 ],
   alphaCSR[ 199 ][ 279 ],
   alphaCSR[ 199 ][ 280 ],
   alphaCSR[ 199 ][ 281 ],
   alphaCSR[ 199 ][ 282 ],
   alphaCSR[ 199 ][ 283 ],
   alphaCSR[ 199 ][ 284 ],
   alphaCSR[ 199 ][ 285 ],
   alphaCSR[ 199 ][ 286 ],
   alphaCSR[ 199 ][ 287 ],
   alphaCSR[ 199 ][ 288 ],
   alphaCSR[ 199 ][ 289 ],
   alphaCSR[ 199 ][ 290 ],
   alphaCSR[ 199 ][ 291 ],
   alphaCSR[ 199 ][ 292 ],
   alphaCSR[ 199 ][ 293 ],
   alphaCSR[ 199 ][ 294 ],
   alphaCSR[ 199 ][ 295 ],
   alphaCSR[ 199 ][ 296 ],
   alphaCSR[ 199 ][ 297 ],
   alphaCSR[ 199 ][ 298 ],
   alphaCSR[ 199 ][ 299 ],
   alphaCSR[ 199 ][ 300 ],
   alphaCSR[ 199 ][ 301 ],
   alphaCSR[ 199 ][ 302 ],
   alphaCSR[ 199 ][ 303 ],
   alphaCSR[ 199 ][ 304 ],
   alphaCSR[ 199 ][ 305 ],
   alphaCSR[ 199 ][ 306 ],
   alphaCSR[ 199 ][ 307 ],
   alphaCSR[ 199 ][ 308 ],
   alphaCSR[ 199 ][ 309 ],
   alphaCSR[ 199 ][ 310 ],
   alphaCSR[ 199 ][ 311 ],
   alphaCSR[ 199 ][ 312 ],
   alphaCSR[ 199 ][ 313 ],
   alphaCSR[ 199 ][ 314 ],
   alphaCSR[ 199 ][ 315 ],
   alphaCSR[ 199 ][ 316 ],
   alphaCSR[ 199 ][ 317 ],
   alphaCSR[ 199 ][ 318 ],
   alphaCSR[ 199 ][ 319 ],
   alphaCSR[ 199 ][ 320 ],
   alphaCSR[ 199 ][ 321 ],
   alphaCSR[ 199 ][ 322 ],
   alphaCSR[ 199 ][ 323 ],
   alphaCSR[ 199 ][ 324 ],
   alphaCSR[ 199 ][ 325 ],
   alphaCSR[ 199 ][ 326 ],
   alphaCSR[ 199 ][ 327 ],
   alphaCSR[ 199 ][ 328 ],
   alphaCSR[ 199 ][ 329 ],
   alphaCSR[ 199 ][ 330 ],
   alphaCSR[ 199 ][ 331 ],
   alphaCSR[ 199 ][ 332 ],
   alphaCSR[ 199 ][ 333 ],
   alphaCSR[ 199 ][ 334 ],
   alphaCSR[ 199 ][ 335 ],
   alphaCSR[ 199 ][ 336 ],
   alphaCSR[ 199 ][ 337 ],
   alphaCSR[ 199 ][ 338 ],
   alphaCSR[ 199 ][ 339 ],
   alphaCSR[ 199 ][ 340 ],
   alphaCSR[ 199 ][ 341 ],
   alphaCSR[ 199 ][ 342 ],
   alphaCSR[ 199 ][ 343 ],
   alphaCSR[ 199 ][ 344 ],
   alphaCSR[ 199 ][ 345 ],
   alphaCSR[ 199 ][ 346 ],
   alphaCSR[ 199 ][ 347 ],
   alphaCSR[ 199 ][ 348 ],
   alphaCSR[ 199 ][ 349 ],
   alphaCSR[ 199 ][ 350 ],
   alphaCSR[ 199 ][ 351 ],
   alphaCSR[ 199 ][ 352 ],
   alphaCSR[ 199 ][ 353 ],
   alphaCSR[ 199 ][ 354 ],
   alphaCSR[ 199 ][ 355 ],
   alphaCSR[ 199 ][ 356 ],
   alphaCSR[ 199 ][ 357 ],
   alphaCSR[ 199 ][ 358 ],
   alphaCSR[ 199 ][ 359 ],
   alphaCSR[ 199 ][ 360 ],
   alphaCSR[ 199 ][ 361 ],
   alphaCSR[ 199 ][ 362 ],
   alphaCSR[ 199 ][ 363 ],
   alphaCSR[ 199 ][ 364 ],
   alphaCSR[ 199 ][ 365 ],
   alphaCSR[ 199 ][ 366 ],
   alphaCSR[ 199 ][ 367 ],
   alphaCSR[ 199 ][ 368 ],
   alphaCSR[ 199 ][ 369 ],
   alphaCSR[ 199 ][ 370 ],
   alphaCSR[ 199 ][ 371 ],
   alphaCSR[ 199 ][ 372 ],
   alphaCSR[ 199 ][ 373 ],
   alphaCSR[ 199 ][ 374 ],
   alphaCSR[ 199 ][ 375 ],
   alphaCSR[ 199 ][ 376 ],
   alphaCSR[ 199 ][ 377 ],
   alphaCSR[ 199 ][ 378 ],
   alphaCSR[ 199 ][ 379 ],
   alphaCSR[ 199 ][ 380 ],
   alphaCSR[ 199 ][ 381 ],
   alphaCSR[ 199 ][ 382 ],
   alphaCSR[ 199 ][ 383 ],
   alphaCSR[ 200 ][ 0 ],
   alphaCSR[ 200 ][ 1 ],
   alphaCSR[ 200 ][ 2 ],
   alphaCSR[ 200 ][ 3 ],
   alphaCSR[ 200 ][ 4 ],
   alphaCSR[ 200 ][ 5 ],
   alphaCSR[ 200 ][ 6 ],
   alphaCSR[ 200 ][ 7 ],
   alphaCSR[ 200 ][ 8 ],
   alphaCSR[ 200 ][ 9 ],
   alphaCSR[ 200 ][ 10 ],
   alphaCSR[ 200 ][ 11 ],
   alphaCSR[ 200 ][ 12 ],
   alphaCSR[ 200 ][ 13 ],
   alphaCSR[ 200 ][ 14 ],
   alphaCSR[ 200 ][ 15 ],
   alphaCSR[ 200 ][ 16 ],
   alphaCSR[ 200 ][ 17 ],
   alphaCSR[ 200 ][ 18 ],
   alphaCSR[ 200 ][ 19 ],
   alphaCSR[ 200 ][ 20 ],
   alphaCSR[ 200 ][ 21 ],
   alphaCSR[ 200 ][ 22 ],
   alphaCSR[ 200 ][ 23 ],
   alphaCSR[ 200 ][ 24 ],
   alphaCSR[ 200 ][ 25 ],
   alphaCSR[ 200 ][ 26 ],
   alphaCSR[ 200 ][ 27 ],
   alphaCSR[ 200 ][ 28 ],
   alphaCSR[ 200 ][ 29 ],
   alphaCSR[ 200 ][ 30 ],
   alphaCSR[ 200 ][ 31 ],
   alphaCSR[ 200 ][ 32 ],
   alphaCSR[ 200 ][ 33 ],
   alphaCSR[ 200 ][ 34 ],
   alphaCSR[ 200 ][ 35 ],
   alphaCSR[ 200 ][ 36 ],
   alphaCSR[ 200 ][ 37 ],
   alphaCSR[ 200 ][ 38 ],
   alphaCSR[ 200 ][ 39 ],
   alphaCSR[ 200 ][ 40 ],
   alphaCSR[ 200 ][ 41 ],
   alphaCSR[ 200 ][ 42 ],
   alphaCSR[ 200 ][ 43 ],
   alphaCSR[ 200 ][ 44 ],
   alphaCSR[ 200 ][ 45 ],
   alphaCSR[ 200 ][ 46 ],
   alphaCSR[ 200 ][ 47 ],
   alphaCSR[ 200 ][ 48 ],
   alphaCSR[ 200 ][ 49 ],
   alphaCSR[ 200 ][ 50 ],
   alphaCSR[ 200 ][ 51 ],
   alphaCSR[ 200 ][ 52 ],
   alphaCSR[ 200 ][ 53 ],
   alphaCSR[ 200 ][ 54 ],
   alphaCSR[ 200 ][ 55 ],
   alphaCSR[ 200 ][ 56 ],
   alphaCSR[ 200 ][ 57 ],
   alphaCSR[ 200 ][ 58 ],
   alphaCSR[ 200 ][ 59 ],
   alphaCSR[ 200 ][ 60 ],
   alphaCSR[ 200 ][ 61 ],
   alphaCSR[ 200 ][ 62 ],
   alphaCSR[ 200 ][ 63 ],
   alphaCSR[ 200 ][ 64 ],
   alphaCSR[ 200 ][ 65 ],
   alphaCSR[ 200 ][ 66 ],
   alphaCSR[ 200 ][ 67 ],
   alphaCSR[ 200 ][ 68 ],
   alphaCSR[ 200 ][ 69 ],
   alphaCSR[ 200 ][ 70 ],
   alphaCSR[ 200 ][ 71 ],
   alphaCSR[ 200 ][ 72 ],
   alphaCSR[ 200 ][ 73 ],
   alphaCSR[ 200 ][ 74 ],
   alphaCSR[ 200 ][ 75 ],
   alphaCSR[ 200 ][ 76 ],
   alphaCSR[ 200 ][ 77 ],
   alphaCSR[ 200 ][ 78 ],
   alphaCSR[ 200 ][ 79 ],
   alphaCSR[ 200 ][ 80 ],
   alphaCSR[ 200 ][ 81 ],
   alphaCSR[ 200 ][ 82 ],
   alphaCSR[ 200 ][ 83 ],
   alphaCSR[ 200 ][ 84 ],
   alphaCSR[ 200 ][ 85 ],
   alphaCSR[ 200 ][ 86 ],
   alphaCSR[ 200 ][ 87 ],
   alphaCSR[ 200 ][ 88 ],
   alphaCSR[ 200 ][ 89 ],
   alphaCSR[ 200 ][ 90 ],
   alphaCSR[ 200 ][ 91 ],
   alphaCSR[ 200 ][ 92 ],
   alphaCSR[ 200 ][ 93 ],
   alphaCSR[ 200 ][ 94 ],
   alphaCSR[ 200 ][ 95 ],
   alphaCSR[ 200 ][ 96 ],
   alphaCSR[ 200 ][ 97 ],
   alphaCSR[ 200 ][ 98 ],
   alphaCSR[ 200 ][ 99 ],
   alphaCSR[ 200 ][ 100 ],
   alphaCSR[ 200 ][ 101 ],
   alphaCSR[ 200 ][ 102 ],
   alphaCSR[ 200 ][ 103 ],
   alphaCSR[ 200 ][ 104 ],
   alphaCSR[ 200 ][ 105 ],
   alphaCSR[ 200 ][ 106 ],
   alphaCSR[ 200 ][ 107 ],
   alphaCSR[ 200 ][ 108 ],
   alphaCSR[ 200 ][ 109 ],
   alphaCSR[ 200 ][ 110 ],
   alphaCSR[ 200 ][ 111 ],
   alphaCSR[ 200 ][ 112 ],
   alphaCSR[ 200 ][ 113 ],
   alphaCSR[ 200 ][ 114 ],
   alphaCSR[ 200 ][ 115 ],
   alphaCSR[ 200 ][ 116 ],
   alphaCSR[ 200 ][ 117 ],
   alphaCSR[ 200 ][ 118 ],
   alphaCSR[ 200 ][ 119 ],
   alphaCSR[ 200 ][ 120 ],
   alphaCSR[ 200 ][ 121 ],
   alphaCSR[ 200 ][ 122 ],
   alphaCSR[ 200 ][ 123 ],
   alphaCSR[ 200 ][ 124 ],
   alphaCSR[ 200 ][ 125 ],
   alphaCSR[ 200 ][ 126 ],
   alphaCSR[ 200 ][ 127 ],
   alphaCSR[ 200 ][ 128 ],
   alphaCSR[ 200 ][ 129 ],
   alphaCSR[ 200 ][ 130 ],
   alphaCSR[ 200 ][ 131 ],
   alphaCSR[ 200 ][ 132 ],
   alphaCSR[ 200 ][ 133 ],
   alphaCSR[ 200 ][ 134 ],
   alphaCSR[ 200 ][ 135 ],
   alphaCSR[ 200 ][ 136 ],
   alphaCSR[ 200 ][ 137 ],
   alphaCSR[ 200 ][ 138 ],
   alphaCSR[ 200 ][ 139 ],
   alphaCSR[ 200 ][ 140 ],
   alphaCSR[ 200 ][ 141 ],
   alphaCSR[ 200 ][ 142 ],
   alphaCSR[ 200 ][ 143 ],
   alphaCSR[ 200 ][ 144 ],
   alphaCSR[ 200 ][ 145 ],
   alphaCSR[ 200 ][ 146 ],
   alphaCSR[ 200 ][ 147 ],
   alphaCSR[ 200 ][ 148 ],
   alphaCSR[ 200 ][ 149 ],
   alphaCSR[ 200 ][ 150 ],
   alphaCSR[ 200 ][ 151 ],
   alphaCSR[ 200 ][ 152 ],
   alphaCSR[ 200 ][ 153 ],
   alphaCSR[ 200 ][ 154 ],
   alphaCSR[ 200 ][ 155 ],
   alphaCSR[ 200 ][ 156 ],
   alphaCSR[ 200 ][ 157 ],
   alphaCSR[ 200 ][ 158 ],
   alphaCSR[ 200 ][ 159 ],
   alphaCSR[ 200 ][ 160 ],
   alphaCSR[ 200 ][ 161 ],
   alphaCSR[ 200 ][ 162 ],
   alphaCSR[ 200 ][ 163 ],
   alphaCSR[ 200 ][ 164 ],
   alphaCSR[ 200 ][ 165 ],
   alphaCSR[ 200 ][ 166 ],
   alphaCSR[ 200 ][ 167 ],
   alphaCSR[ 200 ][ 168 ],
   alphaCSR[ 200 ][ 169 ],
   alphaCSR[ 200 ][ 170 ],
   alphaCSR[ 200 ][ 171 ],
   alphaCSR[ 200 ][ 172 ],
   alphaCSR[ 200 ][ 173 ],
   alphaCSR[ 200 ][ 174 ],
   alphaCSR[ 200 ][ 175 ],
   alphaCSR[ 200 ][ 176 ],
   alphaCSR[ 200 ][ 177 ],
   alphaCSR[ 200 ][ 178 ],
   alphaCSR[ 200 ][ 179 ],
   alphaCSR[ 200 ][ 180 ],
   alphaCSR[ 200 ][ 181 ],
   alphaCSR[ 200 ][ 182 ],
   alphaCSR[ 200 ][ 183 ],
   alphaCSR[ 200 ][ 184 ],
   alphaCSR[ 200 ][ 185 ],
   alphaCSR[ 200 ][ 186 ],
   alphaCSR[ 200 ][ 187 ],
   alphaCSR[ 200 ][ 188 ],
   alphaCSR[ 200 ][ 189 ],
   alphaCSR[ 200 ][ 190 ],
   alphaCSR[ 200 ][ 191 ],
   alphaCSR[ 200 ][ 192 ],
   alphaCSR[ 200 ][ 193 ],
   alphaCSR[ 200 ][ 194 ],
   alphaCSR[ 200 ][ 195 ],
   alphaCSR[ 200 ][ 196 ],
   alphaCSR[ 200 ][ 197 ],
   alphaCSR[ 200 ][ 198 ],
   alphaCSR[ 200 ][ 199 ],
   alphaCSR[ 200 ][ 200 ],
   alphaCSR[ 200 ][ 201 ],
   alphaCSR[ 200 ][ 202 ],
   alphaCSR[ 200 ][ 203 ],
   alphaCSR[ 200 ][ 204 ],
   alphaCSR[ 200 ][ 205 ],
   alphaCSR[ 200 ][ 206 ],
   alphaCSR[ 200 ][ 207 ],
   alphaCSR[ 200 ][ 208 ],
   alphaCSR[ 200 ][ 209 ],
   alphaCSR[ 200 ][ 210 ],
   alphaCSR[ 200 ][ 211 ],
   alphaCSR[ 200 ][ 212 ],
   alphaCSR[ 200 ][ 213 ],
   alphaCSR[ 200 ][ 214 ],
   alphaCSR[ 200 ][ 215 ],
   alphaCSR[ 200 ][ 216 ],
   alphaCSR[ 200 ][ 217 ],
   alphaCSR[ 200 ][ 218 ],
   alphaCSR[ 200 ][ 219 ],
   alphaCSR[ 200 ][ 220 ],
   alphaCSR[ 200 ][ 221 ],
   alphaCSR[ 200 ][ 222 ],
   alphaCSR[ 200 ][ 223 ],
   alphaCSR[ 200 ][ 224 ],
   alphaCSR[ 200 ][ 225 ],
   alphaCSR[ 200 ][ 226 ],
   alphaCSR[ 200 ][ 227 ],
   alphaCSR[ 200 ][ 228 ],
   alphaCSR[ 200 ][ 229 ],
   alphaCSR[ 200 ][ 230 ],
   alphaCSR[ 200 ][ 231 ],
   alphaCSR[ 200 ][ 232 ],
   alphaCSR[ 200 ][ 233 ],
   alphaCSR[ 200 ][ 234 ],
   alphaCSR[ 200 ][ 235 ],
   alphaCSR[ 200 ][ 236 ],
   alphaCSR[ 200 ][ 237 ],
   alphaCSR[ 200 ][ 238 ],
   alphaCSR[ 200 ][ 239 ],
   alphaCSR[ 200 ][ 240 ],
   alphaCSR[ 200 ][ 241 ],
   alphaCSR[ 200 ][ 242 ],
   alphaCSR[ 200 ][ 243 ],
   alphaCSR[ 200 ][ 244 ],
   alphaCSR[ 200 ][ 245 ],
   alphaCSR[ 200 ][ 246 ],
   alphaCSR[ 200 ][ 247 ],
   alphaCSR[ 200 ][ 248 ],
   alphaCSR[ 200 ][ 249 ],
   alphaCSR[ 200 ][ 250 ],
   alphaCSR[ 200 ][ 251 ],
   alphaCSR[ 200 ][ 252 ],
   alphaCSR[ 200 ][ 253 ],
   alphaCSR[ 200 ][ 254 ],
   alphaCSR[ 200 ][ 255 ],
   alphaCSR[ 200 ][ 256 ],
   alphaCSR[ 200 ][ 257 ],
   alphaCSR[ 200 ][ 258 ],
   alphaCSR[ 200 ][ 259 ],
   alphaCSR[ 200 ][ 260 ],
   alphaCSR[ 200 ][ 261 ],
   alphaCSR[ 200 ][ 262 ],
   alphaCSR[ 200 ][ 263 ],
   alphaCSR[ 200 ][ 264 ],
   alphaCSR[ 200 ][ 265 ],
   alphaCSR[ 200 ][ 266 ],
   alphaCSR[ 200 ][ 267 ],
   alphaCSR[ 200 ][ 268 ],
   alphaCSR[ 200 ][ 269 ],
   alphaCSR[ 200 ][ 270 ],
   alphaCSR[ 200 ][ 271 ],
   alphaCSR[ 200 ][ 272 ],
   alphaCSR[ 200 ][ 273 ],
   alphaCSR[ 200 ][ 274 ],
   alphaCSR[ 200 ][ 275 ],
   alphaCSR[ 200 ][ 276 ],
   alphaCSR[ 200 ][ 277 ],
   alphaCSR[ 200 ][ 278 ],
   alphaCSR[ 200 ][ 279 ],
   alphaCSR[ 200 ][ 280 ],
   alphaCSR[ 200 ][ 281 ],
   alphaCSR[ 200 ][ 282 ],
   alphaCSR[ 200 ][ 283 ],
   alphaCSR[ 200 ][ 284 ],
   alphaCSR[ 200 ][ 285 ],
   alphaCSR[ 200 ][ 286 ],
   alphaCSR[ 200 ][ 287 ],
   alphaCSR[ 200 ][ 288 ],
   alphaCSR[ 200 ][ 289 ],
   alphaCSR[ 200 ][ 290 ],
   alphaCSR[ 200 ][ 291 ],
   alphaCSR[ 200 ][ 292 ],
   alphaCSR[ 200 ][ 293 ],
   alphaCSR[ 200 ][ 294 ],
   alphaCSR[ 200 ][ 295 ],
   alphaCSR[ 200 ][ 296 ],
   alphaCSR[ 200 ][ 297 ],
   alphaCSR[ 200 ][ 298 ],
   alphaCSR[ 200 ][ 299 ],
   alphaCSR[ 200 ][ 300 ],
   alphaCSR[ 200 ][ 301 ],
   alphaCSR[ 200 ][ 302 ],
   alphaCSR[ 200 ][ 303 ],
   alphaCSR[ 200 ][ 304 ],
   alphaCSR[ 200 ][ 305 ],
   alphaCSR[ 200 ][ 306 ],
   alphaCSR[ 200 ][ 307 ],
   alphaCSR[ 200 ][ 308 ],
   alphaCSR[ 200 ][ 309 ],
   alphaCSR[ 200 ][ 310 ],
   alphaCSR[ 200 ][ 311 ],
   alphaCSR[ 200 ][ 312 ],
   alphaCSR[ 200 ][ 313 ],
   alphaCSR[ 200 ][ 314 ],
   alphaCSR[ 200 ][ 315 ],
   alphaCSR[ 200 ][ 316 ],
   alphaCSR[ 200 ][ 317 ],
   alphaCSR[ 200 ][ 318 ],
   alphaCSR[ 200 ][ 319 ],
   alphaCSR[ 200 ][ 320 ],
   alphaCSR[ 200 ][ 321 ],
   alphaCSR[ 200 ][ 322 ],
   alphaCSR[ 200 ][ 323 ],
   alphaCSR[ 200 ][ 324 ],
   alphaCSR[ 200 ][ 325 ],
   alphaCSR[ 200 ][ 326 ],
   alphaCSR[ 200 ][ 327 ],
   alphaCSR[ 200 ][ 328 ],
   alphaCSR[ 200 ][ 329 ],
   alphaCSR[ 200 ][ 330 ],
   alphaCSR[ 200 ][ 331 ],
   alphaCSR[ 200 ][ 332 ],
   alphaCSR[ 200 ][ 333 ],
   alphaCSR[ 200 ][ 334 ],
   alphaCSR[ 200 ][ 335 ],
   alphaCSR[ 200 ][ 336 ],
   alphaCSR[ 200 ][ 337 ],
   alphaCSR[ 200 ][ 338 ],
   alphaCSR[ 200 ][ 339 ],
   alphaCSR[ 200 ][ 340 ],
   alphaCSR[ 200 ][ 341 ],
   alphaCSR[ 200 ][ 342 ],
   alphaCSR[ 200 ][ 343 ],
   alphaCSR[ 200 ][ 344 ],
   alphaCSR[ 200 ][ 345 ],
   alphaCSR[ 200 ][ 346 ],
   alphaCSR[ 200 ][ 347 ],
   alphaCSR[ 200 ][ 348 ],
   alphaCSR[ 200 ][ 349 ],
   alphaCSR[ 200 ][ 350 ],
   alphaCSR[ 200 ][ 351 ],
   alphaCSR[ 200 ][ 352 ],
   alphaCSR[ 200 ][ 353 ],
   alphaCSR[ 200 ][ 354 ],
   alphaCSR[ 200 ][ 355 ],
   alphaCSR[ 200 ][ 356 ],
   alphaCSR[ 200 ][ 357 ],
   alphaCSR[ 200 ][ 358 ],
   alphaCSR[ 200 ][ 359 ],
   alphaCSR[ 200 ][ 360 ],
   alphaCSR[ 200 ][ 361 ],
   alphaCSR[ 200 ][ 362 ],
   alphaCSR[ 200 ][ 363 ],
   alphaCSR[ 200 ][ 364 ],
   alphaCSR[ 200 ][ 365 ],
   alphaCSR[ 200 ][ 366 ],
   alphaCSR[ 200 ][ 367 ],
   alphaCSR[ 200 ][ 368 ],
   alphaCSR[ 200 ][ 369 ],
   alphaCSR[ 200 ][ 370 ],
   alphaCSR[ 200 ][ 371 ],
   alphaCSR[ 200 ][ 372 ],
   alphaCSR[ 200 ][ 373 ],
   alphaCSR[ 200 ][ 374 ],
   alphaCSR[ 200 ][ 375 ],
   alphaCSR[ 200 ][ 376 ],
   alphaCSR[ 200 ][ 377 ],
   alphaCSR[ 200 ][ 378 ],
   alphaCSR[ 200 ][ 379 ],
   alphaCSR[ 200 ][ 380 ],
   alphaCSR[ 200 ][ 381 ],
   alphaCSR[ 200 ][ 382 ],
   alphaCSR[ 200 ][ 383 ],
   alphaCSR[ 201 ][ 0 ],
   alphaCSR[ 201 ][ 1 ],
   alphaCSR[ 201 ][ 2 ],
   alphaCSR[ 201 ][ 3 ],
   alphaCSR[ 201 ][ 4 ],
   alphaCSR[ 201 ][ 5 ],
   alphaCSR[ 201 ][ 6 ],
   alphaCSR[ 201 ][ 7 ],
   alphaCSR[ 201 ][ 8 ],
   alphaCSR[ 201 ][ 9 ],
   alphaCSR[ 201 ][ 10 ],
   alphaCSR[ 201 ][ 11 ],
   alphaCSR[ 201 ][ 12 ],
   alphaCSR[ 201 ][ 13 ],
   alphaCSR[ 201 ][ 14 ],
   alphaCSR[ 201 ][ 15 ],
   alphaCSR[ 201 ][ 16 ],
   alphaCSR[ 201 ][ 17 ],
   alphaCSR[ 201 ][ 18 ],
   alphaCSR[ 201 ][ 19 ],
   alphaCSR[ 201 ][ 20 ],
   alphaCSR[ 201 ][ 21 ],
   alphaCSR[ 201 ][ 22 ],
   alphaCSR[ 201 ][ 23 ],
   alphaCSR[ 201 ][ 24 ],
   alphaCSR[ 201 ][ 25 ],
   alphaCSR[ 201 ][ 26 ],
   alphaCSR[ 201 ][ 27 ],
   alphaCSR[ 201 ][ 28 ],
   alphaCSR[ 201 ][ 29 ],
   alphaCSR[ 201 ][ 30 ],
   alphaCSR[ 201 ][ 31 ],
   alphaCSR[ 201 ][ 32 ],
   alphaCSR[ 201 ][ 33 ],
   alphaCSR[ 201 ][ 34 ],
   alphaCSR[ 201 ][ 35 ],
   alphaCSR[ 201 ][ 36 ],
   alphaCSR[ 201 ][ 37 ],
   alphaCSR[ 201 ][ 38 ],
   alphaCSR[ 201 ][ 39 ],
   alphaCSR[ 201 ][ 40 ],
   alphaCSR[ 201 ][ 41 ],
   alphaCSR[ 201 ][ 42 ],
   alphaCSR[ 201 ][ 43 ],
   alphaCSR[ 201 ][ 44 ],
   alphaCSR[ 201 ][ 45 ],
   alphaCSR[ 201 ][ 46 ],
   alphaCSR[ 201 ][ 47 ],
   alphaCSR[ 201 ][ 48 ],
   alphaCSR[ 201 ][ 49 ],
   alphaCSR[ 201 ][ 50 ],
   alphaCSR[ 201 ][ 51 ],
   alphaCSR[ 201 ][ 52 ],
   alphaCSR[ 201 ][ 53 ],
   alphaCSR[ 201 ][ 54 ],
   alphaCSR[ 201 ][ 55 ],
   alphaCSR[ 201 ][ 56 ],
   alphaCSR[ 201 ][ 57 ],
   alphaCSR[ 201 ][ 58 ],
   alphaCSR[ 201 ][ 59 ],
   alphaCSR[ 201 ][ 60 ],
   alphaCSR[ 201 ][ 61 ],
   alphaCSR[ 201 ][ 62 ],
   alphaCSR[ 201 ][ 63 ],
   alphaCSR[ 201 ][ 64 ],
   alphaCSR[ 201 ][ 65 ],
   alphaCSR[ 201 ][ 66 ],
   alphaCSR[ 201 ][ 67 ],
   alphaCSR[ 201 ][ 68 ],
   alphaCSR[ 201 ][ 69 ],
   alphaCSR[ 201 ][ 70 ],
   alphaCSR[ 201 ][ 71 ],
   alphaCSR[ 201 ][ 72 ],
   alphaCSR[ 201 ][ 73 ],
   alphaCSR[ 201 ][ 74 ],
   alphaCSR[ 201 ][ 75 ],
   alphaCSR[ 201 ][ 76 ],
   alphaCSR[ 201 ][ 77 ],
   alphaCSR[ 201 ][ 78 ],
   alphaCSR[ 201 ][ 79 ],
   alphaCSR[ 201 ][ 80 ],
   alphaCSR[ 201 ][ 81 ],
   alphaCSR[ 201 ][ 82 ],
   alphaCSR[ 201 ][ 83 ],
   alphaCSR[ 201 ][ 84 ],
   alphaCSR[ 201 ][ 85 ],
   alphaCSR[ 201 ][ 86 ],
   alphaCSR[ 201 ][ 87 ],
   alphaCSR[ 201 ][ 88 ],
   alphaCSR[ 201 ][ 89 ],
   alphaCSR[ 201 ][ 90 ],
   alphaCSR[ 201 ][ 91 ],
   alphaCSR[ 201 ][ 92 ],
   alphaCSR[ 201 ][ 93 ],
   alphaCSR[ 201 ][ 94 ],
   alphaCSR[ 201 ][ 95 ],
   alphaCSR[ 201 ][ 96 ],
   alphaCSR[ 201 ][ 97 ],
   alphaCSR[ 201 ][ 98 ],
   alphaCSR[ 201 ][ 99 ],
   alphaCSR[ 201 ][ 100 ],
   alphaCSR[ 201 ][ 101 ],
   alphaCSR[ 201 ][ 102 ],
   alphaCSR[ 201 ][ 103 ],
   alphaCSR[ 201 ][ 104 ],
   alphaCSR[ 201 ][ 105 ],
   alphaCSR[ 201 ][ 106 ],
   alphaCSR[ 201 ][ 107 ],
   alphaCSR[ 201 ][ 108 ],
   alphaCSR[ 201 ][ 109 ],
   alphaCSR[ 201 ][ 110 ],
   alphaCSR[ 201 ][ 111 ],
   alphaCSR[ 201 ][ 112 ],
   alphaCSR[ 201 ][ 113 ],
   alphaCSR[ 201 ][ 114 ],
   alphaCSR[ 201 ][ 115 ],
   alphaCSR[ 201 ][ 116 ],
   alphaCSR[ 201 ][ 117 ],
   alphaCSR[ 201 ][ 118 ],
   alphaCSR[ 201 ][ 119 ],
   alphaCSR[ 201 ][ 120 ],
   alphaCSR[ 201 ][ 121 ],
   alphaCSR[ 201 ][ 122 ],
   alphaCSR[ 201 ][ 123 ],
   alphaCSR[ 201 ][ 124 ],
   alphaCSR[ 201 ][ 125 ],
   alphaCSR[ 201 ][ 126 ],
   alphaCSR[ 201 ][ 127 ],
   alphaCSR[ 201 ][ 128 ],
   alphaCSR[ 201 ][ 129 ],
   alphaCSR[ 201 ][ 130 ],
   alphaCSR[ 201 ][ 131 ],
   alphaCSR[ 201 ][ 132 ],
   alphaCSR[ 201 ][ 133 ],
   alphaCSR[ 201 ][ 134 ],
   alphaCSR[ 201 ][ 135 ],
   alphaCSR[ 201 ][ 136 ],
   alphaCSR[ 201 ][ 137 ],
   alphaCSR[ 201 ][ 138 ],
   alphaCSR[ 201 ][ 139 ],
   alphaCSR[ 201 ][ 140 ],
   alphaCSR[ 201 ][ 141 ],
   alphaCSR[ 201 ][ 142 ],
   alphaCSR[ 201 ][ 143 ],
   alphaCSR[ 201 ][ 144 ],
   alphaCSR[ 201 ][ 145 ],
   alphaCSR[ 201 ][ 146 ],
   alphaCSR[ 201 ][ 147 ],
   alphaCSR[ 201 ][ 148 ],
   alphaCSR[ 201 ][ 149 ],
   alphaCSR[ 201 ][ 150 ],
   alphaCSR[ 201 ][ 151 ],
   alphaCSR[ 201 ][ 152 ],
   alphaCSR[ 201 ][ 153 ],
   alphaCSR[ 201 ][ 154 ],
   alphaCSR[ 201 ][ 155 ],
   alphaCSR[ 201 ][ 156 ],
   alphaCSR[ 201 ][ 157 ],
   alphaCSR[ 201 ][ 158 ],
   alphaCSR[ 201 ][ 159 ],
   alphaCSR[ 201 ][ 160 ],
   alphaCSR[ 201 ][ 161 ],
   alphaCSR[ 201 ][ 162 ],
   alphaCSR[ 201 ][ 163 ],
   alphaCSR[ 201 ][ 164 ],
   alphaCSR[ 201 ][ 165 ],
   alphaCSR[ 201 ][ 166 ],
   alphaCSR[ 201 ][ 167 ],
   alphaCSR[ 201 ][ 168 ],
   alphaCSR[ 201 ][ 169 ],
   alphaCSR[ 201 ][ 170 ],
   alphaCSR[ 201 ][ 171 ],
   alphaCSR[ 201 ][ 172 ],
   alphaCSR[ 201 ][ 173 ],
   alphaCSR[ 201 ][ 174 ],
   alphaCSR[ 201 ][ 175 ],
   alphaCSR[ 201 ][ 176 ],
   alphaCSR[ 201 ][ 177 ],
   alphaCSR[ 201 ][ 178 ],
   alphaCSR[ 201 ][ 179 ],
   alphaCSR[ 201 ][ 180 ],
   alphaCSR[ 201 ][ 181 ],
   alphaCSR[ 201 ][ 182 ],
   alphaCSR[ 201 ][ 183 ],
   alphaCSR[ 201 ][ 184 ],
   alphaCSR[ 201 ][ 185 ],
   alphaCSR[ 201 ][ 186 ],
   alphaCSR[ 201 ][ 187 ],
   alphaCSR[ 201 ][ 188 ],
   alphaCSR[ 201 ][ 189 ],
   alphaCSR[ 201 ][ 190 ],
   alphaCSR[ 201 ][ 191 ],
   alphaCSR[ 201 ][ 192 ],
   alphaCSR[ 201 ][ 193 ],
   alphaCSR[ 201 ][ 194 ],
   alphaCSR[ 201 ][ 195 ],
   alphaCSR[ 201 ][ 196 ],
   alphaCSR[ 201 ][ 197 ],
   alphaCSR[ 201 ][ 198 ],
   alphaCSR[ 201 ][ 199 ],
   alphaCSR[ 201 ][ 200 ],
   alphaCSR[ 201 ][ 201 ],
   alphaCSR[ 201 ][ 202 ],
   alphaCSR[ 201 ][ 203 ],
   alphaCSR[ 201 ][ 204 ],
   alphaCSR[ 201 ][ 205 ],
   alphaCSR[ 201 ][ 206 ],
   alphaCSR[ 201 ][ 207 ],
   alphaCSR[ 201 ][ 208 ],
   alphaCSR[ 201 ][ 209 ],
   alphaCSR[ 201 ][ 210 ],
   alphaCSR[ 201 ][ 211 ],
   alphaCSR[ 201 ][ 212 ],
   alphaCSR[ 201 ][ 213 ],
   alphaCSR[ 201 ][ 214 ],
   alphaCSR[ 201 ][ 215 ],
   alphaCSR[ 201 ][ 216 ],
   alphaCSR[ 201 ][ 217 ],
   alphaCSR[ 201 ][ 218 ],
   alphaCSR[ 201 ][ 219 ],
   alphaCSR[ 201 ][ 220 ],
   alphaCSR[ 201 ][ 221 ],
   alphaCSR[ 201 ][ 222 ],
   alphaCSR[ 201 ][ 223 ],
   alphaCSR[ 201 ][ 224 ],
   alphaCSR[ 201 ][ 225 ],
   alphaCSR[ 201 ][ 226 ],
   alphaCSR[ 201 ][ 227 ],
   alphaCSR[ 201 ][ 228 ],
   alphaCSR[ 201 ][ 229 ],
   alphaCSR[ 201 ][ 230 ],
   alphaCSR[ 201 ][ 231 ],
   alphaCSR[ 201 ][ 232 ],
   alphaCSR[ 201 ][ 233 ],
   alphaCSR[ 201 ][ 234 ],
   alphaCSR[ 201 ][ 235 ],
   alphaCSR[ 201 ][ 236 ],
   alphaCSR[ 201 ][ 237 ],
   alphaCSR[ 201 ][ 238 ],
   alphaCSR[ 201 ][ 239 ],
   alphaCSR[ 201 ][ 240 ],
   alphaCSR[ 201 ][ 241 ],
   alphaCSR[ 201 ][ 242 ],
   alphaCSR[ 201 ][ 243 ],
   alphaCSR[ 201 ][ 244 ],
   alphaCSR[ 201 ][ 245 ],
   alphaCSR[ 201 ][ 246 ],
   alphaCSR[ 201 ][ 247 ],
   alphaCSR[ 201 ][ 248 ],
   alphaCSR[ 201 ][ 249 ],
   alphaCSR[ 201 ][ 250 ],
   alphaCSR[ 201 ][ 251 ],
   alphaCSR[ 201 ][ 252 ],
   alphaCSR[ 201 ][ 253 ],
   alphaCSR[ 201 ][ 254 ],
   alphaCSR[ 201 ][ 255 ],
   alphaCSR[ 201 ][ 256 ],
   alphaCSR[ 201 ][ 257 ],
   alphaCSR[ 201 ][ 258 ],
   alphaCSR[ 201 ][ 259 ],
   alphaCSR[ 201 ][ 260 ],
   alphaCSR[ 201 ][ 261 ],
   alphaCSR[ 201 ][ 262 ],
   alphaCSR[ 201 ][ 263 ],
   alphaCSR[ 201 ][ 264 ],
   alphaCSR[ 201 ][ 265 ],
   alphaCSR[ 201 ][ 266 ],
   alphaCSR[ 201 ][ 267 ],
   alphaCSR[ 201 ][ 268 ],
   alphaCSR[ 201 ][ 269 ],
   alphaCSR[ 201 ][ 270 ],
   alphaCSR[ 201 ][ 271 ],
   alphaCSR[ 201 ][ 272 ],
   alphaCSR[ 201 ][ 273 ],
   alphaCSR[ 201 ][ 274 ],
   alphaCSR[ 201 ][ 275 ],
   alphaCSR[ 201 ][ 276 ],
   alphaCSR[ 201 ][ 277 ],
   alphaCSR[ 201 ][ 278 ],
   alphaCSR[ 201 ][ 279 ],
   alphaCSR[ 201 ][ 280 ],
   alphaCSR[ 201 ][ 281 ],
   alphaCSR[ 201 ][ 282 ],
   alphaCSR[ 201 ][ 283 ],
   alphaCSR[ 201 ][ 284 ],
   alphaCSR[ 201 ][ 285 ],
   alphaCSR[ 201 ][ 286 ],
   alphaCSR[ 201 ][ 287 ],
   alphaCSR[ 201 ][ 288 ],
   alphaCSR[ 201 ][ 289 ],
   alphaCSR[ 201 ][ 290 ],
   alphaCSR[ 201 ][ 291 ],
   alphaCSR[ 201 ][ 292 ],
   alphaCSR[ 201 ][ 293 ],
   alphaCSR[ 201 ][ 294 ],
   alphaCSR[ 201 ][ 295 ],
   alphaCSR[ 201 ][ 296 ],
   alphaCSR[ 201 ][ 297 ],
   alphaCSR[ 201 ][ 298 ],
   alphaCSR[ 201 ][ 299 ],
   alphaCSR[ 201 ][ 300 ],
   alphaCSR[ 201 ][ 301 ],
   alphaCSR[ 201 ][ 302 ],
   alphaCSR[ 201 ][ 303 ],
   alphaCSR[ 201 ][ 304 ],
   alphaCSR[ 201 ][ 305 ],
   alphaCSR[ 201 ][ 306 ],
   alphaCSR[ 201 ][ 307 ],
   alphaCSR[ 201 ][ 308 ],
   alphaCSR[ 201 ][ 309 ],
   alphaCSR[ 201 ][ 310 ],
   alphaCSR[ 201 ][ 311 ],
   alphaCSR[ 201 ][ 312 ],
   alphaCSR[ 201 ][ 313 ],
   alphaCSR[ 201 ][ 314 ],
   alphaCSR[ 201 ][ 315 ],
   alphaCSR[ 201 ][ 316 ],
   alphaCSR[ 201 ][ 317 ],
   alphaCSR[ 201 ][ 318 ],
   alphaCSR[ 201 ][ 319 ],
   alphaCSR[ 201 ][ 320 ],
   alphaCSR[ 201 ][ 321 ],
   alphaCSR[ 201 ][ 322 ],
   alphaCSR[ 201 ][ 323 ],
   alphaCSR[ 201 ][ 324 ],
   alphaCSR[ 201 ][ 325 ],
   alphaCSR[ 201 ][ 326 ],
   alphaCSR[ 201 ][ 327 ],
   alphaCSR[ 201 ][ 328 ],
   alphaCSR[ 201 ][ 329 ],
   alphaCSR[ 201 ][ 330 ],
   alphaCSR[ 201 ][ 331 ],
   alphaCSR[ 201 ][ 332 ],
   alphaCSR[ 201 ][ 333 ],
   alphaCSR[ 201 ][ 334 ],
   alphaCSR[ 201 ][ 335 ],
   alphaCSR[ 201 ][ 336 ],
   alphaCSR[ 201 ][ 337 ],
   alphaCSR[ 201 ][ 338 ],
   alphaCSR[ 201 ][ 339 ],
   alphaCSR[ 201 ][ 340 ],
   alphaCSR[ 201 ][ 341 ],
   alphaCSR[ 201 ][ 342 ],
   alphaCSR[ 201 ][ 343 ],
   alphaCSR[ 201 ][ 344 ],
   alphaCSR[ 201 ][ 345 ],
   alphaCSR[ 201 ][ 346 ],
   alphaCSR[ 201 ][ 347 ],
   alphaCSR[ 201 ][ 348 ],
   alphaCSR[ 201 ][ 349 ],
   alphaCSR[ 201 ][ 350 ],
   alphaCSR[ 201 ][ 351 ],
   alphaCSR[ 201 ][ 352 ],
   alphaCSR[ 201 ][ 353 ],
   alphaCSR[ 201 ][ 354 ],
   alphaCSR[ 201 ][ 355 ],
   alphaCSR[ 201 ][ 356 ],
   alphaCSR[ 201 ][ 357 ],
   alphaCSR[ 201 ][ 358 ],
   alphaCSR[ 201 ][ 359 ],
   alphaCSR[ 201 ][ 360 ],
   alphaCSR[ 201 ][ 361 ],
   alphaCSR[ 201 ][ 362 ],
   alphaCSR[ 201 ][ 363 ],
   alphaCSR[ 201 ][ 364 ],
   alphaCSR[ 201 ][ 365 ],
   alphaCSR[ 201 ][ 366 ],
   alphaCSR[ 201 ][ 367 ],
   alphaCSR[ 201 ][ 368 ],
   alphaCSR[ 201 ][ 369 ],
   alphaCSR[ 201 ][ 370 ],
   alphaCSR[ 201 ][ 371 ],
   alphaCSR[ 201 ][ 372 ],
   alphaCSR[ 201 ][ 373 ],
   alphaCSR[ 201 ][ 374 ],
   alphaCSR[ 201 ][ 375 ],
   alphaCSR[ 201 ][ 376 ],
   alphaCSR[ 201 ][ 377 ],
   alphaCSR[ 201 ][ 378 ],
   alphaCSR[ 201 ][ 379 ],
   alphaCSR[ 201 ][ 380 ],
   alphaCSR[ 201 ][ 381 ],
   alphaCSR[ 201 ][ 382 ],
   alphaCSR[ 201 ][ 383 ],
   alphaCSR[ 202 ][ 0 ],
   alphaCSR[ 202 ][ 1 ],
   alphaCSR[ 202 ][ 2 ],
   alphaCSR[ 202 ][ 3 ],
   alphaCSR[ 202 ][ 4 ],
   alphaCSR[ 202 ][ 5 ],
   alphaCSR[ 202 ][ 6 ],
   alphaCSR[ 202 ][ 7 ],
   alphaCSR[ 202 ][ 8 ],
   alphaCSR[ 202 ][ 9 ],
   alphaCSR[ 202 ][ 10 ],
   alphaCSR[ 202 ][ 11 ],
   alphaCSR[ 202 ][ 12 ],
   alphaCSR[ 202 ][ 13 ],
   alphaCSR[ 202 ][ 14 ],
   alphaCSR[ 202 ][ 15 ],
   alphaCSR[ 202 ][ 16 ],
   alphaCSR[ 202 ][ 17 ],
   alphaCSR[ 202 ][ 18 ],
   alphaCSR[ 202 ][ 19 ],
   alphaCSR[ 202 ][ 20 ],
   alphaCSR[ 202 ][ 21 ],
   alphaCSR[ 202 ][ 22 ],
   alphaCSR[ 202 ][ 23 ],
   alphaCSR[ 202 ][ 24 ],
   alphaCSR[ 202 ][ 25 ],
   alphaCSR[ 202 ][ 26 ],
   alphaCSR[ 202 ][ 27 ],
   alphaCSR[ 202 ][ 28 ],
   alphaCSR[ 202 ][ 29 ],
   alphaCSR[ 202 ][ 30 ],
   alphaCSR[ 202 ][ 31 ],
   alphaCSR[ 202 ][ 32 ],
   alphaCSR[ 202 ][ 33 ],
   alphaCSR[ 202 ][ 34 ],
   alphaCSR[ 202 ][ 35 ],
   alphaCSR[ 202 ][ 36 ],
   alphaCSR[ 202 ][ 37 ],
   alphaCSR[ 202 ][ 38 ],
   alphaCSR[ 202 ][ 39 ],
   alphaCSR[ 202 ][ 40 ],
   alphaCSR[ 202 ][ 41 ],
   alphaCSR[ 202 ][ 42 ],
   alphaCSR[ 202 ][ 43 ],
   alphaCSR[ 202 ][ 44 ],
   alphaCSR[ 202 ][ 45 ],
   alphaCSR[ 202 ][ 46 ],
   alphaCSR[ 202 ][ 47 ],
   alphaCSR[ 202 ][ 48 ],
   alphaCSR[ 202 ][ 49 ],
   alphaCSR[ 202 ][ 50 ],
   alphaCSR[ 202 ][ 51 ],
   alphaCSR[ 202 ][ 52 ],
   alphaCSR[ 202 ][ 53 ],
   alphaCSR[ 202 ][ 54 ],
   alphaCSR[ 202 ][ 55 ],
   alphaCSR[ 202 ][ 56 ],
   alphaCSR[ 202 ][ 57 ],
   alphaCSR[ 202 ][ 58 ],
   alphaCSR[ 202 ][ 59 ],
   alphaCSR[ 202 ][ 60 ],
   alphaCSR[ 202 ][ 61 ],
   alphaCSR[ 202 ][ 62 ],
   alphaCSR[ 202 ][ 63 ],
   alphaCSR[ 202 ][ 64 ],
   alphaCSR[ 202 ][ 65 ],
   alphaCSR[ 202 ][ 66 ],
   alphaCSR[ 202 ][ 67 ],
   alphaCSR[ 202 ][ 68 ],
   alphaCSR[ 202 ][ 69 ],
   alphaCSR[ 202 ][ 70 ],
   alphaCSR[ 202 ][ 71 ],
   alphaCSR[ 202 ][ 72 ],
   alphaCSR[ 202 ][ 73 ],
   alphaCSR[ 202 ][ 74 ],
   alphaCSR[ 202 ][ 75 ],
   alphaCSR[ 202 ][ 76 ],
   alphaCSR[ 202 ][ 77 ],
   alphaCSR[ 202 ][ 78 ],
   alphaCSR[ 202 ][ 79 ],
   alphaCSR[ 202 ][ 80 ],
   alphaCSR[ 202 ][ 81 ],
   alphaCSR[ 202 ][ 82 ],
   alphaCSR[ 202 ][ 83 ],
   alphaCSR[ 202 ][ 84 ],
   alphaCSR[ 202 ][ 85 ],
   alphaCSR[ 202 ][ 86 ],
   alphaCSR[ 202 ][ 87 ],
   alphaCSR[ 202 ][ 88 ],
   alphaCSR[ 202 ][ 89 ],
   alphaCSR[ 202 ][ 90 ],
   alphaCSR[ 202 ][ 91 ],
   alphaCSR[ 202 ][ 92 ],
   alphaCSR[ 202 ][ 93 ],
   alphaCSR[ 202 ][ 94 ],
   alphaCSR[ 202 ][ 95 ],
   alphaCSR[ 202 ][ 96 ],
   alphaCSR[ 202 ][ 97 ],
   alphaCSR[ 202 ][ 98 ],
   alphaCSR[ 202 ][ 99 ],
   alphaCSR[ 202 ][ 100 ],
   alphaCSR[ 202 ][ 101 ],
   alphaCSR[ 202 ][ 102 ],
   alphaCSR[ 202 ][ 103 ],
   alphaCSR[ 202 ][ 104 ],
   alphaCSR[ 202 ][ 105 ],
   alphaCSR[ 202 ][ 106 ],
   alphaCSR[ 202 ][ 107 ],
   alphaCSR[ 202 ][ 108 ],
   alphaCSR[ 202 ][ 109 ],
   alphaCSR[ 202 ][ 110 ],
   alphaCSR[ 202 ][ 111 ],
   alphaCSR[ 202 ][ 112 ],
   alphaCSR[ 202 ][ 113 ],
   alphaCSR[ 202 ][ 114 ],
   alphaCSR[ 202 ][ 115 ],
   alphaCSR[ 202 ][ 116 ],
   alphaCSR[ 202 ][ 117 ],
   alphaCSR[ 202 ][ 118 ],
   alphaCSR[ 202 ][ 119 ],
   alphaCSR[ 202 ][ 120 ],
   alphaCSR[ 202 ][ 121 ],
   alphaCSR[ 202 ][ 122 ],
   alphaCSR[ 202 ][ 123 ],
   alphaCSR[ 202 ][ 124 ],
   alphaCSR[ 202 ][ 125 ],
   alphaCSR[ 202 ][ 126 ],
   alphaCSR[ 202 ][ 127 ],
   alphaCSR[ 202 ][ 128 ],
   alphaCSR[ 202 ][ 129 ],
   alphaCSR[ 202 ][ 130 ],
   alphaCSR[ 202 ][ 131 ],
   alphaCSR[ 202 ][ 132 ],
   alphaCSR[ 202 ][ 133 ],
   alphaCSR[ 202 ][ 134 ],
   alphaCSR[ 202 ][ 135 ],
   alphaCSR[ 202 ][ 136 ],
   alphaCSR[ 202 ][ 137 ],
   alphaCSR[ 202 ][ 138 ],
   alphaCSR[ 202 ][ 139 ],
   alphaCSR[ 202 ][ 140 ],
   alphaCSR[ 202 ][ 141 ],
   alphaCSR[ 202 ][ 142 ],
   alphaCSR[ 202 ][ 143 ],
   alphaCSR[ 202 ][ 144 ],
   alphaCSR[ 202 ][ 145 ],
   alphaCSR[ 202 ][ 146 ],
   alphaCSR[ 202 ][ 147 ],
   alphaCSR[ 202 ][ 148 ],
   alphaCSR[ 202 ][ 149 ],
   alphaCSR[ 202 ][ 150 ],
   alphaCSR[ 202 ][ 151 ],
   alphaCSR[ 202 ][ 152 ],
   alphaCSR[ 202 ][ 153 ],
   alphaCSR[ 202 ][ 154 ],
   alphaCSR[ 202 ][ 155 ],
   alphaCSR[ 202 ][ 156 ],
   alphaCSR[ 202 ][ 157 ],
   alphaCSR[ 202 ][ 158 ],
   alphaCSR[ 202 ][ 159 ],
   alphaCSR[ 202 ][ 160 ],
   alphaCSR[ 202 ][ 161 ],
   alphaCSR[ 202 ][ 162 ],
   alphaCSR[ 202 ][ 163 ],
   alphaCSR[ 202 ][ 164 ],
   alphaCSR[ 202 ][ 165 ],
   alphaCSR[ 202 ][ 166 ],
   alphaCSR[ 202 ][ 167 ],
   alphaCSR[ 202 ][ 168 ],
   alphaCSR[ 202 ][ 169 ],
   alphaCSR[ 202 ][ 170 ],
   alphaCSR[ 202 ][ 171 ],
   alphaCSR[ 202 ][ 172 ],
   alphaCSR[ 202 ][ 173 ],
   alphaCSR[ 202 ][ 174 ],
   alphaCSR[ 202 ][ 175 ],
   alphaCSR[ 202 ][ 176 ],
   alphaCSR[ 202 ][ 177 ],
   alphaCSR[ 202 ][ 178 ],
   alphaCSR[ 202 ][ 179 ],
   alphaCSR[ 202 ][ 180 ],
   alphaCSR[ 202 ][ 181 ],
   alphaCSR[ 202 ][ 182 ],
   alphaCSR[ 202 ][ 183 ],
   alphaCSR[ 202 ][ 184 ],
   alphaCSR[ 202 ][ 185 ],
   alphaCSR[ 202 ][ 186 ],
   alphaCSR[ 202 ][ 187 ],
   alphaCSR[ 202 ][ 188 ],
   alphaCSR[ 202 ][ 189 ],
   alphaCSR[ 202 ][ 190 ],
   alphaCSR[ 202 ][ 191 ],
   alphaCSR[ 202 ][ 192 ],
   alphaCSR[ 202 ][ 193 ],
   alphaCSR[ 202 ][ 194 ],
   alphaCSR[ 202 ][ 195 ],
   alphaCSR[ 202 ][ 196 ],
   alphaCSR[ 202 ][ 197 ],
   alphaCSR[ 202 ][ 198 ],
   alphaCSR[ 202 ][ 199 ],
   alphaCSR[ 202 ][ 200 ],
   alphaCSR[ 202 ][ 201 ],
   alphaCSR[ 202 ][ 202 ],
   alphaCSR[ 202 ][ 203 ],
   alphaCSR[ 202 ][ 204 ],
   alphaCSR[ 202 ][ 205 ],
   alphaCSR[ 202 ][ 206 ],
   alphaCSR[ 202 ][ 207 ],
   alphaCSR[ 202 ][ 208 ],
   alphaCSR[ 202 ][ 209 ],
   alphaCSR[ 202 ][ 210 ],
   alphaCSR[ 202 ][ 211 ],
   alphaCSR[ 202 ][ 212 ],
   alphaCSR[ 202 ][ 213 ],
   alphaCSR[ 202 ][ 214 ],
   alphaCSR[ 202 ][ 215 ],
   alphaCSR[ 202 ][ 216 ],
   alphaCSR[ 202 ][ 217 ],
   alphaCSR[ 202 ][ 218 ],
   alphaCSR[ 202 ][ 219 ],
   alphaCSR[ 202 ][ 220 ],
   alphaCSR[ 202 ][ 221 ],
   alphaCSR[ 202 ][ 222 ],
   alphaCSR[ 202 ][ 223 ],
   alphaCSR[ 202 ][ 224 ],
   alphaCSR[ 202 ][ 225 ],
   alphaCSR[ 202 ][ 226 ],
   alphaCSR[ 202 ][ 227 ],
   alphaCSR[ 202 ][ 228 ],
   alphaCSR[ 202 ][ 229 ],
   alphaCSR[ 202 ][ 230 ],
   alphaCSR[ 202 ][ 231 ],
   alphaCSR[ 202 ][ 232 ],
   alphaCSR[ 202 ][ 233 ],
   alphaCSR[ 202 ][ 234 ],
   alphaCSR[ 202 ][ 235 ],
   alphaCSR[ 202 ][ 236 ],
   alphaCSR[ 202 ][ 237 ],
   alphaCSR[ 202 ][ 238 ],
   alphaCSR[ 202 ][ 239 ],
   alphaCSR[ 202 ][ 240 ],
   alphaCSR[ 202 ][ 241 ],
   alphaCSR[ 202 ][ 242 ],
   alphaCSR[ 202 ][ 243 ],
   alphaCSR[ 202 ][ 244 ],
   alphaCSR[ 202 ][ 245 ],
   alphaCSR[ 202 ][ 246 ],
   alphaCSR[ 202 ][ 247 ],
   alphaCSR[ 202 ][ 248 ],
   alphaCSR[ 202 ][ 249 ],
   alphaCSR[ 202 ][ 250 ],
   alphaCSR[ 202 ][ 251 ],
   alphaCSR[ 202 ][ 252 ],
   alphaCSR[ 202 ][ 253 ],
   alphaCSR[ 202 ][ 254 ],
   alphaCSR[ 202 ][ 255 ],
   alphaCSR[ 202 ][ 256 ],
   alphaCSR[ 202 ][ 257 ],
   alphaCSR[ 202 ][ 258 ],
   alphaCSR[ 202 ][ 259 ],
   alphaCSR[ 202 ][ 260 ],
   alphaCSR[ 202 ][ 261 ],
   alphaCSR[ 202 ][ 262 ],
   alphaCSR[ 202 ][ 263 ],
   alphaCSR[ 202 ][ 264 ],
   alphaCSR[ 202 ][ 265 ],
   alphaCSR[ 202 ][ 266 ],
   alphaCSR[ 202 ][ 267 ],
   alphaCSR[ 202 ][ 268 ],
   alphaCSR[ 202 ][ 269 ],
   alphaCSR[ 202 ][ 270 ],
   alphaCSR[ 202 ][ 271 ],
   alphaCSR[ 202 ][ 272 ],
   alphaCSR[ 202 ][ 273 ],
   alphaCSR[ 202 ][ 274 ],
   alphaCSR[ 202 ][ 275 ],
   alphaCSR[ 202 ][ 276 ],
   alphaCSR[ 202 ][ 277 ],
   alphaCSR[ 202 ][ 278 ],
   alphaCSR[ 202 ][ 279 ],
   alphaCSR[ 202 ][ 280 ],
   alphaCSR[ 202 ][ 281 ],
   alphaCSR[ 202 ][ 282 ],
   alphaCSR[ 202 ][ 283 ],
   alphaCSR[ 202 ][ 284 ],
   alphaCSR[ 202 ][ 285 ],
   alphaCSR[ 202 ][ 286 ],
   alphaCSR[ 202 ][ 287 ],
   alphaCSR[ 202 ][ 288 ],
   alphaCSR[ 202 ][ 289 ],
   alphaCSR[ 202 ][ 290 ],
   alphaCSR[ 202 ][ 291 ],
   alphaCSR[ 202 ][ 292 ],
   alphaCSR[ 202 ][ 293 ],
   alphaCSR[ 202 ][ 294 ],
   alphaCSR[ 202 ][ 295 ],
   alphaCSR[ 202 ][ 296 ],
   alphaCSR[ 202 ][ 297 ],
   alphaCSR[ 202 ][ 298 ],
   alphaCSR[ 202 ][ 299 ],
   alphaCSR[ 202 ][ 300 ],
   alphaCSR[ 202 ][ 301 ],
   alphaCSR[ 202 ][ 302 ],
   alphaCSR[ 202 ][ 303 ],
   alphaCSR[ 202 ][ 304 ],
   alphaCSR[ 202 ][ 305 ],
   alphaCSR[ 202 ][ 306 ],
   alphaCSR[ 202 ][ 307 ],
   alphaCSR[ 202 ][ 308 ],
   alphaCSR[ 202 ][ 309 ],
   alphaCSR[ 202 ][ 310 ],
   alphaCSR[ 202 ][ 311 ],
   alphaCSR[ 202 ][ 312 ],
   alphaCSR[ 202 ][ 313 ],
   alphaCSR[ 202 ][ 314 ],
   alphaCSR[ 202 ][ 315 ],
   alphaCSR[ 202 ][ 316 ],
   alphaCSR[ 202 ][ 317 ],
   alphaCSR[ 202 ][ 318 ],
   alphaCSR[ 202 ][ 319 ],
   alphaCSR[ 202 ][ 320 ],
   alphaCSR[ 202 ][ 321 ],
   alphaCSR[ 202 ][ 322 ],
   alphaCSR[ 202 ][ 323 ],
   alphaCSR[ 202 ][ 324 ],
   alphaCSR[ 202 ][ 325 ],
   alphaCSR[ 202 ][ 326 ],
   alphaCSR[ 202 ][ 327 ],
   alphaCSR[ 202 ][ 328 ],
   alphaCSR[ 202 ][ 329 ],
   alphaCSR[ 202 ][ 330 ],
   alphaCSR[ 202 ][ 331 ],
   alphaCSR[ 202 ][ 332 ],
   alphaCSR[ 202 ][ 333 ],
   alphaCSR[ 202 ][ 334 ],
   alphaCSR[ 202 ][ 335 ],
   alphaCSR[ 202 ][ 336 ],
   alphaCSR[ 202 ][ 337 ],
   alphaCSR[ 202 ][ 338 ],
   alphaCSR[ 202 ][ 339 ],
   alphaCSR[ 202 ][ 340 ],
   alphaCSR[ 202 ][ 341 ],
   alphaCSR[ 202 ][ 342 ],
   alphaCSR[ 202 ][ 343 ],
   alphaCSR[ 202 ][ 344 ],
   alphaCSR[ 202 ][ 345 ],
   alphaCSR[ 202 ][ 346 ],
   alphaCSR[ 202 ][ 347 ],
   alphaCSR[ 202 ][ 348 ],
   alphaCSR[ 202 ][ 349 ],
   alphaCSR[ 202 ][ 350 ],
   alphaCSR[ 202 ][ 351 ],
   alphaCSR[ 202 ][ 352 ],
   alphaCSR[ 202 ][ 353 ],
   alphaCSR[ 202 ][ 354 ],
   alphaCSR[ 202 ][ 355 ],
   alphaCSR[ 202 ][ 356 ],
   alphaCSR[ 202 ][ 357 ],
   alphaCSR[ 202 ][ 358 ],
   alphaCSR[ 202 ][ 359 ],
   alphaCSR[ 202 ][ 360 ],
   alphaCSR[ 202 ][ 361 ],
   alphaCSR[ 202 ][ 362 ],
   alphaCSR[ 202 ][ 363 ],
   alphaCSR[ 202 ][ 364 ],
   alphaCSR[ 202 ][ 365 ],
   alphaCSR[ 202 ][ 366 ],
   alphaCSR[ 202 ][ 367 ],
   alphaCSR[ 202 ][ 368 ],
   alphaCSR[ 202 ][ 369 ],
   alphaCSR[ 202 ][ 370 ],
   alphaCSR[ 202 ][ 371 ],
   alphaCSR[ 202 ][ 372 ],
   alphaCSR[ 202 ][ 373 ],
   alphaCSR[ 202 ][ 374 ],
   alphaCSR[ 202 ][ 375 ],
   alphaCSR[ 202 ][ 376 ],
   alphaCSR[ 202 ][ 377 ],
   alphaCSR[ 202 ][ 378 ],
   alphaCSR[ 202 ][ 379 ],
   alphaCSR[ 202 ][ 380 ],
   alphaCSR[ 202 ][ 381 ],
   alphaCSR[ 202 ][ 382 ],
   alphaCSR[ 202 ][ 383 ],
   alphaCSR[ 203 ][ 0 ],
   alphaCSR[ 203 ][ 1 ],
   alphaCSR[ 203 ][ 2 ],
   alphaCSR[ 203 ][ 3 ],
   alphaCSR[ 203 ][ 4 ],
   alphaCSR[ 203 ][ 5 ],
   alphaCSR[ 203 ][ 6 ],
   alphaCSR[ 203 ][ 7 ],
   alphaCSR[ 203 ][ 8 ],
   alphaCSR[ 203 ][ 9 ],
   alphaCSR[ 203 ][ 10 ],
   alphaCSR[ 203 ][ 11 ],
   alphaCSR[ 203 ][ 12 ],
   alphaCSR[ 203 ][ 13 ],
   alphaCSR[ 203 ][ 14 ],
   alphaCSR[ 203 ][ 15 ],
   alphaCSR[ 203 ][ 16 ],
   alphaCSR[ 203 ][ 17 ],
   alphaCSR[ 203 ][ 18 ],
   alphaCSR[ 203 ][ 19 ],
   alphaCSR[ 203 ][ 20 ],
   alphaCSR[ 203 ][ 21 ],
   alphaCSR[ 203 ][ 22 ],
   alphaCSR[ 203 ][ 23 ],
   alphaCSR[ 203 ][ 24 ],
   alphaCSR[ 203 ][ 25 ],
   alphaCSR[ 203 ][ 26 ],
   alphaCSR[ 203 ][ 27 ],
   alphaCSR[ 203 ][ 28 ],
   alphaCSR[ 203 ][ 29 ],
   alphaCSR[ 203 ][ 30 ],
   alphaCSR[ 203 ][ 31 ],
   alphaCSR[ 203 ][ 32 ],
   alphaCSR[ 203 ][ 33 ],
   alphaCSR[ 203 ][ 34 ],
   alphaCSR[ 203 ][ 35 ],
   alphaCSR[ 203 ][ 36 ],
   alphaCSR[ 203 ][ 37 ],
   alphaCSR[ 203 ][ 38 ],
   alphaCSR[ 203 ][ 39 ],
   alphaCSR[ 203 ][ 40 ],
   alphaCSR[ 203 ][ 41 ],
   alphaCSR[ 203 ][ 42 ],
   alphaCSR[ 203 ][ 43 ],
   alphaCSR[ 203 ][ 44 ],
   alphaCSR[ 203 ][ 45 ],
   alphaCSR[ 203 ][ 46 ],
   alphaCSR[ 203 ][ 47 ],
   alphaCSR[ 203 ][ 48 ],
   alphaCSR[ 203 ][ 49 ],
   alphaCSR[ 203 ][ 50 ],
   alphaCSR[ 203 ][ 51 ],
   alphaCSR[ 203 ][ 52 ],
   alphaCSR[ 203 ][ 53 ],
   alphaCSR[ 203 ][ 54 ],
   alphaCSR[ 203 ][ 55 ],
   alphaCSR[ 203 ][ 56 ],
   alphaCSR[ 203 ][ 57 ],
   alphaCSR[ 203 ][ 58 ],
   alphaCSR[ 203 ][ 59 ],
   alphaCSR[ 203 ][ 60 ],
   alphaCSR[ 203 ][ 61 ],
   alphaCSR[ 203 ][ 62 ],
   alphaCSR[ 203 ][ 63 ],
   alphaCSR[ 203 ][ 64 ],
   alphaCSR[ 203 ][ 65 ],
   alphaCSR[ 203 ][ 66 ],
   alphaCSR[ 203 ][ 67 ],
   alphaCSR[ 203 ][ 68 ],
   alphaCSR[ 203 ][ 69 ],
   alphaCSR[ 203 ][ 70 ],
   alphaCSR[ 203 ][ 71 ],
   alphaCSR[ 203 ][ 72 ],
   alphaCSR[ 203 ][ 73 ],
   alphaCSR[ 203 ][ 74 ],
   alphaCSR[ 203 ][ 75 ],
   alphaCSR[ 203 ][ 76 ],
   alphaCSR[ 203 ][ 77 ],
   alphaCSR[ 203 ][ 78 ],
   alphaCSR[ 203 ][ 79 ],
   alphaCSR[ 203 ][ 80 ],
   alphaCSR[ 203 ][ 81 ],
   alphaCSR[ 203 ][ 82 ],
   alphaCSR[ 203 ][ 83 ],
   alphaCSR[ 203 ][ 84 ],
   alphaCSR[ 203 ][ 85 ],
   alphaCSR[ 203 ][ 86 ],
   alphaCSR[ 203 ][ 87 ],
   alphaCSR[ 203 ][ 88 ],
   alphaCSR[ 203 ][ 89 ],
   alphaCSR[ 203 ][ 90 ],
   alphaCSR[ 203 ][ 91 ],
   alphaCSR[ 203 ][ 92 ],
   alphaCSR[ 203 ][ 93 ],
   alphaCSR[ 203 ][ 94 ],
   alphaCSR[ 203 ][ 95 ],
   alphaCSR[ 203 ][ 96 ],
   alphaCSR[ 203 ][ 97 ],
   alphaCSR[ 203 ][ 98 ],
   alphaCSR[ 203 ][ 99 ],
   alphaCSR[ 203 ][ 100 ],
   alphaCSR[ 203 ][ 101 ],
   alphaCSR[ 203 ][ 102 ],
   alphaCSR[ 203 ][ 103 ],
   alphaCSR[ 203 ][ 104 ],
   alphaCSR[ 203 ][ 105 ],
   alphaCSR[ 203 ][ 106 ],
   alphaCSR[ 203 ][ 107 ],
   alphaCSR[ 203 ][ 108 ],
   alphaCSR[ 203 ][ 109 ],
   alphaCSR[ 203 ][ 110 ],
   alphaCSR[ 203 ][ 111 ],
   alphaCSR[ 203 ][ 112 ],
   alphaCSR[ 203 ][ 113 ],
   alphaCSR[ 203 ][ 114 ],
   alphaCSR[ 203 ][ 115 ],
   alphaCSR[ 203 ][ 116 ],
   alphaCSR[ 203 ][ 117 ],
   alphaCSR[ 203 ][ 118 ],
   alphaCSR[ 203 ][ 119 ],
   alphaCSR[ 203 ][ 120 ],
   alphaCSR[ 203 ][ 121 ],
   alphaCSR[ 203 ][ 122 ],
   alphaCSR[ 203 ][ 123 ],
   alphaCSR[ 203 ][ 124 ],
   alphaCSR[ 203 ][ 125 ],
   alphaCSR[ 203 ][ 126 ],
   alphaCSR[ 203 ][ 127 ],
   alphaCSR[ 203 ][ 128 ],
   alphaCSR[ 203 ][ 129 ],
   alphaCSR[ 203 ][ 130 ],
   alphaCSR[ 203 ][ 131 ],
   alphaCSR[ 203 ][ 132 ],
   alphaCSR[ 203 ][ 133 ],
   alphaCSR[ 203 ][ 134 ],
   alphaCSR[ 203 ][ 135 ],
   alphaCSR[ 203 ][ 136 ],
   alphaCSR[ 203 ][ 137 ],
   alphaCSR[ 203 ][ 138 ],
   alphaCSR[ 203 ][ 139 ],
   alphaCSR[ 203 ][ 140 ],
   alphaCSR[ 203 ][ 141 ],
   alphaCSR[ 203 ][ 142 ],
   alphaCSR[ 203 ][ 143 ],
   alphaCSR[ 203 ][ 144 ],
   alphaCSR[ 203 ][ 145 ],
   alphaCSR[ 203 ][ 146 ],
   alphaCSR[ 203 ][ 147 ],
   alphaCSR[ 203 ][ 148 ],
   alphaCSR[ 203 ][ 149 ],
   alphaCSR[ 203 ][ 150 ],
   alphaCSR[ 203 ][ 151 ],
   alphaCSR[ 203 ][ 152 ],
   alphaCSR[ 203 ][ 153 ],
   alphaCSR[ 203 ][ 154 ],
   alphaCSR[ 203 ][ 155 ],
   alphaCSR[ 203 ][ 156 ],
   alphaCSR[ 203 ][ 157 ],
   alphaCSR[ 203 ][ 158 ],
   alphaCSR[ 203 ][ 159 ],
   alphaCSR[ 203 ][ 160 ],
   alphaCSR[ 203 ][ 161 ],
   alphaCSR[ 203 ][ 162 ],
   alphaCSR[ 203 ][ 163 ],
   alphaCSR[ 203 ][ 164 ],
   alphaCSR[ 203 ][ 165 ],
   alphaCSR[ 203 ][ 166 ],
   alphaCSR[ 203 ][ 167 ],
   alphaCSR[ 203 ][ 168 ],
   alphaCSR[ 203 ][ 169 ],
   alphaCSR[ 203 ][ 170 ],
   alphaCSR[ 203 ][ 171 ],
   alphaCSR[ 203 ][ 172 ],
   alphaCSR[ 203 ][ 173 ],
   alphaCSR[ 203 ][ 174 ],
   alphaCSR[ 203 ][ 175 ],
   alphaCSR[ 203 ][ 176 ],
   alphaCSR[ 203 ][ 177 ],
   alphaCSR[ 203 ][ 178 ],
   alphaCSR[ 203 ][ 179 ],
   alphaCSR[ 203 ][ 180 ],
   alphaCSR[ 203 ][ 181 ],
   alphaCSR[ 203 ][ 182 ],
   alphaCSR[ 203 ][ 183 ],
   alphaCSR[ 203 ][ 184 ],
   alphaCSR[ 203 ][ 185 ],
   alphaCSR[ 203 ][ 186 ],
   alphaCSR[ 203 ][ 187 ],
   alphaCSR[ 203 ][ 188 ],
   alphaCSR[ 203 ][ 189 ],
   alphaCSR[ 203 ][ 190 ],
   alphaCSR[ 203 ][ 191 ],
   alphaCSR[ 203 ][ 192 ],
   alphaCSR[ 203 ][ 193 ],
   alphaCSR[ 203 ][ 194 ],
   alphaCSR[ 203 ][ 195 ],
   alphaCSR[ 203 ][ 196 ],
   alphaCSR[ 203 ][ 197 ],
   alphaCSR[ 203 ][ 198 ],
   alphaCSR[ 203 ][ 199 ],
   alphaCSR[ 203 ][ 200 ],
   alphaCSR[ 203 ][ 201 ],
   alphaCSR[ 203 ][ 202 ],
   alphaCSR[ 203 ][ 203 ],
   alphaCSR[ 203 ][ 204 ],
   alphaCSR[ 203 ][ 205 ],
   alphaCSR[ 203 ][ 206 ],
   alphaCSR[ 203 ][ 207 ],
   alphaCSR[ 203 ][ 208 ],
   alphaCSR[ 203 ][ 209 ],
   alphaCSR[ 203 ][ 210 ],
   alphaCSR[ 203 ][ 211 ],
   alphaCSR[ 203 ][ 212 ],
   alphaCSR[ 203 ][ 213 ],
   alphaCSR[ 203 ][ 214 ],
   alphaCSR[ 203 ][ 215 ],
   alphaCSR[ 203 ][ 216 ],
   alphaCSR[ 203 ][ 217 ],
   alphaCSR[ 203 ][ 218 ],
   alphaCSR[ 203 ][ 219 ],
   alphaCSR[ 203 ][ 220 ],
   alphaCSR[ 203 ][ 221 ],
   alphaCSR[ 203 ][ 222 ],
   alphaCSR[ 203 ][ 223 ],
   alphaCSR[ 203 ][ 224 ],
   alphaCSR[ 203 ][ 225 ],
   alphaCSR[ 203 ][ 226 ],
   alphaCSR[ 203 ][ 227 ],
   alphaCSR[ 203 ][ 228 ],
   alphaCSR[ 203 ][ 229 ],
   alphaCSR[ 203 ][ 230 ],
   alphaCSR[ 203 ][ 231 ],
   alphaCSR[ 203 ][ 232 ],
   alphaCSR[ 203 ][ 233 ],
   alphaCSR[ 203 ][ 234 ],
   alphaCSR[ 203 ][ 235 ],
   alphaCSR[ 203 ][ 236 ],
   alphaCSR[ 203 ][ 237 ],
   alphaCSR[ 203 ][ 238 ],
   alphaCSR[ 203 ][ 239 ],
   alphaCSR[ 203 ][ 240 ],
   alphaCSR[ 203 ][ 241 ],
   alphaCSR[ 203 ][ 242 ],
   alphaCSR[ 203 ][ 243 ],
   alphaCSR[ 203 ][ 244 ],
   alphaCSR[ 203 ][ 245 ],
   alphaCSR[ 203 ][ 246 ],
   alphaCSR[ 203 ][ 247 ],
   alphaCSR[ 203 ][ 248 ],
   alphaCSR[ 203 ][ 249 ],
   alphaCSR[ 203 ][ 250 ],
   alphaCSR[ 203 ][ 251 ],
   alphaCSR[ 203 ][ 252 ],
   alphaCSR[ 203 ][ 253 ],
   alphaCSR[ 203 ][ 254 ],
   alphaCSR[ 203 ][ 255 ],
   alphaCSR[ 203 ][ 256 ],
   alphaCSR[ 203 ][ 257 ],
   alphaCSR[ 203 ][ 258 ],
   alphaCSR[ 203 ][ 259 ],
   alphaCSR[ 203 ][ 260 ],
   alphaCSR[ 203 ][ 261 ],
   alphaCSR[ 203 ][ 262 ],
   alphaCSR[ 203 ][ 263 ],
   alphaCSR[ 203 ][ 264 ],
   alphaCSR[ 203 ][ 265 ],
   alphaCSR[ 203 ][ 266 ],
   alphaCSR[ 203 ][ 267 ],
   alphaCSR[ 203 ][ 268 ],
   alphaCSR[ 203 ][ 269 ],
   alphaCSR[ 203 ][ 270 ],
   alphaCSR[ 203 ][ 271 ],
   alphaCSR[ 203 ][ 272 ],
   alphaCSR[ 203 ][ 273 ],
   alphaCSR[ 203 ][ 274 ],
   alphaCSR[ 203 ][ 275 ],
   alphaCSR[ 203 ][ 276 ],
   alphaCSR[ 203 ][ 277 ],
   alphaCSR[ 203 ][ 278 ],
   alphaCSR[ 203 ][ 279 ],
   alphaCSR[ 203 ][ 280 ],
   alphaCSR[ 203 ][ 281 ],
   alphaCSR[ 203 ][ 282 ],
   alphaCSR[ 203 ][ 283 ],
   alphaCSR[ 203 ][ 284 ],
   alphaCSR[ 203 ][ 285 ],
   alphaCSR[ 203 ][ 286 ],
   alphaCSR[ 203 ][ 287 ],
   alphaCSR[ 203 ][ 288 ],
   alphaCSR[ 203 ][ 289 ],
   alphaCSR[ 203 ][ 290 ],
   alphaCSR[ 203 ][ 291 ],
   alphaCSR[ 203 ][ 292 ],
   alphaCSR[ 203 ][ 293 ],
   alphaCSR[ 203 ][ 294 ],
   alphaCSR[ 203 ][ 295 ],
   alphaCSR[ 203 ][ 296 ],
   alphaCSR[ 203 ][ 297 ],
   alphaCSR[ 203 ][ 298 ],
   alphaCSR[ 203 ][ 299 ],
   alphaCSR[ 203 ][ 300 ],
   alphaCSR[ 203 ][ 301 ],
   alphaCSR[ 203 ][ 302 ],
   alphaCSR[ 203 ][ 303 ],
   alphaCSR[ 203 ][ 304 ],
   alphaCSR[ 203 ][ 305 ],
   alphaCSR[ 203 ][ 306 ],
   alphaCSR[ 203 ][ 307 ],
   alphaCSR[ 203 ][ 308 ],
   alphaCSR[ 203 ][ 309 ],
   alphaCSR[ 203 ][ 310 ],
   alphaCSR[ 203 ][ 311 ],
   alphaCSR[ 203 ][ 312 ],
   alphaCSR[ 203 ][ 313 ],
   alphaCSR[ 203 ][ 314 ],
   alphaCSR[ 203 ][ 315 ],
   alphaCSR[ 203 ][ 316 ],
   alphaCSR[ 203 ][ 317 ],
   alphaCSR[ 203 ][ 318 ],
   alphaCSR[ 203 ][ 319 ],
   alphaCSR[ 203 ][ 320 ],
   alphaCSR[ 203 ][ 321 ],
   alphaCSR[ 203 ][ 322 ],
   alphaCSR[ 203 ][ 323 ],
   alphaCSR[ 203 ][ 324 ],
   alphaCSR[ 203 ][ 325 ],
   alphaCSR[ 203 ][ 326 ],
   alphaCSR[ 203 ][ 327 ],
   alphaCSR[ 203 ][ 328 ],
   alphaCSR[ 203 ][ 329 ],
   alphaCSR[ 203 ][ 330 ],
   alphaCSR[ 203 ][ 331 ],
   alphaCSR[ 203 ][ 332 ],
   alphaCSR[ 203 ][ 333 ],
   alphaCSR[ 203 ][ 334 ],
   alphaCSR[ 203 ][ 335 ],
   alphaCSR[ 203 ][ 336 ],
   alphaCSR[ 203 ][ 337 ],
   alphaCSR[ 203 ][ 338 ],
   alphaCSR[ 203 ][ 339 ],
   alphaCSR[ 203 ][ 340 ],
   alphaCSR[ 203 ][ 341 ],
   alphaCSR[ 203 ][ 342 ],
   alphaCSR[ 203 ][ 343 ],
   alphaCSR[ 203 ][ 344 ],
   alphaCSR[ 203 ][ 345 ],
   alphaCSR[ 203 ][ 346 ],
   alphaCSR[ 203 ][ 347 ],
   alphaCSR[ 203 ][ 348 ],
   alphaCSR[ 203 ][ 349 ],
   alphaCSR[ 203 ][ 350 ],
   alphaCSR[ 203 ][ 351 ],
   alphaCSR[ 203 ][ 352 ],
   alphaCSR[ 203 ][ 353 ],
   alphaCSR[ 203 ][ 354 ],
   alphaCSR[ 203 ][ 355 ],
   alphaCSR[ 203 ][ 356 ],
   alphaCSR[ 203 ][ 357 ],
   alphaCSR[ 203 ][ 358 ],
   alphaCSR[ 203 ][ 359 ],
   alphaCSR[ 203 ][ 360 ],
   alphaCSR[ 203 ][ 361 ],
   alphaCSR[ 203 ][ 362 ],
   alphaCSR[ 203 ][ 363 ],
   alphaCSR[ 203 ][ 364 ],
   alphaCSR[ 203 ][ 365 ],
   alphaCSR[ 203 ][ 366 ],
   alphaCSR[ 203 ][ 367 ],
   alphaCSR[ 203 ][ 368 ],
   alphaCSR[ 203 ][ 369 ],
   alphaCSR[ 203 ][ 370 ],
   alphaCSR[ 203 ][ 371 ],
   alphaCSR[ 203 ][ 372 ],
   alphaCSR[ 203 ][ 373 ],
   alphaCSR[ 203 ][ 374 ],
   alphaCSR[ 203 ][ 375 ],
   alphaCSR[ 203 ][ 376 ],
   alphaCSR[ 203 ][ 377 ],
   alphaCSR[ 203 ][ 378 ],
   alphaCSR[ 203 ][ 379 ],
   alphaCSR[ 203 ][ 380 ],
   alphaCSR[ 203 ][ 381 ],
   alphaCSR[ 203 ][ 382 ],
   alphaCSR[ 203 ][ 383 ],
   alphaCSR[ 204 ][ 0 ],
   alphaCSR[ 204 ][ 1 ],
   alphaCSR[ 204 ][ 2 ],
   alphaCSR[ 204 ][ 3 ],
   alphaCSR[ 204 ][ 4 ],
   alphaCSR[ 204 ][ 5 ],
   alphaCSR[ 204 ][ 6 ],
   alphaCSR[ 204 ][ 7 ],
   alphaCSR[ 204 ][ 8 ],
   alphaCSR[ 204 ][ 9 ],
   alphaCSR[ 204 ][ 10 ],
   alphaCSR[ 204 ][ 11 ],
   alphaCSR[ 204 ][ 12 ],
   alphaCSR[ 204 ][ 13 ],
   alphaCSR[ 204 ][ 14 ],
   alphaCSR[ 204 ][ 15 ],
   alphaCSR[ 204 ][ 16 ],
   alphaCSR[ 204 ][ 17 ],
   alphaCSR[ 204 ][ 18 ],
   alphaCSR[ 204 ][ 19 ],
   alphaCSR[ 204 ][ 20 ],
   alphaCSR[ 204 ][ 21 ],
   alphaCSR[ 204 ][ 22 ],
   alphaCSR[ 204 ][ 23 ],
   alphaCSR[ 204 ][ 24 ],
   alphaCSR[ 204 ][ 25 ],
   alphaCSR[ 204 ][ 26 ],
   alphaCSR[ 204 ][ 27 ],
   alphaCSR[ 204 ][ 28 ],
   alphaCSR[ 204 ][ 29 ],
   alphaCSR[ 204 ][ 30 ],
   alphaCSR[ 204 ][ 31 ],
   alphaCSR[ 204 ][ 32 ],
   alphaCSR[ 204 ][ 33 ],
   alphaCSR[ 204 ][ 34 ],
   alphaCSR[ 204 ][ 35 ],
   alphaCSR[ 204 ][ 36 ],
   alphaCSR[ 204 ][ 37 ],
   alphaCSR[ 204 ][ 38 ],
   alphaCSR[ 204 ][ 39 ],
   alphaCSR[ 204 ][ 40 ],
   alphaCSR[ 204 ][ 41 ],
   alphaCSR[ 204 ][ 42 ],
   alphaCSR[ 204 ][ 43 ],
   alphaCSR[ 204 ][ 44 ],
   alphaCSR[ 204 ][ 45 ],
   alphaCSR[ 204 ][ 46 ],
   alphaCSR[ 204 ][ 47 ],
   alphaCSR[ 204 ][ 48 ],
   alphaCSR[ 204 ][ 49 ],
   alphaCSR[ 204 ][ 50 ],
   alphaCSR[ 204 ][ 51 ],
   alphaCSR[ 204 ][ 52 ],
   alphaCSR[ 204 ][ 53 ],
   alphaCSR[ 204 ][ 54 ],
   alphaCSR[ 204 ][ 55 ],
   alphaCSR[ 204 ][ 56 ],
   alphaCSR[ 204 ][ 57 ],
   alphaCSR[ 204 ][ 58 ],
   alphaCSR[ 204 ][ 59 ],
   alphaCSR[ 204 ][ 60 ],
   alphaCSR[ 204 ][ 61 ],
   alphaCSR[ 204 ][ 62 ],
   alphaCSR[ 204 ][ 63 ],
   alphaCSR[ 204 ][ 64 ],
   alphaCSR[ 204 ][ 65 ],
   alphaCSR[ 204 ][ 66 ],
   alphaCSR[ 204 ][ 67 ],
   alphaCSR[ 204 ][ 68 ],
   alphaCSR[ 204 ][ 69 ],
   alphaCSR[ 204 ][ 70 ],
   alphaCSR[ 204 ][ 71 ],
   alphaCSR[ 204 ][ 72 ],
   alphaCSR[ 204 ][ 73 ],
   alphaCSR[ 204 ][ 74 ],
   alphaCSR[ 204 ][ 75 ],
   alphaCSR[ 204 ][ 76 ],
   alphaCSR[ 204 ][ 77 ],
   alphaCSR[ 204 ][ 78 ],
   alphaCSR[ 204 ][ 79 ],
   alphaCSR[ 204 ][ 80 ],
   alphaCSR[ 204 ][ 81 ],
   alphaCSR[ 204 ][ 82 ],
   alphaCSR[ 204 ][ 83 ],
   alphaCSR[ 204 ][ 84 ],
   alphaCSR[ 204 ][ 85 ],
   alphaCSR[ 204 ][ 86 ],
   alphaCSR[ 204 ][ 87 ],
   alphaCSR[ 204 ][ 88 ],
   alphaCSR[ 204 ][ 89 ],
   alphaCSR[ 204 ][ 90 ],
   alphaCSR[ 204 ][ 91 ],
   alphaCSR[ 204 ][ 92 ],
   alphaCSR[ 204 ][ 93 ],
   alphaCSR[ 204 ][ 94 ],
   alphaCSR[ 204 ][ 95 ],
   alphaCSR[ 204 ][ 96 ],
   alphaCSR[ 204 ][ 97 ],
   alphaCSR[ 204 ][ 98 ],
   alphaCSR[ 204 ][ 99 ],
   alphaCSR[ 204 ][ 100 ],
   alphaCSR[ 204 ][ 101 ],
   alphaCSR[ 204 ][ 102 ],
   alphaCSR[ 204 ][ 103 ],
   alphaCSR[ 204 ][ 104 ],
   alphaCSR[ 204 ][ 105 ],
   alphaCSR[ 204 ][ 106 ],
   alphaCSR[ 204 ][ 107 ],
   alphaCSR[ 204 ][ 108 ],
   alphaCSR[ 204 ][ 109 ],
   alphaCSR[ 204 ][ 110 ],
   alphaCSR[ 204 ][ 111 ],
   alphaCSR[ 204 ][ 112 ],
   alphaCSR[ 204 ][ 113 ],
   alphaCSR[ 204 ][ 114 ],
   alphaCSR[ 204 ][ 115 ],
   alphaCSR[ 204 ][ 116 ],
   alphaCSR[ 204 ][ 117 ],
   alphaCSR[ 204 ][ 118 ],
   alphaCSR[ 204 ][ 119 ],
   alphaCSR[ 204 ][ 120 ],
   alphaCSR[ 204 ][ 121 ],
   alphaCSR[ 204 ][ 122 ],
   alphaCSR[ 204 ][ 123 ],
   alphaCSR[ 204 ][ 124 ],
   alphaCSR[ 204 ][ 125 ],
   alphaCSR[ 204 ][ 126 ],
   alphaCSR[ 204 ][ 127 ],
   alphaCSR[ 204 ][ 128 ],
   alphaCSR[ 204 ][ 129 ],
   alphaCSR[ 204 ][ 130 ],
   alphaCSR[ 204 ][ 131 ],
   alphaCSR[ 204 ][ 132 ],
   alphaCSR[ 204 ][ 133 ],
   alphaCSR[ 204 ][ 134 ],
   alphaCSR[ 204 ][ 135 ],
   alphaCSR[ 204 ][ 136 ],
   alphaCSR[ 204 ][ 137 ],
   alphaCSR[ 204 ][ 138 ],
   alphaCSR[ 204 ][ 139 ],
   alphaCSR[ 204 ][ 140 ],
   alphaCSR[ 204 ][ 141 ],
   alphaCSR[ 204 ][ 142 ],
   alphaCSR[ 204 ][ 143 ],
   alphaCSR[ 204 ][ 144 ],
   alphaCSR[ 204 ][ 145 ],
   alphaCSR[ 204 ][ 146 ],
   alphaCSR[ 204 ][ 147 ],
   alphaCSR[ 204 ][ 148 ],
   alphaCSR[ 204 ][ 149 ],
   alphaCSR[ 204 ][ 150 ],
   alphaCSR[ 204 ][ 151 ],
   alphaCSR[ 204 ][ 152 ],
   alphaCSR[ 204 ][ 153 ],
   alphaCSR[ 204 ][ 154 ],
   alphaCSR[ 204 ][ 155 ],
   alphaCSR[ 204 ][ 156 ],
   alphaCSR[ 204 ][ 157 ],
   alphaCSR[ 204 ][ 158 ],
   alphaCSR[ 204 ][ 159 ],
   alphaCSR[ 204 ][ 160 ],
   alphaCSR[ 204 ][ 161 ],
   alphaCSR[ 204 ][ 162 ],
   alphaCSR[ 204 ][ 163 ],
   alphaCSR[ 204 ][ 164 ],
   alphaCSR[ 204 ][ 165 ],
   alphaCSR[ 204 ][ 166 ],
   alphaCSR[ 204 ][ 167 ],
   alphaCSR[ 204 ][ 168 ],
   alphaCSR[ 204 ][ 169 ],
   alphaCSR[ 204 ][ 170 ],
   alphaCSR[ 204 ][ 171 ],
   alphaCSR[ 204 ][ 172 ],
   alphaCSR[ 204 ][ 173 ],
   alphaCSR[ 204 ][ 174 ],
   alphaCSR[ 204 ][ 175 ],
   alphaCSR[ 204 ][ 176 ],
   alphaCSR[ 204 ][ 177 ],
   alphaCSR[ 204 ][ 178 ],
   alphaCSR[ 204 ][ 179 ],
   alphaCSR[ 204 ][ 180 ],
   alphaCSR[ 204 ][ 181 ],
   alphaCSR[ 204 ][ 182 ],
   alphaCSR[ 204 ][ 183 ],
   alphaCSR[ 204 ][ 184 ],
   alphaCSR[ 204 ][ 185 ],
   alphaCSR[ 204 ][ 186 ],
   alphaCSR[ 204 ][ 187 ],
   alphaCSR[ 204 ][ 188 ],
   alphaCSR[ 204 ][ 189 ],
   alphaCSR[ 204 ][ 190 ],
   alphaCSR[ 204 ][ 191 ],
   alphaCSR[ 204 ][ 192 ],
   alphaCSR[ 204 ][ 193 ],
   alphaCSR[ 204 ][ 194 ],
   alphaCSR[ 204 ][ 195 ],
   alphaCSR[ 204 ][ 196 ],
   alphaCSR[ 204 ][ 197 ],
   alphaCSR[ 204 ][ 198 ],
   alphaCSR[ 204 ][ 199 ],
   alphaCSR[ 204 ][ 200 ],
   alphaCSR[ 204 ][ 201 ],
   alphaCSR[ 204 ][ 202 ],
   alphaCSR[ 204 ][ 203 ],
   alphaCSR[ 204 ][ 204 ],
   alphaCSR[ 204 ][ 205 ],
   alphaCSR[ 204 ][ 206 ],
   alphaCSR[ 204 ][ 207 ],
   alphaCSR[ 204 ][ 208 ],
   alphaCSR[ 204 ][ 209 ],
   alphaCSR[ 204 ][ 210 ],
   alphaCSR[ 204 ][ 211 ],
   alphaCSR[ 204 ][ 212 ],
   alphaCSR[ 204 ][ 213 ],
   alphaCSR[ 204 ][ 214 ],
   alphaCSR[ 204 ][ 215 ],
   alphaCSR[ 204 ][ 216 ],
   alphaCSR[ 204 ][ 217 ],
   alphaCSR[ 204 ][ 218 ],
   alphaCSR[ 204 ][ 219 ],
   alphaCSR[ 204 ][ 220 ],
   alphaCSR[ 204 ][ 221 ],
   alphaCSR[ 204 ][ 222 ],
   alphaCSR[ 204 ][ 223 ],
   alphaCSR[ 204 ][ 224 ],
   alphaCSR[ 204 ][ 225 ],
   alphaCSR[ 204 ][ 226 ],
   alphaCSR[ 204 ][ 227 ],
   alphaCSR[ 204 ][ 228 ],
   alphaCSR[ 204 ][ 229 ],
   alphaCSR[ 204 ][ 230 ],
   alphaCSR[ 204 ][ 231 ],
   alphaCSR[ 204 ][ 232 ],
   alphaCSR[ 204 ][ 233 ],
   alphaCSR[ 204 ][ 234 ],
   alphaCSR[ 204 ][ 235 ],
   alphaCSR[ 204 ][ 236 ],
   alphaCSR[ 204 ][ 237 ],
   alphaCSR[ 204 ][ 238 ],
   alphaCSR[ 204 ][ 239 ],
   alphaCSR[ 204 ][ 240 ],
   alphaCSR[ 204 ][ 241 ],
   alphaCSR[ 204 ][ 242 ],
   alphaCSR[ 204 ][ 243 ],
   alphaCSR[ 204 ][ 244 ],
   alphaCSR[ 204 ][ 245 ],
   alphaCSR[ 204 ][ 246 ],
   alphaCSR[ 204 ][ 247 ],
   alphaCSR[ 204 ][ 248 ],
   alphaCSR[ 204 ][ 249 ],
   alphaCSR[ 204 ][ 250 ],
   alphaCSR[ 204 ][ 251 ],
   alphaCSR[ 204 ][ 252 ],
   alphaCSR[ 204 ][ 253 ],
   alphaCSR[ 204 ][ 254 ],
   alphaCSR[ 204 ][ 255 ],
   alphaCSR[ 204 ][ 256 ],
   alphaCSR[ 204 ][ 257 ],
   alphaCSR[ 204 ][ 258 ],
   alphaCSR[ 204 ][ 259 ],
   alphaCSR[ 204 ][ 260 ],
   alphaCSR[ 204 ][ 261 ],
   alphaCSR[ 204 ][ 262 ],
   alphaCSR[ 204 ][ 263 ],
   alphaCSR[ 204 ][ 264 ],
   alphaCSR[ 204 ][ 265 ],
   alphaCSR[ 204 ][ 266 ],
   alphaCSR[ 204 ][ 267 ],
   alphaCSR[ 204 ][ 268 ],
   alphaCSR[ 204 ][ 269 ],
   alphaCSR[ 204 ][ 270 ],
   alphaCSR[ 204 ][ 271 ],
   alphaCSR[ 204 ][ 272 ],
   alphaCSR[ 204 ][ 273 ],
   alphaCSR[ 204 ][ 274 ],
   alphaCSR[ 204 ][ 275 ],
   alphaCSR[ 204 ][ 276 ],
   alphaCSR[ 204 ][ 277 ],
   alphaCSR[ 204 ][ 278 ],
   alphaCSR[ 204 ][ 279 ],
   alphaCSR[ 204 ][ 280 ],
   alphaCSR[ 204 ][ 281 ],
   alphaCSR[ 204 ][ 282 ],
   alphaCSR[ 204 ][ 283 ],
   alphaCSR[ 204 ][ 284 ],
   alphaCSR[ 204 ][ 285 ],
   alphaCSR[ 204 ][ 286 ],
   alphaCSR[ 204 ][ 287 ],
   alphaCSR[ 204 ][ 288 ],
   alphaCSR[ 204 ][ 289 ],
   alphaCSR[ 204 ][ 290 ],
   alphaCSR[ 204 ][ 291 ],
   alphaCSR[ 204 ][ 292 ],
   alphaCSR[ 204 ][ 293 ],
   alphaCSR[ 204 ][ 294 ],
   alphaCSR[ 204 ][ 295 ],
   alphaCSR[ 204 ][ 296 ],
   alphaCSR[ 204 ][ 297 ],
   alphaCSR[ 204 ][ 298 ],
   alphaCSR[ 204 ][ 299 ],
   alphaCSR[ 204 ][ 300 ],
   alphaCSR[ 204 ][ 301 ],
   alphaCSR[ 204 ][ 302 ],
   alphaCSR[ 204 ][ 303 ],
   alphaCSR[ 204 ][ 304 ],
   alphaCSR[ 204 ][ 305 ],
   alphaCSR[ 204 ][ 306 ],
   alphaCSR[ 204 ][ 307 ],
   alphaCSR[ 204 ][ 308 ],
   alphaCSR[ 204 ][ 309 ],
   alphaCSR[ 204 ][ 310 ],
   alphaCSR[ 204 ][ 311 ],
   alphaCSR[ 204 ][ 312 ],
   alphaCSR[ 204 ][ 313 ],
   alphaCSR[ 204 ][ 314 ],
   alphaCSR[ 204 ][ 315 ],
   alphaCSR[ 204 ][ 316 ],
   alphaCSR[ 204 ][ 317 ],
   alphaCSR[ 204 ][ 318 ],
   alphaCSR[ 204 ][ 319 ],
   alphaCSR[ 204 ][ 320 ],
   alphaCSR[ 204 ][ 321 ],
   alphaCSR[ 204 ][ 322 ],
   alphaCSR[ 204 ][ 323 ],
   alphaCSR[ 204 ][ 324 ],
   alphaCSR[ 204 ][ 325 ],
   alphaCSR[ 204 ][ 326 ],
   alphaCSR[ 204 ][ 327 ],
   alphaCSR[ 204 ][ 328 ],
   alphaCSR[ 204 ][ 329 ],
   alphaCSR[ 204 ][ 330 ],
   alphaCSR[ 204 ][ 331 ],
   alphaCSR[ 204 ][ 332 ],
   alphaCSR[ 204 ][ 333 ],
   alphaCSR[ 204 ][ 334 ],
   alphaCSR[ 204 ][ 335 ],
   alphaCSR[ 204 ][ 336 ],
   alphaCSR[ 204 ][ 337 ],
   alphaCSR[ 204 ][ 338 ],
   alphaCSR[ 204 ][ 339 ],
   alphaCSR[ 204 ][ 340 ],
   alphaCSR[ 204 ][ 341 ],
   alphaCSR[ 204 ][ 342 ],
   alphaCSR[ 204 ][ 343 ],
   alphaCSR[ 204 ][ 344 ],
   alphaCSR[ 204 ][ 345 ],
   alphaCSR[ 204 ][ 346 ],
   alphaCSR[ 204 ][ 347 ],
   alphaCSR[ 204 ][ 348 ],
   alphaCSR[ 204 ][ 349 ],
   alphaCSR[ 204 ][ 350 ],
   alphaCSR[ 204 ][ 351 ],
   alphaCSR[ 204 ][ 352 ],
   alphaCSR[ 204 ][ 353 ],
   alphaCSR[ 204 ][ 354 ],
   alphaCSR[ 204 ][ 355 ],
   alphaCSR[ 204 ][ 356 ],
   alphaCSR[ 204 ][ 357 ],
   alphaCSR[ 204 ][ 358 ],
   alphaCSR[ 204 ][ 359 ],
   alphaCSR[ 204 ][ 360 ],
   alphaCSR[ 204 ][ 361 ],
   alphaCSR[ 204 ][ 362 ],
   alphaCSR[ 204 ][ 363 ],
   alphaCSR[ 204 ][ 364 ],
   alphaCSR[ 204 ][ 365 ],
   alphaCSR[ 204 ][ 366 ],
   alphaCSR[ 204 ][ 367 ],
   alphaCSR[ 204 ][ 368 ],
   alphaCSR[ 204 ][ 369 ],
   alphaCSR[ 204 ][ 370 ],
   alphaCSR[ 204 ][ 371 ],
   alphaCSR[ 204 ][ 372 ],
   alphaCSR[ 204 ][ 373 ],
   alphaCSR[ 204 ][ 374 ],
   alphaCSR[ 204 ][ 375 ],
   alphaCSR[ 204 ][ 376 ],
   alphaCSR[ 204 ][ 377 ],
   alphaCSR[ 204 ][ 378 ],
   alphaCSR[ 204 ][ 379 ],
   alphaCSR[ 204 ][ 380 ],
   alphaCSR[ 204 ][ 381 ],
   alphaCSR[ 204 ][ 382 ],
   alphaCSR[ 204 ][ 383 ],
   alphaCSR[ 205 ][ 0 ],
   alphaCSR[ 205 ][ 1 ],
   alphaCSR[ 205 ][ 2 ],
   alphaCSR[ 205 ][ 3 ],
   alphaCSR[ 205 ][ 4 ],
   alphaCSR[ 205 ][ 5 ],
   alphaCSR[ 205 ][ 6 ],
   alphaCSR[ 205 ][ 7 ],
   alphaCSR[ 205 ][ 8 ],
   alphaCSR[ 205 ][ 9 ],
   alphaCSR[ 205 ][ 10 ],
   alphaCSR[ 205 ][ 11 ],
   alphaCSR[ 205 ][ 12 ],
   alphaCSR[ 205 ][ 13 ],
   alphaCSR[ 205 ][ 14 ],
   alphaCSR[ 205 ][ 15 ],
   alphaCSR[ 205 ][ 16 ],
   alphaCSR[ 205 ][ 17 ],
   alphaCSR[ 205 ][ 18 ],
   alphaCSR[ 205 ][ 19 ],
   alphaCSR[ 205 ][ 20 ],
   alphaCSR[ 205 ][ 21 ],
   alphaCSR[ 205 ][ 22 ],
   alphaCSR[ 205 ][ 23 ],
   alphaCSR[ 205 ][ 24 ],
   alphaCSR[ 205 ][ 25 ],
   alphaCSR[ 205 ][ 26 ],
   alphaCSR[ 205 ][ 27 ],
   alphaCSR[ 205 ][ 28 ],
   alphaCSR[ 205 ][ 29 ],
   alphaCSR[ 205 ][ 30 ],
   alphaCSR[ 205 ][ 31 ],
   alphaCSR[ 205 ][ 32 ],
   alphaCSR[ 205 ][ 33 ],
   alphaCSR[ 205 ][ 34 ],
   alphaCSR[ 205 ][ 35 ],
   alphaCSR[ 205 ][ 36 ],
   alphaCSR[ 205 ][ 37 ],
   alphaCSR[ 205 ][ 38 ],
   alphaCSR[ 205 ][ 39 ],
   alphaCSR[ 205 ][ 40 ],
   alphaCSR[ 205 ][ 41 ],
   alphaCSR[ 205 ][ 42 ],
   alphaCSR[ 205 ][ 43 ],
   alphaCSR[ 205 ][ 44 ],
   alphaCSR[ 205 ][ 45 ],
   alphaCSR[ 205 ][ 46 ],
   alphaCSR[ 205 ][ 47 ],
   alphaCSR[ 205 ][ 48 ],
   alphaCSR[ 205 ][ 49 ],
   alphaCSR[ 205 ][ 50 ],
   alphaCSR[ 205 ][ 51 ],
   alphaCSR[ 205 ][ 52 ],
   alphaCSR[ 205 ][ 53 ],
   alphaCSR[ 205 ][ 54 ],
   alphaCSR[ 205 ][ 55 ],
   alphaCSR[ 205 ][ 56 ],
   alphaCSR[ 205 ][ 57 ],
   alphaCSR[ 205 ][ 58 ],
   alphaCSR[ 205 ][ 59 ],
   alphaCSR[ 205 ][ 60 ],
   alphaCSR[ 205 ][ 61 ],
   alphaCSR[ 205 ][ 62 ],
   alphaCSR[ 205 ][ 63 ],
   alphaCSR[ 205 ][ 64 ],
   alphaCSR[ 205 ][ 65 ],
   alphaCSR[ 205 ][ 66 ],
   alphaCSR[ 205 ][ 67 ],
   alphaCSR[ 205 ][ 68 ],
   alphaCSR[ 205 ][ 69 ],
   alphaCSR[ 205 ][ 70 ],
   alphaCSR[ 205 ][ 71 ],
   alphaCSR[ 205 ][ 72 ],
   alphaCSR[ 205 ][ 73 ],
   alphaCSR[ 205 ][ 74 ],
   alphaCSR[ 205 ][ 75 ],
   alphaCSR[ 205 ][ 76 ],
   alphaCSR[ 205 ][ 77 ],
   alphaCSR[ 205 ][ 78 ],
   alphaCSR[ 205 ][ 79 ],
   alphaCSR[ 205 ][ 80 ],
   alphaCSR[ 205 ][ 81 ],
   alphaCSR[ 205 ][ 82 ],
   alphaCSR[ 205 ][ 83 ],
   alphaCSR[ 205 ][ 84 ],
   alphaCSR[ 205 ][ 85 ],
   alphaCSR[ 205 ][ 86 ],
   alphaCSR[ 205 ][ 87 ],
   alphaCSR[ 205 ][ 88 ],
   alphaCSR[ 205 ][ 89 ],
   alphaCSR[ 205 ][ 90 ],
   alphaCSR[ 205 ][ 91 ],
   alphaCSR[ 205 ][ 92 ],
   alphaCSR[ 205 ][ 93 ],
   alphaCSR[ 205 ][ 94 ],
   alphaCSR[ 205 ][ 95 ],
   alphaCSR[ 205 ][ 96 ],
   alphaCSR[ 205 ][ 97 ],
   alphaCSR[ 205 ][ 98 ],
   alphaCSR[ 205 ][ 99 ],
   alphaCSR[ 205 ][ 100 ],
   alphaCSR[ 205 ][ 101 ],
   alphaCSR[ 205 ][ 102 ],
   alphaCSR[ 205 ][ 103 ],
   alphaCSR[ 205 ][ 104 ],
   alphaCSR[ 205 ][ 105 ],
   alphaCSR[ 205 ][ 106 ],
   alphaCSR[ 205 ][ 107 ],
   alphaCSR[ 205 ][ 108 ],
   alphaCSR[ 205 ][ 109 ],
   alphaCSR[ 205 ][ 110 ],
   alphaCSR[ 205 ][ 111 ],
   alphaCSR[ 205 ][ 112 ],
   alphaCSR[ 205 ][ 113 ],
   alphaCSR[ 205 ][ 114 ],
   alphaCSR[ 205 ][ 115 ],
   alphaCSR[ 205 ][ 116 ],
   alphaCSR[ 205 ][ 117 ],
   alphaCSR[ 205 ][ 118 ],
   alphaCSR[ 205 ][ 119 ],
   alphaCSR[ 205 ][ 120 ],
   alphaCSR[ 205 ][ 121 ],
   alphaCSR[ 205 ][ 122 ],
   alphaCSR[ 205 ][ 123 ],
   alphaCSR[ 205 ][ 124 ],
   alphaCSR[ 205 ][ 125 ],
   alphaCSR[ 205 ][ 126 ],
   alphaCSR[ 205 ][ 127 ],
   alphaCSR[ 205 ][ 128 ],
   alphaCSR[ 205 ][ 129 ],
   alphaCSR[ 205 ][ 130 ],
   alphaCSR[ 205 ][ 131 ],
   alphaCSR[ 205 ][ 132 ],
   alphaCSR[ 205 ][ 133 ],
   alphaCSR[ 205 ][ 134 ],
   alphaCSR[ 205 ][ 135 ],
   alphaCSR[ 205 ][ 136 ],
   alphaCSR[ 205 ][ 137 ],
   alphaCSR[ 205 ][ 138 ],
   alphaCSR[ 205 ][ 139 ],
   alphaCSR[ 205 ][ 140 ],
   alphaCSR[ 205 ][ 141 ],
   alphaCSR[ 205 ][ 142 ],
   alphaCSR[ 205 ][ 143 ],
   alphaCSR[ 205 ][ 144 ],
   alphaCSR[ 205 ][ 145 ],
   alphaCSR[ 205 ][ 146 ],
   alphaCSR[ 205 ][ 147 ],
   alphaCSR[ 205 ][ 148 ],
   alphaCSR[ 205 ][ 149 ],
   alphaCSR[ 205 ][ 150 ],
   alphaCSR[ 205 ][ 151 ],
   alphaCSR[ 205 ][ 152 ],
   alphaCSR[ 205 ][ 153 ],
   alphaCSR[ 205 ][ 154 ],
   alphaCSR[ 205 ][ 155 ],
   alphaCSR[ 205 ][ 156 ],
   alphaCSR[ 205 ][ 157 ],
   alphaCSR[ 205 ][ 158 ],
   alphaCSR[ 205 ][ 159 ],
   alphaCSR[ 205 ][ 160 ],
   alphaCSR[ 205 ][ 161 ],
   alphaCSR[ 205 ][ 162 ],
   alphaCSR[ 205 ][ 163 ],
   alphaCSR[ 205 ][ 164 ],
   alphaCSR[ 205 ][ 165 ],
   alphaCSR[ 205 ][ 166 ],
   alphaCSR[ 205 ][ 167 ],
   alphaCSR[ 205 ][ 168 ],
   alphaCSR[ 205 ][ 169 ],
   alphaCSR[ 205 ][ 170 ],
   alphaCSR[ 205 ][ 171 ],
   alphaCSR[ 205 ][ 172 ],
   alphaCSR[ 205 ][ 173 ],
   alphaCSR[ 205 ][ 174 ],
   alphaCSR[ 205 ][ 175 ],
   alphaCSR[ 205 ][ 176 ],
   alphaCSR[ 205 ][ 177 ],
   alphaCSR[ 205 ][ 178 ],
   alphaCSR[ 205 ][ 179 ],
   alphaCSR[ 205 ][ 180 ],
   alphaCSR[ 205 ][ 181 ],
   alphaCSR[ 205 ][ 182 ],
   alphaCSR[ 205 ][ 183 ],
   alphaCSR[ 205 ][ 184 ],
   alphaCSR[ 205 ][ 185 ],
   alphaCSR[ 205 ][ 186 ],
   alphaCSR[ 205 ][ 187 ],
   alphaCSR[ 205 ][ 188 ],
   alphaCSR[ 205 ][ 189 ],
   alphaCSR[ 205 ][ 190 ],
   alphaCSR[ 205 ][ 191 ],
   alphaCSR[ 205 ][ 192 ],
   alphaCSR[ 205 ][ 193 ],
   alphaCSR[ 205 ][ 194 ],
   alphaCSR[ 205 ][ 195 ],
   alphaCSR[ 205 ][ 196 ],
   alphaCSR[ 205 ][ 197 ],
   alphaCSR[ 205 ][ 198 ],
   alphaCSR[ 205 ][ 199 ],
   alphaCSR[ 205 ][ 200 ],
   alphaCSR[ 205 ][ 201 ],
   alphaCSR[ 205 ][ 202 ],
   alphaCSR[ 205 ][ 203 ],
   alphaCSR[ 205 ][ 204 ],
   alphaCSR[ 205 ][ 205 ],
   alphaCSR[ 205 ][ 206 ],
   alphaCSR[ 205 ][ 207 ],
   alphaCSR[ 205 ][ 208 ],
   alphaCSR[ 205 ][ 209 ],
   alphaCSR[ 205 ][ 210 ],
   alphaCSR[ 205 ][ 211 ],
   alphaCSR[ 205 ][ 212 ],
   alphaCSR[ 205 ][ 213 ],
   alphaCSR[ 205 ][ 214 ],
   alphaCSR[ 205 ][ 215 ],
   alphaCSR[ 205 ][ 216 ],
   alphaCSR[ 205 ][ 217 ],
   alphaCSR[ 205 ][ 218 ],
   alphaCSR[ 205 ][ 219 ],
   alphaCSR[ 205 ][ 220 ],
   alphaCSR[ 205 ][ 221 ],
   alphaCSR[ 205 ][ 222 ],
   alphaCSR[ 205 ][ 223 ],
   alphaCSR[ 205 ][ 224 ],
   alphaCSR[ 205 ][ 225 ],
   alphaCSR[ 205 ][ 226 ],
   alphaCSR[ 205 ][ 227 ],
   alphaCSR[ 205 ][ 228 ],
   alphaCSR[ 205 ][ 229 ],
   alphaCSR[ 205 ][ 230 ],
   alphaCSR[ 205 ][ 231 ],
   alphaCSR[ 205 ][ 232 ],
   alphaCSR[ 205 ][ 233 ],
   alphaCSR[ 205 ][ 234 ],
   alphaCSR[ 205 ][ 235 ],
   alphaCSR[ 205 ][ 236 ],
   alphaCSR[ 205 ][ 237 ],
   alphaCSR[ 205 ][ 238 ],
   alphaCSR[ 205 ][ 239 ],
   alphaCSR[ 205 ][ 240 ],
   alphaCSR[ 205 ][ 241 ],
   alphaCSR[ 205 ][ 242 ],
   alphaCSR[ 205 ][ 243 ],
   alphaCSR[ 205 ][ 244 ],
   alphaCSR[ 205 ][ 245 ],
   alphaCSR[ 205 ][ 246 ],
   alphaCSR[ 205 ][ 247 ],
   alphaCSR[ 205 ][ 248 ],
   alphaCSR[ 205 ][ 249 ],
   alphaCSR[ 205 ][ 250 ],
   alphaCSR[ 205 ][ 251 ],
   alphaCSR[ 205 ][ 252 ],
   alphaCSR[ 205 ][ 253 ],
   alphaCSR[ 205 ][ 254 ],
   alphaCSR[ 205 ][ 255 ],
   alphaCSR[ 205 ][ 256 ],
   alphaCSR[ 205 ][ 257 ],
   alphaCSR[ 205 ][ 258 ],
   alphaCSR[ 205 ][ 259 ],
   alphaCSR[ 205 ][ 260 ],
   alphaCSR[ 205 ][ 261 ],
   alphaCSR[ 205 ][ 262 ],
   alphaCSR[ 205 ][ 263 ],
   alphaCSR[ 205 ][ 264 ],
   alphaCSR[ 205 ][ 265 ],
   alphaCSR[ 205 ][ 266 ],
   alphaCSR[ 205 ][ 267 ],
   alphaCSR[ 205 ][ 268 ],
   alphaCSR[ 205 ][ 269 ],
   alphaCSR[ 205 ][ 270 ],
   alphaCSR[ 205 ][ 271 ],
   alphaCSR[ 205 ][ 272 ],
   alphaCSR[ 205 ][ 273 ],
   alphaCSR[ 205 ][ 274 ],
   alphaCSR[ 205 ][ 275 ],
   alphaCSR[ 205 ][ 276 ],
   alphaCSR[ 205 ][ 277 ],
   alphaCSR[ 205 ][ 278 ],
   alphaCSR[ 205 ][ 279 ],
   alphaCSR[ 205 ][ 280 ],
   alphaCSR[ 205 ][ 281 ],
   alphaCSR[ 205 ][ 282 ],
   alphaCSR[ 205 ][ 283 ],
   alphaCSR[ 205 ][ 284 ],
   alphaCSR[ 205 ][ 285 ],
   alphaCSR[ 205 ][ 286 ],
   alphaCSR[ 205 ][ 287 ],
   alphaCSR[ 205 ][ 288 ],
   alphaCSR[ 205 ][ 289 ],
   alphaCSR[ 205 ][ 290 ],
   alphaCSR[ 205 ][ 291 ],
   alphaCSR[ 205 ][ 292 ],
   alphaCSR[ 205 ][ 293 ],
   alphaCSR[ 205 ][ 294 ],
   alphaCSR[ 205 ][ 295 ],
   alphaCSR[ 205 ][ 296 ],
   alphaCSR[ 205 ][ 297 ],
   alphaCSR[ 205 ][ 298 ],
   alphaCSR[ 205 ][ 299 ],
   alphaCSR[ 205 ][ 300 ],
   alphaCSR[ 205 ][ 301 ],
   alphaCSR[ 205 ][ 302 ],
   alphaCSR[ 205 ][ 303 ],
   alphaCSR[ 205 ][ 304 ],
   alphaCSR[ 205 ][ 305 ],
   alphaCSR[ 205 ][ 306 ],
   alphaCSR[ 205 ][ 307 ],
   alphaCSR[ 205 ][ 308 ],
   alphaCSR[ 205 ][ 309 ],
   alphaCSR[ 205 ][ 310 ],
   alphaCSR[ 205 ][ 311 ],
   alphaCSR[ 205 ][ 312 ],
   alphaCSR[ 205 ][ 313 ],
   alphaCSR[ 205 ][ 314 ],
   alphaCSR[ 205 ][ 315 ],
   alphaCSR[ 205 ][ 316 ],
   alphaCSR[ 205 ][ 317 ],
   alphaCSR[ 205 ][ 318 ],
   alphaCSR[ 205 ][ 319 ],
   alphaCSR[ 205 ][ 320 ],
   alphaCSR[ 205 ][ 321 ],
   alphaCSR[ 205 ][ 322 ],
   alphaCSR[ 205 ][ 323 ],
   alphaCSR[ 205 ][ 324 ],
   alphaCSR[ 205 ][ 325 ],
   alphaCSR[ 205 ][ 326 ],
   alphaCSR[ 205 ][ 327 ],
   alphaCSR[ 205 ][ 328 ],
   alphaCSR[ 205 ][ 329 ],
   alphaCSR[ 205 ][ 330 ],
   alphaCSR[ 205 ][ 331 ],
   alphaCSR[ 205 ][ 332 ],
   alphaCSR[ 205 ][ 333 ],
   alphaCSR[ 205 ][ 334 ],
   alphaCSR[ 205 ][ 335 ],
   alphaCSR[ 205 ][ 336 ],
   alphaCSR[ 205 ][ 337 ],
   alphaCSR[ 205 ][ 338 ],
   alphaCSR[ 205 ][ 339 ],
   alphaCSR[ 205 ][ 340 ],
   alphaCSR[ 205 ][ 341 ],
   alphaCSR[ 205 ][ 342 ],
   alphaCSR[ 205 ][ 343 ],
   alphaCSR[ 205 ][ 344 ],
   alphaCSR[ 205 ][ 345 ],
   alphaCSR[ 205 ][ 346 ],
   alphaCSR[ 205 ][ 347 ],
   alphaCSR[ 205 ][ 348 ],
   alphaCSR[ 205 ][ 349 ],
   alphaCSR[ 205 ][ 350 ],
   alphaCSR[ 205 ][ 351 ],
   alphaCSR[ 205 ][ 352 ],
   alphaCSR[ 205 ][ 353 ],
   alphaCSR[ 205 ][ 354 ],
   alphaCSR[ 205 ][ 355 ],
   alphaCSR[ 205 ][ 356 ],
   alphaCSR[ 205 ][ 357 ],
   alphaCSR[ 205 ][ 358 ],
   alphaCSR[ 205 ][ 359 ],
   alphaCSR[ 205 ][ 360 ],
   alphaCSR[ 205 ][ 361 ],
   alphaCSR[ 205 ][ 362 ],
   alphaCSR[ 205 ][ 363 ],
   alphaCSR[ 205 ][ 364 ],
   alphaCSR[ 205 ][ 365 ],
   alphaCSR[ 205 ][ 366 ],
   alphaCSR[ 205 ][ 367 ],
   alphaCSR[ 205 ][ 368 ],
   alphaCSR[ 205 ][ 369 ],
   alphaCSR[ 205 ][ 370 ],
   alphaCSR[ 205 ][ 371 ],
   alphaCSR[ 205 ][ 372 ],
   alphaCSR[ 205 ][ 373 ],
   alphaCSR[ 205 ][ 374 ],
   alphaCSR[ 205 ][ 375 ],
   alphaCSR[ 205 ][ 376 ],
   alphaCSR[ 205 ][ 377 ],
   alphaCSR[ 205 ][ 378 ],
   alphaCSR[ 205 ][ 379 ],
   alphaCSR[ 205 ][ 380 ],
   alphaCSR[ 205 ][ 381 ],
   alphaCSR[ 205 ][ 382 ],
   alphaCSR[ 205 ][ 383 ],
   alphaCSR[ 206 ][ 0 ],
   alphaCSR[ 206 ][ 1 ],
   alphaCSR[ 206 ][ 2 ],
   alphaCSR[ 206 ][ 3 ],
   alphaCSR[ 206 ][ 4 ],
   alphaCSR[ 206 ][ 5 ],
   alphaCSR[ 206 ][ 6 ],
   alphaCSR[ 206 ][ 7 ],
   alphaCSR[ 206 ][ 8 ],
   alphaCSR[ 206 ][ 9 ],
   alphaCSR[ 206 ][ 10 ],
   alphaCSR[ 206 ][ 11 ],
   alphaCSR[ 206 ][ 12 ],
   alphaCSR[ 206 ][ 13 ],
   alphaCSR[ 206 ][ 14 ],
   alphaCSR[ 206 ][ 15 ],
   alphaCSR[ 206 ][ 16 ],
   alphaCSR[ 206 ][ 17 ],
   alphaCSR[ 206 ][ 18 ],
   alphaCSR[ 206 ][ 19 ],
   alphaCSR[ 206 ][ 20 ],
   alphaCSR[ 206 ][ 21 ],
   alphaCSR[ 206 ][ 22 ],
   alphaCSR[ 206 ][ 23 ],
   alphaCSR[ 206 ][ 24 ],
   alphaCSR[ 206 ][ 25 ],
   alphaCSR[ 206 ][ 26 ],
   alphaCSR[ 206 ][ 27 ],
   alphaCSR[ 206 ][ 28 ],
   alphaCSR[ 206 ][ 29 ],
   alphaCSR[ 206 ][ 30 ],
   alphaCSR[ 206 ][ 31 ],
   alphaCSR[ 206 ][ 32 ],
   alphaCSR[ 206 ][ 33 ],
   alphaCSR[ 206 ][ 34 ],
   alphaCSR[ 206 ][ 35 ],
   alphaCSR[ 206 ][ 36 ],
   alphaCSR[ 206 ][ 37 ],
   alphaCSR[ 206 ][ 38 ],
   alphaCSR[ 206 ][ 39 ],
   alphaCSR[ 206 ][ 40 ],
   alphaCSR[ 206 ][ 41 ],
   alphaCSR[ 206 ][ 42 ],
   alphaCSR[ 206 ][ 43 ],
   alphaCSR[ 206 ][ 44 ],
   alphaCSR[ 206 ][ 45 ],
   alphaCSR[ 206 ][ 46 ],
   alphaCSR[ 206 ][ 47 ],
   alphaCSR[ 206 ][ 48 ],
   alphaCSR[ 206 ][ 49 ],
   alphaCSR[ 206 ][ 50 ],
   alphaCSR[ 206 ][ 51 ],
   alphaCSR[ 206 ][ 52 ],
   alphaCSR[ 206 ][ 53 ],
   alphaCSR[ 206 ][ 54 ],
   alphaCSR[ 206 ][ 55 ],
   alphaCSR[ 206 ][ 56 ],
   alphaCSR[ 206 ][ 57 ],
   alphaCSR[ 206 ][ 58 ],
   alphaCSR[ 206 ][ 59 ],
   alphaCSR[ 206 ][ 60 ],
   alphaCSR[ 206 ][ 61 ],
   alphaCSR[ 206 ][ 62 ],
   alphaCSR[ 206 ][ 63 ],
   alphaCSR[ 206 ][ 64 ],
   alphaCSR[ 206 ][ 65 ],
   alphaCSR[ 206 ][ 66 ],
   alphaCSR[ 206 ][ 67 ],
   alphaCSR[ 206 ][ 68 ],
   alphaCSR[ 206 ][ 69 ],
   alphaCSR[ 206 ][ 70 ],
   alphaCSR[ 206 ][ 71 ],
   alphaCSR[ 206 ][ 72 ],
   alphaCSR[ 206 ][ 73 ],
   alphaCSR[ 206 ][ 74 ],
   alphaCSR[ 206 ][ 75 ],
   alphaCSR[ 206 ][ 76 ],
   alphaCSR[ 206 ][ 77 ],
   alphaCSR[ 206 ][ 78 ],
   alphaCSR[ 206 ][ 79 ],
   alphaCSR[ 206 ][ 80 ],
   alphaCSR[ 206 ][ 81 ],
   alphaCSR[ 206 ][ 82 ],
   alphaCSR[ 206 ][ 83 ],
   alphaCSR[ 206 ][ 84 ],
   alphaCSR[ 206 ][ 85 ],
   alphaCSR[ 206 ][ 86 ],
   alphaCSR[ 206 ][ 87 ],
   alphaCSR[ 206 ][ 88 ],
   alphaCSR[ 206 ][ 89 ],
   alphaCSR[ 206 ][ 90 ],
   alphaCSR[ 206 ][ 91 ],
   alphaCSR[ 206 ][ 92 ],
   alphaCSR[ 206 ][ 93 ],
   alphaCSR[ 206 ][ 94 ],
   alphaCSR[ 206 ][ 95 ],
   alphaCSR[ 206 ][ 96 ],
   alphaCSR[ 206 ][ 97 ],
   alphaCSR[ 206 ][ 98 ],
   alphaCSR[ 206 ][ 99 ],
   alphaCSR[ 206 ][ 100 ],
   alphaCSR[ 206 ][ 101 ],
   alphaCSR[ 206 ][ 102 ],
   alphaCSR[ 206 ][ 103 ],
   alphaCSR[ 206 ][ 104 ],
   alphaCSR[ 206 ][ 105 ],
   alphaCSR[ 206 ][ 106 ],
   alphaCSR[ 206 ][ 107 ],
   alphaCSR[ 206 ][ 108 ],
   alphaCSR[ 206 ][ 109 ],
   alphaCSR[ 206 ][ 110 ],
   alphaCSR[ 206 ][ 111 ],
   alphaCSR[ 206 ][ 112 ],
   alphaCSR[ 206 ][ 113 ],
   alphaCSR[ 206 ][ 114 ],
   alphaCSR[ 206 ][ 115 ],
   alphaCSR[ 206 ][ 116 ],
   alphaCSR[ 206 ][ 117 ],
   alphaCSR[ 206 ][ 118 ],
   alphaCSR[ 206 ][ 119 ],
   alphaCSR[ 206 ][ 120 ],
   alphaCSR[ 206 ][ 121 ],
   alphaCSR[ 206 ][ 122 ],
   alphaCSR[ 206 ][ 123 ],
   alphaCSR[ 206 ][ 124 ],
   alphaCSR[ 206 ][ 125 ],
   alphaCSR[ 206 ][ 126 ],
   alphaCSR[ 206 ][ 127 ],
   alphaCSR[ 206 ][ 128 ],
   alphaCSR[ 206 ][ 129 ],
   alphaCSR[ 206 ][ 130 ],
   alphaCSR[ 206 ][ 131 ],
   alphaCSR[ 206 ][ 132 ],
   alphaCSR[ 206 ][ 133 ],
   alphaCSR[ 206 ][ 134 ],
   alphaCSR[ 206 ][ 135 ],
   alphaCSR[ 206 ][ 136 ],
   alphaCSR[ 206 ][ 137 ],
   alphaCSR[ 206 ][ 138 ],
   alphaCSR[ 206 ][ 139 ],
   alphaCSR[ 206 ][ 140 ],
   alphaCSR[ 206 ][ 141 ],
   alphaCSR[ 206 ][ 142 ],
   alphaCSR[ 206 ][ 143 ],
   alphaCSR[ 206 ][ 144 ],
   alphaCSR[ 206 ][ 145 ],
   alphaCSR[ 206 ][ 146 ],
   alphaCSR[ 206 ][ 147 ],
   alphaCSR[ 206 ][ 148 ],
   alphaCSR[ 206 ][ 149 ],
   alphaCSR[ 206 ][ 150 ],
   alphaCSR[ 206 ][ 151 ],
   alphaCSR[ 206 ][ 152 ],
   alphaCSR[ 206 ][ 153 ],
   alphaCSR[ 206 ][ 154 ],
   alphaCSR[ 206 ][ 155 ],
   alphaCSR[ 206 ][ 156 ],
   alphaCSR[ 206 ][ 157 ],
   alphaCSR[ 206 ][ 158 ],
   alphaCSR[ 206 ][ 159 ],
   alphaCSR[ 206 ][ 160 ],
   alphaCSR[ 206 ][ 161 ],
   alphaCSR[ 206 ][ 162 ],
   alphaCSR[ 206 ][ 163 ],
   alphaCSR[ 206 ][ 164 ],
   alphaCSR[ 206 ][ 165 ],
   alphaCSR[ 206 ][ 166 ],
   alphaCSR[ 206 ][ 167 ],
   alphaCSR[ 206 ][ 168 ],
   alphaCSR[ 206 ][ 169 ],
   alphaCSR[ 206 ][ 170 ],
   alphaCSR[ 206 ][ 171 ],
   alphaCSR[ 206 ][ 172 ],
   alphaCSR[ 206 ][ 173 ],
   alphaCSR[ 206 ][ 174 ],
   alphaCSR[ 206 ][ 175 ],
   alphaCSR[ 206 ][ 176 ],
   alphaCSR[ 206 ][ 177 ],
   alphaCSR[ 206 ][ 178 ],
   alphaCSR[ 206 ][ 179 ],
   alphaCSR[ 206 ][ 180 ],
   alphaCSR[ 206 ][ 181 ],
   alphaCSR[ 206 ][ 182 ],
   alphaCSR[ 206 ][ 183 ],
   alphaCSR[ 206 ][ 184 ],
   alphaCSR[ 206 ][ 185 ],
   alphaCSR[ 206 ][ 186 ],
   alphaCSR[ 206 ][ 187 ],
   alphaCSR[ 206 ][ 188 ],
   alphaCSR[ 206 ][ 189 ],
   alphaCSR[ 206 ][ 190 ],
   alphaCSR[ 206 ][ 191 ],
   alphaCSR[ 206 ][ 192 ],
   alphaCSR[ 206 ][ 193 ],
   alphaCSR[ 206 ][ 194 ],
   alphaCSR[ 206 ][ 195 ],
   alphaCSR[ 206 ][ 196 ],
   alphaCSR[ 206 ][ 197 ],
   alphaCSR[ 206 ][ 198 ],
   alphaCSR[ 206 ][ 199 ],
   alphaCSR[ 206 ][ 200 ],
   alphaCSR[ 206 ][ 201 ],
   alphaCSR[ 206 ][ 202 ],
   alphaCSR[ 206 ][ 203 ],
   alphaCSR[ 206 ][ 204 ],
   alphaCSR[ 206 ][ 205 ],
   alphaCSR[ 206 ][ 206 ],
   alphaCSR[ 206 ][ 207 ],
   alphaCSR[ 206 ][ 208 ],
   alphaCSR[ 206 ][ 209 ],
   alphaCSR[ 206 ][ 210 ],
   alphaCSR[ 206 ][ 211 ],
   alphaCSR[ 206 ][ 212 ],
   alphaCSR[ 206 ][ 213 ],
   alphaCSR[ 206 ][ 214 ],
   alphaCSR[ 206 ][ 215 ],
   alphaCSR[ 206 ][ 216 ],
   alphaCSR[ 206 ][ 217 ],
   alphaCSR[ 206 ][ 218 ],
   alphaCSR[ 206 ][ 219 ],
   alphaCSR[ 206 ][ 220 ],
   alphaCSR[ 206 ][ 221 ],
   alphaCSR[ 206 ][ 222 ],
   alphaCSR[ 206 ][ 223 ],
   alphaCSR[ 206 ][ 224 ],
   alphaCSR[ 206 ][ 225 ],
   alphaCSR[ 206 ][ 226 ],
   alphaCSR[ 206 ][ 227 ],
   alphaCSR[ 206 ][ 228 ],
   alphaCSR[ 206 ][ 229 ],
   alphaCSR[ 206 ][ 230 ],
   alphaCSR[ 206 ][ 231 ],
   alphaCSR[ 206 ][ 232 ],
   alphaCSR[ 206 ][ 233 ],
   alphaCSR[ 206 ][ 234 ],
   alphaCSR[ 206 ][ 235 ],
   alphaCSR[ 206 ][ 236 ],
   alphaCSR[ 206 ][ 237 ],
   alphaCSR[ 206 ][ 238 ],
   alphaCSR[ 206 ][ 239 ],
   alphaCSR[ 206 ][ 240 ],
   alphaCSR[ 206 ][ 241 ],
   alphaCSR[ 206 ][ 242 ],
   alphaCSR[ 206 ][ 243 ],
   alphaCSR[ 206 ][ 244 ],
   alphaCSR[ 206 ][ 245 ],
   alphaCSR[ 206 ][ 246 ],
   alphaCSR[ 206 ][ 247 ],
   alphaCSR[ 206 ][ 248 ],
   alphaCSR[ 206 ][ 249 ],
   alphaCSR[ 206 ][ 250 ],
   alphaCSR[ 206 ][ 251 ],
   alphaCSR[ 206 ][ 252 ],
   alphaCSR[ 206 ][ 253 ],
   alphaCSR[ 206 ][ 254 ],
   alphaCSR[ 206 ][ 255 ],
   alphaCSR[ 206 ][ 256 ],
   alphaCSR[ 206 ][ 257 ],
   alphaCSR[ 206 ][ 258 ],
   alphaCSR[ 206 ][ 259 ],
   alphaCSR[ 206 ][ 260 ],
   alphaCSR[ 206 ][ 261 ],
   alphaCSR[ 206 ][ 262 ],
   alphaCSR[ 206 ][ 263 ],
   alphaCSR[ 206 ][ 264 ],
   alphaCSR[ 206 ][ 265 ],
   alphaCSR[ 206 ][ 266 ],
   alphaCSR[ 206 ][ 267 ],
   alphaCSR[ 206 ][ 268 ],
   alphaCSR[ 206 ][ 269 ],
   alphaCSR[ 206 ][ 270 ],
   alphaCSR[ 206 ][ 271 ],
   alphaCSR[ 206 ][ 272 ],
   alphaCSR[ 206 ][ 273 ],
   alphaCSR[ 206 ][ 274 ],
   alphaCSR[ 206 ][ 275 ],
   alphaCSR[ 206 ][ 276 ],
   alphaCSR[ 206 ][ 277 ],
   alphaCSR[ 206 ][ 278 ],
   alphaCSR[ 206 ][ 279 ],
   alphaCSR[ 206 ][ 280 ],
   alphaCSR[ 206 ][ 281 ],
   alphaCSR[ 206 ][ 282 ],
   alphaCSR[ 206 ][ 283 ],
   alphaCSR[ 206 ][ 284 ],
   alphaCSR[ 206 ][ 285 ],
   alphaCSR[ 206 ][ 286 ],
   alphaCSR[ 206 ][ 287 ],
   alphaCSR[ 206 ][ 288 ],
   alphaCSR[ 206 ][ 289 ],
   alphaCSR[ 206 ][ 290 ],
   alphaCSR[ 206 ][ 291 ],
   alphaCSR[ 206 ][ 292 ],
   alphaCSR[ 206 ][ 293 ],
   alphaCSR[ 206 ][ 294 ],
   alphaCSR[ 206 ][ 295 ],
   alphaCSR[ 206 ][ 296 ],
   alphaCSR[ 206 ][ 297 ],
   alphaCSR[ 206 ][ 298 ],
   alphaCSR[ 206 ][ 299 ],
   alphaCSR[ 206 ][ 300 ],
   alphaCSR[ 206 ][ 301 ],
   alphaCSR[ 206 ][ 302 ],
   alphaCSR[ 206 ][ 303 ],
   alphaCSR[ 206 ][ 304 ],
   alphaCSR[ 206 ][ 305 ],
   alphaCSR[ 206 ][ 306 ],
   alphaCSR[ 206 ][ 307 ],
   alphaCSR[ 206 ][ 308 ],
   alphaCSR[ 206 ][ 309 ],
   alphaCSR[ 206 ][ 310 ],
   alphaCSR[ 206 ][ 311 ],
   alphaCSR[ 206 ][ 312 ],
   alphaCSR[ 206 ][ 313 ],
   alphaCSR[ 206 ][ 314 ],
   alphaCSR[ 206 ][ 315 ],
   alphaCSR[ 206 ][ 316 ],
   alphaCSR[ 206 ][ 317 ],
   alphaCSR[ 206 ][ 318 ],
   alphaCSR[ 206 ][ 319 ],
   alphaCSR[ 206 ][ 320 ],
   alphaCSR[ 206 ][ 321 ],
   alphaCSR[ 206 ][ 322 ],
   alphaCSR[ 206 ][ 323 ],
   alphaCSR[ 206 ][ 324 ],
   alphaCSR[ 206 ][ 325 ],
   alphaCSR[ 206 ][ 326 ],
   alphaCSR[ 206 ][ 327 ],
   alphaCSR[ 206 ][ 328 ],
   alphaCSR[ 206 ][ 329 ],
   alphaCSR[ 206 ][ 330 ],
   alphaCSR[ 206 ][ 331 ],
   alphaCSR[ 206 ][ 332 ],
   alphaCSR[ 206 ][ 333 ],
   alphaCSR[ 206 ][ 334 ],
   alphaCSR[ 206 ][ 335 ],
   alphaCSR[ 206 ][ 336 ],
   alphaCSR[ 206 ][ 337 ],
   alphaCSR[ 206 ][ 338 ],
   alphaCSR[ 206 ][ 339 ],
   alphaCSR[ 206 ][ 340 ],
   alphaCSR[ 206 ][ 341 ],
   alphaCSR[ 206 ][ 342 ],
   alphaCSR[ 206 ][ 343 ],
   alphaCSR[ 206 ][ 344 ],
   alphaCSR[ 206 ][ 345 ],
   alphaCSR[ 206 ][ 346 ],
   alphaCSR[ 206 ][ 347 ],
   alphaCSR[ 206 ][ 348 ],
   alphaCSR[ 206 ][ 349 ],
   alphaCSR[ 206 ][ 350 ],
   alphaCSR[ 206 ][ 351 ],
   alphaCSR[ 206 ][ 352 ],
   alphaCSR[ 206 ][ 353 ],
   alphaCSR[ 206 ][ 354 ],
   alphaCSR[ 206 ][ 355 ],
   alphaCSR[ 206 ][ 356 ],
   alphaCSR[ 206 ][ 357 ],
   alphaCSR[ 206 ][ 358 ],
   alphaCSR[ 206 ][ 359 ],
   alphaCSR[ 206 ][ 360 ],
   alphaCSR[ 206 ][ 361 ],
   alphaCSR[ 206 ][ 362 ],
   alphaCSR[ 206 ][ 363 ],
   alphaCSR[ 206 ][ 364 ],
   alphaCSR[ 206 ][ 365 ],
   alphaCSR[ 206 ][ 366 ],
   alphaCSR[ 206 ][ 367 ],
   alphaCSR[ 206 ][ 368 ],
   alphaCSR[ 206 ][ 369 ],
   alphaCSR[ 206 ][ 370 ],
   alphaCSR[ 206 ][ 371 ],
   alphaCSR[ 206 ][ 372 ],
   alphaCSR[ 206 ][ 373 ],
   alphaCSR[ 206 ][ 374 ],
   alphaCSR[ 206 ][ 375 ],
   alphaCSR[ 206 ][ 376 ],
   alphaCSR[ 206 ][ 377 ],
   alphaCSR[ 206 ][ 378 ],
   alphaCSR[ 206 ][ 379 ],
   alphaCSR[ 206 ][ 380 ],
   alphaCSR[ 206 ][ 381 ],
   alphaCSR[ 206 ][ 382 ],
   alphaCSR[ 206 ][ 383 ],
   alphaCSR[ 207 ][ 0 ],
   alphaCSR[ 207 ][ 1 ],
   alphaCSR[ 207 ][ 2 ],
   alphaCSR[ 207 ][ 3 ],
   alphaCSR[ 207 ][ 4 ],
   alphaCSR[ 207 ][ 5 ],
   alphaCSR[ 207 ][ 6 ],
   alphaCSR[ 207 ][ 7 ],
   alphaCSR[ 207 ][ 8 ],
   alphaCSR[ 207 ][ 9 ],
   alphaCSR[ 207 ][ 10 ],
   alphaCSR[ 207 ][ 11 ],
   alphaCSR[ 207 ][ 12 ],
   alphaCSR[ 207 ][ 13 ],
   alphaCSR[ 207 ][ 14 ],
   alphaCSR[ 207 ][ 15 ],
   alphaCSR[ 207 ][ 16 ],
   alphaCSR[ 207 ][ 17 ],
   alphaCSR[ 207 ][ 18 ],
   alphaCSR[ 207 ][ 19 ],
   alphaCSR[ 207 ][ 20 ],
   alphaCSR[ 207 ][ 21 ],
   alphaCSR[ 207 ][ 22 ],
   alphaCSR[ 207 ][ 23 ],
   alphaCSR[ 207 ][ 24 ],
   alphaCSR[ 207 ][ 25 ],
   alphaCSR[ 207 ][ 26 ],
   alphaCSR[ 207 ][ 27 ],
   alphaCSR[ 207 ][ 28 ],
   alphaCSR[ 207 ][ 29 ],
   alphaCSR[ 207 ][ 30 ],
   alphaCSR[ 207 ][ 31 ],
   alphaCSR[ 207 ][ 32 ],
   alphaCSR[ 207 ][ 33 ],
   alphaCSR[ 207 ][ 34 ],
   alphaCSR[ 207 ][ 35 ],
   alphaCSR[ 207 ][ 36 ],
   alphaCSR[ 207 ][ 37 ],
   alphaCSR[ 207 ][ 38 ],
   alphaCSR[ 207 ][ 39 ],
   alphaCSR[ 207 ][ 40 ],
   alphaCSR[ 207 ][ 41 ],
   alphaCSR[ 207 ][ 42 ],
   alphaCSR[ 207 ][ 43 ],
   alphaCSR[ 207 ][ 44 ],
   alphaCSR[ 207 ][ 45 ],
   alphaCSR[ 207 ][ 46 ],
   alphaCSR[ 207 ][ 47 ],
   alphaCSR[ 207 ][ 48 ],
   alphaCSR[ 207 ][ 49 ],
   alphaCSR[ 207 ][ 50 ],
   alphaCSR[ 207 ][ 51 ],
   alphaCSR[ 207 ][ 52 ],
   alphaCSR[ 207 ][ 53 ],
   alphaCSR[ 207 ][ 54 ],
   alphaCSR[ 207 ][ 55 ],
   alphaCSR[ 207 ][ 56 ],
   alphaCSR[ 207 ][ 57 ],
   alphaCSR[ 207 ][ 58 ],
   alphaCSR[ 207 ][ 59 ],
   alphaCSR[ 207 ][ 60 ],
   alphaCSR[ 207 ][ 61 ],
   alphaCSR[ 207 ][ 62 ],
   alphaCSR[ 207 ][ 63 ],
   alphaCSR[ 207 ][ 64 ],
   alphaCSR[ 207 ][ 65 ],
   alphaCSR[ 207 ][ 66 ],
   alphaCSR[ 207 ][ 67 ],
   alphaCSR[ 207 ][ 68 ],
   alphaCSR[ 207 ][ 69 ],
   alphaCSR[ 207 ][ 70 ],
   alphaCSR[ 207 ][ 71 ],
   alphaCSR[ 207 ][ 72 ],
   alphaCSR[ 207 ][ 73 ],
   alphaCSR[ 207 ][ 74 ],
   alphaCSR[ 207 ][ 75 ],
   alphaCSR[ 207 ][ 76 ],
   alphaCSR[ 207 ][ 77 ],
   alphaCSR[ 207 ][ 78 ],
   alphaCSR[ 207 ][ 79 ],
   alphaCSR[ 207 ][ 80 ],
   alphaCSR[ 207 ][ 81 ],
   alphaCSR[ 207 ][ 82 ],
   alphaCSR[ 207 ][ 83 ],
   alphaCSR[ 207 ][ 84 ],
   alphaCSR[ 207 ][ 85 ],
   alphaCSR[ 207 ][ 86 ],
   alphaCSR[ 207 ][ 87 ],
   alphaCSR[ 207 ][ 88 ],
   alphaCSR[ 207 ][ 89 ],
   alphaCSR[ 207 ][ 90 ],
   alphaCSR[ 207 ][ 91 ],
   alphaCSR[ 207 ][ 92 ],
   alphaCSR[ 207 ][ 93 ],
   alphaCSR[ 207 ][ 94 ],
   alphaCSR[ 207 ][ 95 ],
   alphaCSR[ 207 ][ 96 ],
   alphaCSR[ 207 ][ 97 ],
   alphaCSR[ 207 ][ 98 ],
   alphaCSR[ 207 ][ 99 ],
   alphaCSR[ 207 ][ 100 ],
   alphaCSR[ 207 ][ 101 ],
   alphaCSR[ 207 ][ 102 ],
   alphaCSR[ 207 ][ 103 ],
   alphaCSR[ 207 ][ 104 ],
   alphaCSR[ 207 ][ 105 ],
   alphaCSR[ 207 ][ 106 ],
   alphaCSR[ 207 ][ 107 ],
   alphaCSR[ 207 ][ 108 ],
   alphaCSR[ 207 ][ 109 ],
   alphaCSR[ 207 ][ 110 ],
   alphaCSR[ 207 ][ 111 ],
   alphaCSR[ 207 ][ 112 ],
   alphaCSR[ 207 ][ 113 ],
   alphaCSR[ 207 ][ 114 ],
   alphaCSR[ 207 ][ 115 ],
   alphaCSR[ 207 ][ 116 ],
   alphaCSR[ 207 ][ 117 ],
   alphaCSR[ 207 ][ 118 ],
   alphaCSR[ 207 ][ 119 ],
   alphaCSR[ 207 ][ 120 ],
   alphaCSR[ 207 ][ 121 ],
   alphaCSR[ 207 ][ 122 ],
   alphaCSR[ 207 ][ 123 ],
   alphaCSR[ 207 ][ 124 ],
   alphaCSR[ 207 ][ 125 ],
   alphaCSR[ 207 ][ 126 ],
   alphaCSR[ 207 ][ 127 ],
   alphaCSR[ 207 ][ 128 ],
   alphaCSR[ 207 ][ 129 ],
   alphaCSR[ 207 ][ 130 ],
   alphaCSR[ 207 ][ 131 ],
   alphaCSR[ 207 ][ 132 ],
   alphaCSR[ 207 ][ 133 ],
   alphaCSR[ 207 ][ 134 ],
   alphaCSR[ 207 ][ 135 ],
   alphaCSR[ 207 ][ 136 ],
   alphaCSR[ 207 ][ 137 ],
   alphaCSR[ 207 ][ 138 ],
   alphaCSR[ 207 ][ 139 ],
   alphaCSR[ 207 ][ 140 ],
   alphaCSR[ 207 ][ 141 ],
   alphaCSR[ 207 ][ 142 ],
   alphaCSR[ 207 ][ 143 ],
   alphaCSR[ 207 ][ 144 ],
   alphaCSR[ 207 ][ 145 ],
   alphaCSR[ 207 ][ 146 ],
   alphaCSR[ 207 ][ 147 ],
   alphaCSR[ 207 ][ 148 ],
   alphaCSR[ 207 ][ 149 ],
   alphaCSR[ 207 ][ 150 ],
   alphaCSR[ 207 ][ 151 ],
   alphaCSR[ 207 ][ 152 ],
   alphaCSR[ 207 ][ 153 ],
   alphaCSR[ 207 ][ 154 ],
   alphaCSR[ 207 ][ 155 ],
   alphaCSR[ 207 ][ 156 ],
   alphaCSR[ 207 ][ 157 ],
   alphaCSR[ 207 ][ 158 ],
   alphaCSR[ 207 ][ 159 ],
   alphaCSR[ 207 ][ 160 ],
   alphaCSR[ 207 ][ 161 ],
   alphaCSR[ 207 ][ 162 ],
   alphaCSR[ 207 ][ 163 ],
   alphaCSR[ 207 ][ 164 ],
   alphaCSR[ 207 ][ 165 ],
   alphaCSR[ 207 ][ 166 ],
   alphaCSR[ 207 ][ 167 ],
   alphaCSR[ 207 ][ 168 ],
   alphaCSR[ 207 ][ 169 ],
   alphaCSR[ 207 ][ 170 ],
   alphaCSR[ 207 ][ 171 ],
   alphaCSR[ 207 ][ 172 ],
   alphaCSR[ 207 ][ 173 ],
   alphaCSR[ 207 ][ 174 ],
   alphaCSR[ 207 ][ 175 ],
   alphaCSR[ 207 ][ 176 ],
   alphaCSR[ 207 ][ 177 ],
   alphaCSR[ 207 ][ 178 ],
   alphaCSR[ 207 ][ 179 ],
   alphaCSR[ 207 ][ 180 ],
   alphaCSR[ 207 ][ 181 ],
   alphaCSR[ 207 ][ 182 ],
   alphaCSR[ 207 ][ 183 ],
   alphaCSR[ 207 ][ 184 ],
   alphaCSR[ 207 ][ 185 ],
   alphaCSR[ 207 ][ 186 ],
   alphaCSR[ 207 ][ 187 ],
   alphaCSR[ 207 ][ 188 ],
   alphaCSR[ 207 ][ 189 ],
   alphaCSR[ 207 ][ 190 ],
   alphaCSR[ 207 ][ 191 ],
   alphaCSR[ 207 ][ 192 ],
   alphaCSR[ 207 ][ 193 ],
   alphaCSR[ 207 ][ 194 ],
   alphaCSR[ 207 ][ 195 ],
   alphaCSR[ 207 ][ 196 ],
   alphaCSR[ 207 ][ 197 ],
   alphaCSR[ 207 ][ 198 ],
   alphaCSR[ 207 ][ 199 ],
   alphaCSR[ 207 ][ 200 ],
   alphaCSR[ 207 ][ 201 ],
   alphaCSR[ 207 ][ 202 ],
   alphaCSR[ 207 ][ 203 ],
   alphaCSR[ 207 ][ 204 ],
   alphaCSR[ 207 ][ 205 ],
   alphaCSR[ 207 ][ 206 ],
   alphaCSR[ 207 ][ 207 ],
   alphaCSR[ 207 ][ 208 ],
   alphaCSR[ 207 ][ 209 ],
   alphaCSR[ 207 ][ 210 ],
   alphaCSR[ 207 ][ 211 ],
   alphaCSR[ 207 ][ 212 ],
   alphaCSR[ 207 ][ 213 ],
   alphaCSR[ 207 ][ 214 ],
   alphaCSR[ 207 ][ 215 ],
   alphaCSR[ 207 ][ 216 ],
   alphaCSR[ 207 ][ 217 ],
   alphaCSR[ 207 ][ 218 ],
   alphaCSR[ 207 ][ 219 ],
   alphaCSR[ 207 ][ 220 ],
   alphaCSR[ 207 ][ 221 ],
   alphaCSR[ 207 ][ 222 ],
   alphaCSR[ 207 ][ 223 ],
   alphaCSR[ 207 ][ 224 ],
   alphaCSR[ 207 ][ 225 ],
   alphaCSR[ 207 ][ 226 ],
   alphaCSR[ 207 ][ 227 ],
   alphaCSR[ 207 ][ 228 ],
   alphaCSR[ 207 ][ 229 ],
   alphaCSR[ 207 ][ 230 ],
   alphaCSR[ 207 ][ 231 ],
   alphaCSR[ 207 ][ 232 ],
   alphaCSR[ 207 ][ 233 ],
   alphaCSR[ 207 ][ 234 ],
   alphaCSR[ 207 ][ 235 ],
   alphaCSR[ 207 ][ 236 ],
   alphaCSR[ 207 ][ 237 ],
   alphaCSR[ 207 ][ 238 ],
   alphaCSR[ 207 ][ 239 ],
   alphaCSR[ 207 ][ 240 ],
   alphaCSR[ 207 ][ 241 ],
   alphaCSR[ 207 ][ 242 ],
   alphaCSR[ 207 ][ 243 ],
   alphaCSR[ 207 ][ 244 ],
   alphaCSR[ 207 ][ 245 ],
   alphaCSR[ 207 ][ 246 ],
   alphaCSR[ 207 ][ 247 ],
   alphaCSR[ 207 ][ 248 ],
   alphaCSR[ 207 ][ 249 ],
   alphaCSR[ 207 ][ 250 ],
   alphaCSR[ 207 ][ 251 ],
   alphaCSR[ 207 ][ 252 ],
   alphaCSR[ 207 ][ 253 ],
   alphaCSR[ 207 ][ 254 ],
   alphaCSR[ 207 ][ 255 ],
   alphaCSR[ 207 ][ 256 ],
   alphaCSR[ 207 ][ 257 ],
   alphaCSR[ 207 ][ 258 ],
   alphaCSR[ 207 ][ 259 ],
   alphaCSR[ 207 ][ 260 ],
   alphaCSR[ 207 ][ 261 ],
   alphaCSR[ 207 ][ 262 ],
   alphaCSR[ 207 ][ 263 ],
   alphaCSR[ 207 ][ 264 ],
   alphaCSR[ 207 ][ 265 ],
   alphaCSR[ 207 ][ 266 ],
   alphaCSR[ 207 ][ 267 ],
   alphaCSR[ 207 ][ 268 ],
   alphaCSR[ 207 ][ 269 ],
   alphaCSR[ 207 ][ 270 ],
   alphaCSR[ 207 ][ 271 ],
   alphaCSR[ 207 ][ 272 ],
   alphaCSR[ 207 ][ 273 ],
   alphaCSR[ 207 ][ 274 ],
   alphaCSR[ 207 ][ 275 ],
   alphaCSR[ 207 ][ 276 ],
   alphaCSR[ 207 ][ 277 ],
   alphaCSR[ 207 ][ 278 ],
   alphaCSR[ 207 ][ 279 ],
   alphaCSR[ 207 ][ 280 ],
   alphaCSR[ 207 ][ 281 ],
   alphaCSR[ 207 ][ 282 ],
   alphaCSR[ 207 ][ 283 ],
   alphaCSR[ 207 ][ 284 ],
   alphaCSR[ 207 ][ 285 ],
   alphaCSR[ 207 ][ 286 ],
   alphaCSR[ 207 ][ 287 ],
   alphaCSR[ 207 ][ 288 ],
   alphaCSR[ 207 ][ 289 ],
   alphaCSR[ 207 ][ 290 ],
   alphaCSR[ 207 ][ 291 ],
   alphaCSR[ 207 ][ 292 ],
   alphaCSR[ 207 ][ 293 ],
   alphaCSR[ 207 ][ 294 ],
   alphaCSR[ 207 ][ 295 ],
   alphaCSR[ 207 ][ 296 ],
   alphaCSR[ 207 ][ 297 ],
   alphaCSR[ 207 ][ 298 ],
   alphaCSR[ 207 ][ 299 ],
   alphaCSR[ 207 ][ 300 ],
   alphaCSR[ 207 ][ 301 ],
   alphaCSR[ 207 ][ 302 ],
   alphaCSR[ 207 ][ 303 ],
   alphaCSR[ 207 ][ 304 ],
   alphaCSR[ 207 ][ 305 ],
   alphaCSR[ 207 ][ 306 ],
   alphaCSR[ 207 ][ 307 ],
   alphaCSR[ 207 ][ 308 ],
   alphaCSR[ 207 ][ 309 ],
   alphaCSR[ 207 ][ 310 ],
   alphaCSR[ 207 ][ 311 ],
   alphaCSR[ 207 ][ 312 ],
   alphaCSR[ 207 ][ 313 ],
   alphaCSR[ 207 ][ 314 ],
   alphaCSR[ 207 ][ 315 ],
   alphaCSR[ 207 ][ 316 ],
   alphaCSR[ 207 ][ 317 ],
   alphaCSR[ 207 ][ 318 ],
   alphaCSR[ 207 ][ 319 ],
   alphaCSR[ 207 ][ 320 ],
   alphaCSR[ 207 ][ 321 ],
   alphaCSR[ 207 ][ 322 ],
   alphaCSR[ 207 ][ 323 ],
   alphaCSR[ 207 ][ 324 ],
   alphaCSR[ 207 ][ 325 ],
   alphaCSR[ 207 ][ 326 ],
   alphaCSR[ 207 ][ 327 ],
   alphaCSR[ 207 ][ 328 ],
   alphaCSR[ 207 ][ 329 ],
   alphaCSR[ 207 ][ 330 ],
   alphaCSR[ 207 ][ 331 ],
   alphaCSR[ 207 ][ 332 ],
   alphaCSR[ 207 ][ 333 ],
   alphaCSR[ 207 ][ 334 ],
   alphaCSR[ 207 ][ 335 ],
   alphaCSR[ 207 ][ 336 ],
   alphaCSR[ 207 ][ 337 ],
   alphaCSR[ 207 ][ 338 ],
   alphaCSR[ 207 ][ 339 ],
   alphaCSR[ 207 ][ 340 ],
   alphaCSR[ 207 ][ 341 ],
   alphaCSR[ 207 ][ 342 ],
   alphaCSR[ 207 ][ 343 ],
   alphaCSR[ 207 ][ 344 ],
   alphaCSR[ 207 ][ 345 ],
   alphaCSR[ 207 ][ 346 ],
   alphaCSR[ 207 ][ 347 ],
   alphaCSR[ 207 ][ 348 ],
   alphaCSR[ 207 ][ 349 ],
   alphaCSR[ 207 ][ 350 ],
   alphaCSR[ 207 ][ 351 ],
   alphaCSR[ 207 ][ 352 ],
   alphaCSR[ 207 ][ 353 ],
   alphaCSR[ 207 ][ 354 ],
   alphaCSR[ 207 ][ 355 ],
   alphaCSR[ 207 ][ 356 ],
   alphaCSR[ 207 ][ 357 ],
   alphaCSR[ 207 ][ 358 ],
   alphaCSR[ 207 ][ 359 ],
   alphaCSR[ 207 ][ 360 ],
   alphaCSR[ 207 ][ 361 ],
   alphaCSR[ 207 ][ 362 ],
   alphaCSR[ 207 ][ 363 ],
   alphaCSR[ 207 ][ 364 ],
   alphaCSR[ 207 ][ 365 ],
   alphaCSR[ 207 ][ 366 ],
   alphaCSR[ 207 ][ 367 ],
   alphaCSR[ 207 ][ 368 ],
   alphaCSR[ 207 ][ 369 ],
   alphaCSR[ 207 ][ 370 ],
   alphaCSR[ 207 ][ 371 ],
   alphaCSR[ 207 ][ 372 ],
   alphaCSR[ 207 ][ 373 ],
   alphaCSR[ 207 ][ 374 ],
   alphaCSR[ 207 ][ 375 ],
   alphaCSR[ 207 ][ 376 ],
   alphaCSR[ 207 ][ 377 ],
   alphaCSR[ 207 ][ 378 ],
   alphaCSR[ 207 ][ 379 ],
   alphaCSR[ 207 ][ 380 ],
   alphaCSR[ 207 ][ 381 ],
   alphaCSR[ 207 ][ 382 ],
   alphaCSR[ 207 ][ 383 ],
   alphaCSR[ 208 ][ 0 ],
   alphaCSR[ 208 ][ 1 ],
   alphaCSR[ 208 ][ 2 ],
   alphaCSR[ 208 ][ 3 ],
   alphaCSR[ 208 ][ 4 ],
   alphaCSR[ 208 ][ 5 ],
   alphaCSR[ 208 ][ 6 ],
   alphaCSR[ 208 ][ 7 ],
   alphaCSR[ 208 ][ 8 ],
   alphaCSR[ 208 ][ 9 ],
   alphaCSR[ 208 ][ 10 ],
   alphaCSR[ 208 ][ 11 ],
   alphaCSR[ 208 ][ 12 ],
   alphaCSR[ 208 ][ 13 ],
   alphaCSR[ 208 ][ 14 ],
   alphaCSR[ 208 ][ 15 ],
   alphaCSR[ 208 ][ 16 ],
   alphaCSR[ 208 ][ 17 ],
   alphaCSR[ 208 ][ 18 ],
   alphaCSR[ 208 ][ 19 ],
   alphaCSR[ 208 ][ 20 ],
   alphaCSR[ 208 ][ 21 ],
   alphaCSR[ 208 ][ 22 ],
   alphaCSR[ 208 ][ 23 ],
   alphaCSR[ 208 ][ 24 ],
   alphaCSR[ 208 ][ 25 ],
   alphaCSR[ 208 ][ 26 ],
   alphaCSR[ 208 ][ 27 ],
   alphaCSR[ 208 ][ 28 ],
   alphaCSR[ 208 ][ 29 ],
   alphaCSR[ 208 ][ 30 ],
   alphaCSR[ 208 ][ 31 ],
   alphaCSR[ 208 ][ 32 ],
   alphaCSR[ 208 ][ 33 ],
   alphaCSR[ 208 ][ 34 ],
   alphaCSR[ 208 ][ 35 ],
   alphaCSR[ 208 ][ 36 ],
   alphaCSR[ 208 ][ 37 ],
   alphaCSR[ 208 ][ 38 ],
   alphaCSR[ 208 ][ 39 ],
   alphaCSR[ 208 ][ 40 ],
   alphaCSR[ 208 ][ 41 ],
   alphaCSR[ 208 ][ 42 ],
   alphaCSR[ 208 ][ 43 ],
   alphaCSR[ 208 ][ 44 ],
   alphaCSR[ 208 ][ 45 ],
   alphaCSR[ 208 ][ 46 ],
   alphaCSR[ 208 ][ 47 ],
   alphaCSR[ 208 ][ 48 ],
   alphaCSR[ 208 ][ 49 ],
   alphaCSR[ 208 ][ 50 ],
   alphaCSR[ 208 ][ 51 ],
   alphaCSR[ 208 ][ 52 ],
   alphaCSR[ 208 ][ 53 ],
   alphaCSR[ 208 ][ 54 ],
   alphaCSR[ 208 ][ 55 ],
   alphaCSR[ 208 ][ 56 ],
   alphaCSR[ 208 ][ 57 ],
   alphaCSR[ 208 ][ 58 ],
   alphaCSR[ 208 ][ 59 ],
   alphaCSR[ 208 ][ 60 ],
   alphaCSR[ 208 ][ 61 ],
   alphaCSR[ 208 ][ 62 ],
   alphaCSR[ 208 ][ 63 ],
   alphaCSR[ 208 ][ 64 ],
   alphaCSR[ 208 ][ 65 ],
   alphaCSR[ 208 ][ 66 ],
   alphaCSR[ 208 ][ 67 ],
   alphaCSR[ 208 ][ 68 ],
   alphaCSR[ 208 ][ 69 ],
   alphaCSR[ 208 ][ 70 ],
   alphaCSR[ 208 ][ 71 ],
   alphaCSR[ 208 ][ 72 ],
   alphaCSR[ 208 ][ 73 ],
   alphaCSR[ 208 ][ 74 ],
   alphaCSR[ 208 ][ 75 ],
   alphaCSR[ 208 ][ 76 ],
   alphaCSR[ 208 ][ 77 ],
   alphaCSR[ 208 ][ 78 ],
   alphaCSR[ 208 ][ 79 ],
   alphaCSR[ 208 ][ 80 ],
   alphaCSR[ 208 ][ 81 ],
   alphaCSR[ 208 ][ 82 ],
   alphaCSR[ 208 ][ 83 ],
   alphaCSR[ 208 ][ 84 ],
   alphaCSR[ 208 ][ 85 ],
   alphaCSR[ 208 ][ 86 ],
   alphaCSR[ 208 ][ 87 ],
   alphaCSR[ 208 ][ 88 ],
   alphaCSR[ 208 ][ 89 ],
   alphaCSR[ 208 ][ 90 ],
   alphaCSR[ 208 ][ 91 ],
   alphaCSR[ 208 ][ 92 ],
   alphaCSR[ 208 ][ 93 ],
   alphaCSR[ 208 ][ 94 ],
   alphaCSR[ 208 ][ 95 ],
   alphaCSR[ 208 ][ 96 ],
   alphaCSR[ 208 ][ 97 ],
   alphaCSR[ 208 ][ 98 ],
   alphaCSR[ 208 ][ 99 ],
   alphaCSR[ 208 ][ 100 ],
   alphaCSR[ 208 ][ 101 ],
   alphaCSR[ 208 ][ 102 ],
   alphaCSR[ 208 ][ 103 ],
   alphaCSR[ 208 ][ 104 ],
   alphaCSR[ 208 ][ 105 ],
   alphaCSR[ 208 ][ 106 ],
   alphaCSR[ 208 ][ 107 ],
   alphaCSR[ 208 ][ 108 ],
   alphaCSR[ 208 ][ 109 ],
   alphaCSR[ 208 ][ 110 ],
   alphaCSR[ 208 ][ 111 ],
   alphaCSR[ 208 ][ 112 ],
   alphaCSR[ 208 ][ 113 ],
   alphaCSR[ 208 ][ 114 ],
   alphaCSR[ 208 ][ 115 ],
   alphaCSR[ 208 ][ 116 ],
   alphaCSR[ 208 ][ 117 ],
   alphaCSR[ 208 ][ 118 ],
   alphaCSR[ 208 ][ 119 ],
   alphaCSR[ 208 ][ 120 ],
   alphaCSR[ 208 ][ 121 ],
   alphaCSR[ 208 ][ 122 ],
   alphaCSR[ 208 ][ 123 ],
   alphaCSR[ 208 ][ 124 ],
   alphaCSR[ 208 ][ 125 ],
   alphaCSR[ 208 ][ 126 ],
   alphaCSR[ 208 ][ 127 ],
   alphaCSR[ 208 ][ 128 ],
   alphaCSR[ 208 ][ 129 ],
   alphaCSR[ 208 ][ 130 ],
   alphaCSR[ 208 ][ 131 ],
   alphaCSR[ 208 ][ 132 ],
   alphaCSR[ 208 ][ 133 ],
   alphaCSR[ 208 ][ 134 ],
   alphaCSR[ 208 ][ 135 ],
   alphaCSR[ 208 ][ 136 ],
   alphaCSR[ 208 ][ 137 ],
   alphaCSR[ 208 ][ 138 ],
   alphaCSR[ 208 ][ 139 ],
   alphaCSR[ 208 ][ 140 ],
   alphaCSR[ 208 ][ 141 ],
   alphaCSR[ 208 ][ 142 ],
   alphaCSR[ 208 ][ 143 ],
   alphaCSR[ 208 ][ 144 ],
   alphaCSR[ 208 ][ 145 ],
   alphaCSR[ 208 ][ 146 ],
   alphaCSR[ 208 ][ 147 ],
   alphaCSR[ 208 ][ 148 ],
   alphaCSR[ 208 ][ 149 ],
   alphaCSR[ 208 ][ 150 ],
   alphaCSR[ 208 ][ 151 ],
   alphaCSR[ 208 ][ 152 ],
   alphaCSR[ 208 ][ 153 ],
   alphaCSR[ 208 ][ 154 ],
   alphaCSR[ 208 ][ 155 ],
   alphaCSR[ 208 ][ 156 ],
   alphaCSR[ 208 ][ 157 ],
   alphaCSR[ 208 ][ 158 ],
   alphaCSR[ 208 ][ 159 ],
   alphaCSR[ 208 ][ 160 ],
   alphaCSR[ 208 ][ 161 ],
   alphaCSR[ 208 ][ 162 ],
   alphaCSR[ 208 ][ 163 ],
   alphaCSR[ 208 ][ 164 ],
   alphaCSR[ 208 ][ 165 ],
   alphaCSR[ 208 ][ 166 ],
   alphaCSR[ 208 ][ 167 ],
   alphaCSR[ 208 ][ 168 ],
   alphaCSR[ 208 ][ 169 ],
   alphaCSR[ 208 ][ 170 ],
   alphaCSR[ 208 ][ 171 ],
   alphaCSR[ 208 ][ 172 ],
   alphaCSR[ 208 ][ 173 ],
   alphaCSR[ 208 ][ 174 ],
   alphaCSR[ 208 ][ 175 ],
   alphaCSR[ 208 ][ 176 ],
   alphaCSR[ 208 ][ 177 ],
   alphaCSR[ 208 ][ 178 ],
   alphaCSR[ 208 ][ 179 ],
   alphaCSR[ 208 ][ 180 ],
   alphaCSR[ 208 ][ 181 ],
   alphaCSR[ 208 ][ 182 ],
   alphaCSR[ 208 ][ 183 ],
   alphaCSR[ 208 ][ 184 ],
   alphaCSR[ 208 ][ 185 ],
   alphaCSR[ 208 ][ 186 ],
   alphaCSR[ 208 ][ 187 ],
   alphaCSR[ 208 ][ 188 ],
   alphaCSR[ 208 ][ 189 ],
   alphaCSR[ 208 ][ 190 ],
   alphaCSR[ 208 ][ 191 ],
   alphaCSR[ 208 ][ 192 ],
   alphaCSR[ 208 ][ 193 ],
   alphaCSR[ 208 ][ 194 ],
   alphaCSR[ 208 ][ 195 ],
   alphaCSR[ 208 ][ 196 ],
   alphaCSR[ 208 ][ 197 ],
   alphaCSR[ 208 ][ 198 ],
   alphaCSR[ 208 ][ 199 ],
   alphaCSR[ 208 ][ 200 ],
   alphaCSR[ 208 ][ 201 ],
   alphaCSR[ 208 ][ 202 ],
   alphaCSR[ 208 ][ 203 ],
   alphaCSR[ 208 ][ 204 ],
   alphaCSR[ 208 ][ 205 ],
   alphaCSR[ 208 ][ 206 ],
   alphaCSR[ 208 ][ 207 ],
   alphaCSR[ 208 ][ 208 ],
   alphaCSR[ 208 ][ 209 ],
   alphaCSR[ 208 ][ 210 ],
   alphaCSR[ 208 ][ 211 ],
   alphaCSR[ 208 ][ 212 ],
   alphaCSR[ 208 ][ 213 ],
   alphaCSR[ 208 ][ 214 ],
   alphaCSR[ 208 ][ 215 ],
   alphaCSR[ 208 ][ 216 ],
   alphaCSR[ 208 ][ 217 ],
   alphaCSR[ 208 ][ 218 ],
   alphaCSR[ 208 ][ 219 ],
   alphaCSR[ 208 ][ 220 ],
   alphaCSR[ 208 ][ 221 ],
   alphaCSR[ 208 ][ 222 ],
   alphaCSR[ 208 ][ 223 ],
   alphaCSR[ 208 ][ 224 ],
   alphaCSR[ 208 ][ 225 ],
   alphaCSR[ 208 ][ 226 ],
   alphaCSR[ 208 ][ 227 ],
   alphaCSR[ 208 ][ 228 ],
   alphaCSR[ 208 ][ 229 ],
   alphaCSR[ 208 ][ 230 ],
   alphaCSR[ 208 ][ 231 ],
   alphaCSR[ 208 ][ 232 ],
   alphaCSR[ 208 ][ 233 ],
   alphaCSR[ 208 ][ 234 ],
   alphaCSR[ 208 ][ 235 ],
   alphaCSR[ 208 ][ 236 ],
   alphaCSR[ 208 ][ 237 ],
   alphaCSR[ 208 ][ 238 ],
   alphaCSR[ 208 ][ 239 ],
   alphaCSR[ 208 ][ 240 ],
   alphaCSR[ 208 ][ 241 ],
   alphaCSR[ 208 ][ 242 ],
   alphaCSR[ 208 ][ 243 ],
   alphaCSR[ 208 ][ 244 ],
   alphaCSR[ 208 ][ 245 ],
   alphaCSR[ 208 ][ 246 ],
   alphaCSR[ 208 ][ 247 ],
   alphaCSR[ 208 ][ 248 ],
   alphaCSR[ 208 ][ 249 ],
   alphaCSR[ 208 ][ 250 ],
   alphaCSR[ 208 ][ 251 ],
   alphaCSR[ 208 ][ 252 ],
   alphaCSR[ 208 ][ 253 ],
   alphaCSR[ 208 ][ 254 ],
   alphaCSR[ 208 ][ 255 ],
   alphaCSR[ 208 ][ 256 ],
   alphaCSR[ 208 ][ 257 ],
   alphaCSR[ 208 ][ 258 ],
   alphaCSR[ 208 ][ 259 ],
   alphaCSR[ 208 ][ 260 ],
   alphaCSR[ 208 ][ 261 ],
   alphaCSR[ 208 ][ 262 ],
   alphaCSR[ 208 ][ 263 ],
   alphaCSR[ 208 ][ 264 ],
   alphaCSR[ 208 ][ 265 ],
   alphaCSR[ 208 ][ 266 ],
   alphaCSR[ 208 ][ 267 ],
   alphaCSR[ 208 ][ 268 ],
   alphaCSR[ 208 ][ 269 ],
   alphaCSR[ 208 ][ 270 ],
   alphaCSR[ 208 ][ 271 ],
   alphaCSR[ 208 ][ 272 ],
   alphaCSR[ 208 ][ 273 ],
   alphaCSR[ 208 ][ 274 ],
   alphaCSR[ 208 ][ 275 ],
   alphaCSR[ 208 ][ 276 ],
   alphaCSR[ 208 ][ 277 ],
   alphaCSR[ 208 ][ 278 ],
   alphaCSR[ 208 ][ 279 ],
   alphaCSR[ 208 ][ 280 ],
   alphaCSR[ 208 ][ 281 ],
   alphaCSR[ 208 ][ 282 ],
   alphaCSR[ 208 ][ 283 ],
   alphaCSR[ 208 ][ 284 ],
   alphaCSR[ 208 ][ 285 ],
   alphaCSR[ 208 ][ 286 ],
   alphaCSR[ 208 ][ 287 ],
   alphaCSR[ 208 ][ 288 ],
   alphaCSR[ 208 ][ 289 ],
   alphaCSR[ 208 ][ 290 ],
   alphaCSR[ 208 ][ 291 ],
   alphaCSR[ 208 ][ 292 ],
   alphaCSR[ 208 ][ 293 ],
   alphaCSR[ 208 ][ 294 ],
   alphaCSR[ 208 ][ 295 ],
   alphaCSR[ 208 ][ 296 ],
   alphaCSR[ 208 ][ 297 ],
   alphaCSR[ 208 ][ 298 ],
   alphaCSR[ 208 ][ 299 ],
   alphaCSR[ 208 ][ 300 ],
   alphaCSR[ 208 ][ 301 ],
   alphaCSR[ 208 ][ 302 ],
   alphaCSR[ 208 ][ 303 ],
   alphaCSR[ 208 ][ 304 ],
   alphaCSR[ 208 ][ 305 ],
   alphaCSR[ 208 ][ 306 ],
   alphaCSR[ 208 ][ 307 ],
   alphaCSR[ 208 ][ 308 ],
   alphaCSR[ 208 ][ 309 ],
   alphaCSR[ 208 ][ 310 ],
   alphaCSR[ 208 ][ 311 ],
   alphaCSR[ 208 ][ 312 ],
   alphaCSR[ 208 ][ 313 ],
   alphaCSR[ 208 ][ 314 ],
   alphaCSR[ 208 ][ 315 ],
   alphaCSR[ 208 ][ 316 ],
   alphaCSR[ 208 ][ 317 ],
   alphaCSR[ 208 ][ 318 ],
   alphaCSR[ 208 ][ 319 ],
   alphaCSR[ 208 ][ 320 ],
   alphaCSR[ 208 ][ 321 ],
   alphaCSR[ 208 ][ 322 ],
   alphaCSR[ 208 ][ 323 ],
   alphaCSR[ 208 ][ 324 ],
   alphaCSR[ 208 ][ 325 ],
   alphaCSR[ 208 ][ 326 ],
   alphaCSR[ 208 ][ 327 ],
   alphaCSR[ 208 ][ 328 ],
   alphaCSR[ 208 ][ 329 ],
   alphaCSR[ 208 ][ 330 ],
   alphaCSR[ 208 ][ 331 ],
   alphaCSR[ 208 ][ 332 ],
   alphaCSR[ 208 ][ 333 ],
   alphaCSR[ 208 ][ 334 ],
   alphaCSR[ 208 ][ 335 ],
   alphaCSR[ 208 ][ 336 ],
   alphaCSR[ 208 ][ 337 ],
   alphaCSR[ 208 ][ 338 ],
   alphaCSR[ 208 ][ 339 ],
   alphaCSR[ 208 ][ 340 ],
   alphaCSR[ 208 ][ 341 ],
   alphaCSR[ 208 ][ 342 ],
   alphaCSR[ 208 ][ 343 ],
   alphaCSR[ 208 ][ 344 ],
   alphaCSR[ 208 ][ 345 ],
   alphaCSR[ 208 ][ 346 ],
   alphaCSR[ 208 ][ 347 ],
   alphaCSR[ 208 ][ 348 ],
   alphaCSR[ 208 ][ 349 ],
   alphaCSR[ 208 ][ 350 ],
   alphaCSR[ 208 ][ 351 ],
   alphaCSR[ 208 ][ 352 ],
   alphaCSR[ 208 ][ 353 ],
   alphaCSR[ 208 ][ 354 ],
   alphaCSR[ 208 ][ 355 ],
   alphaCSR[ 208 ][ 356 ],
   alphaCSR[ 208 ][ 357 ],
   alphaCSR[ 208 ][ 358 ],
   alphaCSR[ 208 ][ 359 ],
   alphaCSR[ 208 ][ 360 ],
   alphaCSR[ 208 ][ 361 ],
   alphaCSR[ 208 ][ 362 ],
   alphaCSR[ 208 ][ 363 ],
   alphaCSR[ 208 ][ 364 ],
   alphaCSR[ 208 ][ 365 ],
   alphaCSR[ 208 ][ 366 ],
   alphaCSR[ 208 ][ 367 ],
   alphaCSR[ 208 ][ 368 ],
   alphaCSR[ 208 ][ 369 ],
   alphaCSR[ 208 ][ 370 ],
   alphaCSR[ 208 ][ 371 ],
   alphaCSR[ 208 ][ 372 ],
   alphaCSR[ 208 ][ 373 ],
   alphaCSR[ 208 ][ 374 ],
   alphaCSR[ 208 ][ 375 ],
   alphaCSR[ 208 ][ 376 ],
   alphaCSR[ 208 ][ 377 ],
   alphaCSR[ 208 ][ 378 ],
   alphaCSR[ 208 ][ 379 ],
   alphaCSR[ 208 ][ 380 ],
   alphaCSR[ 208 ][ 381 ],
   alphaCSR[ 208 ][ 382 ],
   alphaCSR[ 208 ][ 383 ],
   alphaCSR[ 209 ][ 0 ],
   alphaCSR[ 209 ][ 1 ],
   alphaCSR[ 209 ][ 2 ],
   alphaCSR[ 209 ][ 3 ],
   alphaCSR[ 209 ][ 4 ],
   alphaCSR[ 209 ][ 5 ],
   alphaCSR[ 209 ][ 6 ],
   alphaCSR[ 209 ][ 7 ],
   alphaCSR[ 209 ][ 8 ],
   alphaCSR[ 209 ][ 9 ],
   alphaCSR[ 209 ][ 10 ],
   alphaCSR[ 209 ][ 11 ],
   alphaCSR[ 209 ][ 12 ],
   alphaCSR[ 209 ][ 13 ],
   alphaCSR[ 209 ][ 14 ],
   alphaCSR[ 209 ][ 15 ],
   alphaCSR[ 209 ][ 16 ],
   alphaCSR[ 209 ][ 17 ],
   alphaCSR[ 209 ][ 18 ],
   alphaCSR[ 209 ][ 19 ],
   alphaCSR[ 209 ][ 20 ],
   alphaCSR[ 209 ][ 21 ],
   alphaCSR[ 209 ][ 22 ],
   alphaCSR[ 209 ][ 23 ],
   alphaCSR[ 209 ][ 24 ],
   alphaCSR[ 209 ][ 25 ],
   alphaCSR[ 209 ][ 26 ],
   alphaCSR[ 209 ][ 27 ],
   alphaCSR[ 209 ][ 28 ],
   alphaCSR[ 209 ][ 29 ],
   alphaCSR[ 209 ][ 30 ],
   alphaCSR[ 209 ][ 31 ],
   alphaCSR[ 209 ][ 32 ],
   alphaCSR[ 209 ][ 33 ],
   alphaCSR[ 209 ][ 34 ],
   alphaCSR[ 209 ][ 35 ],
   alphaCSR[ 209 ][ 36 ],
   alphaCSR[ 209 ][ 37 ],
   alphaCSR[ 209 ][ 38 ],
   alphaCSR[ 209 ][ 39 ],
   alphaCSR[ 209 ][ 40 ],
   alphaCSR[ 209 ][ 41 ],
   alphaCSR[ 209 ][ 42 ],
   alphaCSR[ 209 ][ 43 ],
   alphaCSR[ 209 ][ 44 ],
   alphaCSR[ 209 ][ 45 ],
   alphaCSR[ 209 ][ 46 ],
   alphaCSR[ 209 ][ 47 ],
   alphaCSR[ 209 ][ 48 ],
   alphaCSR[ 209 ][ 49 ],
   alphaCSR[ 209 ][ 50 ],
   alphaCSR[ 209 ][ 51 ],
   alphaCSR[ 209 ][ 52 ],
   alphaCSR[ 209 ][ 53 ],
   alphaCSR[ 209 ][ 54 ],
   alphaCSR[ 209 ][ 55 ],
   alphaCSR[ 209 ][ 56 ],
   alphaCSR[ 209 ][ 57 ],
   alphaCSR[ 209 ][ 58 ],
   alphaCSR[ 209 ][ 59 ],
   alphaCSR[ 209 ][ 60 ],
   alphaCSR[ 209 ][ 61 ],
   alphaCSR[ 209 ][ 62 ],
   alphaCSR[ 209 ][ 63 ],
   alphaCSR[ 209 ][ 64 ],
   alphaCSR[ 209 ][ 65 ],
   alphaCSR[ 209 ][ 66 ],
   alphaCSR[ 209 ][ 67 ],
   alphaCSR[ 209 ][ 68 ],
   alphaCSR[ 209 ][ 69 ],
   alphaCSR[ 209 ][ 70 ],
   alphaCSR[ 209 ][ 71 ],
   alphaCSR[ 209 ][ 72 ],
   alphaCSR[ 209 ][ 73 ],
   alphaCSR[ 209 ][ 74 ],
   alphaCSR[ 209 ][ 75 ],
   alphaCSR[ 209 ][ 76 ],
   alphaCSR[ 209 ][ 77 ],
   alphaCSR[ 209 ][ 78 ],
   alphaCSR[ 209 ][ 79 ],
   alphaCSR[ 209 ][ 80 ],
   alphaCSR[ 209 ][ 81 ],
   alphaCSR[ 209 ][ 82 ],
   alphaCSR[ 209 ][ 83 ],
   alphaCSR[ 209 ][ 84 ],
   alphaCSR[ 209 ][ 85 ],
   alphaCSR[ 209 ][ 86 ],
   alphaCSR[ 209 ][ 87 ],
   alphaCSR[ 209 ][ 88 ],
   alphaCSR[ 209 ][ 89 ],
   alphaCSR[ 209 ][ 90 ],
   alphaCSR[ 209 ][ 91 ],
   alphaCSR[ 209 ][ 92 ],
   alphaCSR[ 209 ][ 93 ],
   alphaCSR[ 209 ][ 94 ],
   alphaCSR[ 209 ][ 95 ],
   alphaCSR[ 209 ][ 96 ],
   alphaCSR[ 209 ][ 97 ],
   alphaCSR[ 209 ][ 98 ],
   alphaCSR[ 209 ][ 99 ],
   alphaCSR[ 209 ][ 100 ],
   alphaCSR[ 209 ][ 101 ],
   alphaCSR[ 209 ][ 102 ],
   alphaCSR[ 209 ][ 103 ],
   alphaCSR[ 209 ][ 104 ],
   alphaCSR[ 209 ][ 105 ],
   alphaCSR[ 209 ][ 106 ],
   alphaCSR[ 209 ][ 107 ],
   alphaCSR[ 209 ][ 108 ],
   alphaCSR[ 209 ][ 109 ],
   alphaCSR[ 209 ][ 110 ],
   alphaCSR[ 209 ][ 111 ],
   alphaCSR[ 209 ][ 112 ],
   alphaCSR[ 209 ][ 113 ],
   alphaCSR[ 209 ][ 114 ],
   alphaCSR[ 209 ][ 115 ],
   alphaCSR[ 209 ][ 116 ],
   alphaCSR[ 209 ][ 117 ],
   alphaCSR[ 209 ][ 118 ],
   alphaCSR[ 209 ][ 119 ],
   alphaCSR[ 209 ][ 120 ],
   alphaCSR[ 209 ][ 121 ],
   alphaCSR[ 209 ][ 122 ],
   alphaCSR[ 209 ][ 123 ],
   alphaCSR[ 209 ][ 124 ],
   alphaCSR[ 209 ][ 125 ],
   alphaCSR[ 209 ][ 126 ],
   alphaCSR[ 209 ][ 127 ],
   alphaCSR[ 209 ][ 128 ],
   alphaCSR[ 209 ][ 129 ],
   alphaCSR[ 209 ][ 130 ],
   alphaCSR[ 209 ][ 131 ],
   alphaCSR[ 209 ][ 132 ],
   alphaCSR[ 209 ][ 133 ],
   alphaCSR[ 209 ][ 134 ],
   alphaCSR[ 209 ][ 135 ],
   alphaCSR[ 209 ][ 136 ],
   alphaCSR[ 209 ][ 137 ],
   alphaCSR[ 209 ][ 138 ],
   alphaCSR[ 209 ][ 139 ],
   alphaCSR[ 209 ][ 140 ],
   alphaCSR[ 209 ][ 141 ],
   alphaCSR[ 209 ][ 142 ],
   alphaCSR[ 209 ][ 143 ],
   alphaCSR[ 209 ][ 144 ],
   alphaCSR[ 209 ][ 145 ],
   alphaCSR[ 209 ][ 146 ],
   alphaCSR[ 209 ][ 147 ],
   alphaCSR[ 209 ][ 148 ],
   alphaCSR[ 209 ][ 149 ],
   alphaCSR[ 209 ][ 150 ],
   alphaCSR[ 209 ][ 151 ],
   alphaCSR[ 209 ][ 152 ],
   alphaCSR[ 209 ][ 153 ],
   alphaCSR[ 209 ][ 154 ],
   alphaCSR[ 209 ][ 155 ],
   alphaCSR[ 209 ][ 156 ],
   alphaCSR[ 209 ][ 157 ],
   alphaCSR[ 209 ][ 158 ],
   alphaCSR[ 209 ][ 159 ],
   alphaCSR[ 209 ][ 160 ],
   alphaCSR[ 209 ][ 161 ],
   alphaCSR[ 209 ][ 162 ],
   alphaCSR[ 209 ][ 163 ],
   alphaCSR[ 209 ][ 164 ],
   alphaCSR[ 209 ][ 165 ],
   alphaCSR[ 209 ][ 166 ],
   alphaCSR[ 209 ][ 167 ],
   alphaCSR[ 209 ][ 168 ],
   alphaCSR[ 209 ][ 169 ],
   alphaCSR[ 209 ][ 170 ],
   alphaCSR[ 209 ][ 171 ],
   alphaCSR[ 209 ][ 172 ],
   alphaCSR[ 209 ][ 173 ],
   alphaCSR[ 209 ][ 174 ],
   alphaCSR[ 209 ][ 175 ],
   alphaCSR[ 209 ][ 176 ],
   alphaCSR[ 209 ][ 177 ],
   alphaCSR[ 209 ][ 178 ],
   alphaCSR[ 209 ][ 179 ],
   alphaCSR[ 209 ][ 180 ],
   alphaCSR[ 209 ][ 181 ],
   alphaCSR[ 209 ][ 182 ],
   alphaCSR[ 209 ][ 183 ],
   alphaCSR[ 209 ][ 184 ],
   alphaCSR[ 209 ][ 185 ],
   alphaCSR[ 209 ][ 186 ],
   alphaCSR[ 209 ][ 187 ],
   alphaCSR[ 209 ][ 188 ],
   alphaCSR[ 209 ][ 189 ],
   alphaCSR[ 209 ][ 190 ],
   alphaCSR[ 209 ][ 191 ],
   alphaCSR[ 209 ][ 192 ],
   alphaCSR[ 209 ][ 193 ],
   alphaCSR[ 209 ][ 194 ],
   alphaCSR[ 209 ][ 195 ],
   alphaCSR[ 209 ][ 196 ],
   alphaCSR[ 209 ][ 197 ],
   alphaCSR[ 209 ][ 198 ],
   alphaCSR[ 209 ][ 199 ],
   alphaCSR[ 209 ][ 200 ],
   alphaCSR[ 209 ][ 201 ],
   alphaCSR[ 209 ][ 202 ],
   alphaCSR[ 209 ][ 203 ],
   alphaCSR[ 209 ][ 204 ],
   alphaCSR[ 209 ][ 205 ],
   alphaCSR[ 209 ][ 206 ],
   alphaCSR[ 209 ][ 207 ],
   alphaCSR[ 209 ][ 208 ],
   alphaCSR[ 209 ][ 209 ],
   alphaCSR[ 209 ][ 210 ],
   alphaCSR[ 209 ][ 211 ],
   alphaCSR[ 209 ][ 212 ],
   alphaCSR[ 209 ][ 213 ],
   alphaCSR[ 209 ][ 214 ],
   alphaCSR[ 209 ][ 215 ],
   alphaCSR[ 209 ][ 216 ],
   alphaCSR[ 209 ][ 217 ],
   alphaCSR[ 209 ][ 218 ],
   alphaCSR[ 209 ][ 219 ],
   alphaCSR[ 209 ][ 220 ],
   alphaCSR[ 209 ][ 221 ],
   alphaCSR[ 209 ][ 222 ],
   alphaCSR[ 209 ][ 223 ],
   alphaCSR[ 209 ][ 224 ],
   alphaCSR[ 209 ][ 225 ],
   alphaCSR[ 209 ][ 226 ],
   alphaCSR[ 209 ][ 227 ],
   alphaCSR[ 209 ][ 228 ],
   alphaCSR[ 209 ][ 229 ],
   alphaCSR[ 209 ][ 230 ],
   alphaCSR[ 209 ][ 231 ],
   alphaCSR[ 209 ][ 232 ],
   alphaCSR[ 209 ][ 233 ],
   alphaCSR[ 209 ][ 234 ],
   alphaCSR[ 209 ][ 235 ],
   alphaCSR[ 209 ][ 236 ],
   alphaCSR[ 209 ][ 237 ],
   alphaCSR[ 209 ][ 238 ],
   alphaCSR[ 209 ][ 239 ],
   alphaCSR[ 209 ][ 240 ],
   alphaCSR[ 209 ][ 241 ],
   alphaCSR[ 209 ][ 242 ],
   alphaCSR[ 209 ][ 243 ],
   alphaCSR[ 209 ][ 244 ],
   alphaCSR[ 209 ][ 245 ],
   alphaCSR[ 209 ][ 246 ],
   alphaCSR[ 209 ][ 247 ],
   alphaCSR[ 209 ][ 248 ],
   alphaCSR[ 209 ][ 249 ],
   alphaCSR[ 209 ][ 250 ],
   alphaCSR[ 209 ][ 251 ],
   alphaCSR[ 209 ][ 252 ],
   alphaCSR[ 209 ][ 253 ],
   alphaCSR[ 209 ][ 254 ],
   alphaCSR[ 209 ][ 255 ],
   alphaCSR[ 209 ][ 256 ],
   alphaCSR[ 209 ][ 257 ],
   alphaCSR[ 209 ][ 258 ],
   alphaCSR[ 209 ][ 259 ],
   alphaCSR[ 209 ][ 260 ],
   alphaCSR[ 209 ][ 261 ],
   alphaCSR[ 209 ][ 262 ],
   alphaCSR[ 209 ][ 263 ],
   alphaCSR[ 209 ][ 264 ],
   alphaCSR[ 209 ][ 265 ],
   alphaCSR[ 209 ][ 266 ],
   alphaCSR[ 209 ][ 267 ],
   alphaCSR[ 209 ][ 268 ],
   alphaCSR[ 209 ][ 269 ],
   alphaCSR[ 209 ][ 270 ],
   alphaCSR[ 209 ][ 271 ],
   alphaCSR[ 209 ][ 272 ],
   alphaCSR[ 209 ][ 273 ],
   alphaCSR[ 209 ][ 274 ],
   alphaCSR[ 209 ][ 275 ],
   alphaCSR[ 209 ][ 276 ],
   alphaCSR[ 209 ][ 277 ],
   alphaCSR[ 209 ][ 278 ],
   alphaCSR[ 209 ][ 279 ],
   alphaCSR[ 209 ][ 280 ],
   alphaCSR[ 209 ][ 281 ],
   alphaCSR[ 209 ][ 282 ],
   alphaCSR[ 209 ][ 283 ],
   alphaCSR[ 209 ][ 284 ],
   alphaCSR[ 209 ][ 285 ],
   alphaCSR[ 209 ][ 286 ],
   alphaCSR[ 209 ][ 287 ],
   alphaCSR[ 209 ][ 288 ],
   alphaCSR[ 209 ][ 289 ],
   alphaCSR[ 209 ][ 290 ],
   alphaCSR[ 209 ][ 291 ],
   alphaCSR[ 209 ][ 292 ],
   alphaCSR[ 209 ][ 293 ],
   alphaCSR[ 209 ][ 294 ],
   alphaCSR[ 209 ][ 295 ],
   alphaCSR[ 209 ][ 296 ],
   alphaCSR[ 209 ][ 297 ],
   alphaCSR[ 209 ][ 298 ],
   alphaCSR[ 209 ][ 299 ],
   alphaCSR[ 209 ][ 300 ],
   alphaCSR[ 209 ][ 301 ],
   alphaCSR[ 209 ][ 302 ],
   alphaCSR[ 209 ][ 303 ],
   alphaCSR[ 209 ][ 304 ],
   alphaCSR[ 209 ][ 305 ],
   alphaCSR[ 209 ][ 306 ],
   alphaCSR[ 209 ][ 307 ],
   alphaCSR[ 209 ][ 308 ],
   alphaCSR[ 209 ][ 309 ],
   alphaCSR[ 209 ][ 310 ],
   alphaCSR[ 209 ][ 311 ],
   alphaCSR[ 209 ][ 312 ],
   alphaCSR[ 209 ][ 313 ],
   alphaCSR[ 209 ][ 314 ],
   alphaCSR[ 209 ][ 315 ],
   alphaCSR[ 209 ][ 316 ],
   alphaCSR[ 209 ][ 317 ],
   alphaCSR[ 209 ][ 318 ],
   alphaCSR[ 209 ][ 319 ],
   alphaCSR[ 209 ][ 320 ],
   alphaCSR[ 209 ][ 321 ],
   alphaCSR[ 209 ][ 322 ],
   alphaCSR[ 209 ][ 323 ],
   alphaCSR[ 209 ][ 324 ],
   alphaCSR[ 209 ][ 325 ],
   alphaCSR[ 209 ][ 326 ],
   alphaCSR[ 209 ][ 327 ],
   alphaCSR[ 209 ][ 328 ],
   alphaCSR[ 209 ][ 329 ],
   alphaCSR[ 209 ][ 330 ],
   alphaCSR[ 209 ][ 331 ],
   alphaCSR[ 209 ][ 332 ],
   alphaCSR[ 209 ][ 333 ],
   alphaCSR[ 209 ][ 334 ],
   alphaCSR[ 209 ][ 335 ],
   alphaCSR[ 209 ][ 336 ],
   alphaCSR[ 209 ][ 337 ],
   alphaCSR[ 209 ][ 338 ],
   alphaCSR[ 209 ][ 339 ],
   alphaCSR[ 209 ][ 340 ],
   alphaCSR[ 209 ][ 341 ],
   alphaCSR[ 209 ][ 342 ],
   alphaCSR[ 209 ][ 343 ],
   alphaCSR[ 209 ][ 344 ],
   alphaCSR[ 209 ][ 345 ],
   alphaCSR[ 209 ][ 346 ],
   alphaCSR[ 209 ][ 347 ],
   alphaCSR[ 209 ][ 348 ],
   alphaCSR[ 209 ][ 349 ],
   alphaCSR[ 209 ][ 350 ],
   alphaCSR[ 209 ][ 351 ],
   alphaCSR[ 209 ][ 352 ],
   alphaCSR[ 209 ][ 353 ],
   alphaCSR[ 209 ][ 354 ],
   alphaCSR[ 209 ][ 355 ],
   alphaCSR[ 209 ][ 356 ],
   alphaCSR[ 209 ][ 357 ],
   alphaCSR[ 209 ][ 358 ],
   alphaCSR[ 209 ][ 359 ],
   alphaCSR[ 209 ][ 360 ],
   alphaCSR[ 209 ][ 361 ],
   alphaCSR[ 209 ][ 362 ],
   alphaCSR[ 209 ][ 363 ],
   alphaCSR[ 209 ][ 364 ],
   alphaCSR[ 209 ][ 365 ],
   alphaCSR[ 209 ][ 366 ],
   alphaCSR[ 209 ][ 367 ],
   alphaCSR[ 209 ][ 368 ],
   alphaCSR[ 209 ][ 369 ],
   alphaCSR[ 209 ][ 370 ],
   alphaCSR[ 209 ][ 371 ],
   alphaCSR[ 209 ][ 372 ],
   alphaCSR[ 209 ][ 373 ],
   alphaCSR[ 209 ][ 374 ],
   alphaCSR[ 209 ][ 375 ],
   alphaCSR[ 209 ][ 376 ],
   alphaCSR[ 209 ][ 377 ],
   alphaCSR[ 209 ][ 378 ],
   alphaCSR[ 209 ][ 379 ],
   alphaCSR[ 209 ][ 380 ],
   alphaCSR[ 209 ][ 381 ],
   alphaCSR[ 209 ][ 382 ],
   alphaCSR[ 209 ][ 383 ],
   alphaCSR[ 210 ][ 0 ],
   alphaCSR[ 210 ][ 1 ],
   alphaCSR[ 210 ][ 2 ],
   alphaCSR[ 210 ][ 3 ],
   alphaCSR[ 210 ][ 4 ],
   alphaCSR[ 210 ][ 5 ],
   alphaCSR[ 210 ][ 6 ],
   alphaCSR[ 210 ][ 7 ],
   alphaCSR[ 210 ][ 8 ],
   alphaCSR[ 210 ][ 9 ],
   alphaCSR[ 210 ][ 10 ],
   alphaCSR[ 210 ][ 11 ],
   alphaCSR[ 210 ][ 12 ],
   alphaCSR[ 210 ][ 13 ],
   alphaCSR[ 210 ][ 14 ],
   alphaCSR[ 210 ][ 15 ],
   alphaCSR[ 210 ][ 16 ],
   alphaCSR[ 210 ][ 17 ],
   alphaCSR[ 210 ][ 18 ],
   alphaCSR[ 210 ][ 19 ],
   alphaCSR[ 210 ][ 20 ],
   alphaCSR[ 210 ][ 21 ],
   alphaCSR[ 210 ][ 22 ],
   alphaCSR[ 210 ][ 23 ],
   alphaCSR[ 210 ][ 24 ],
   alphaCSR[ 210 ][ 25 ],
   alphaCSR[ 210 ][ 26 ],
   alphaCSR[ 210 ][ 27 ],
   alphaCSR[ 210 ][ 28 ],
   alphaCSR[ 210 ][ 29 ],
   alphaCSR[ 210 ][ 30 ],
   alphaCSR[ 210 ][ 31 ],
   alphaCSR[ 210 ][ 32 ],
   alphaCSR[ 210 ][ 33 ],
   alphaCSR[ 210 ][ 34 ],
   alphaCSR[ 210 ][ 35 ],
   alphaCSR[ 210 ][ 36 ],
   alphaCSR[ 210 ][ 37 ],
   alphaCSR[ 210 ][ 38 ],
   alphaCSR[ 210 ][ 39 ],
   alphaCSR[ 210 ][ 40 ],
   alphaCSR[ 210 ][ 41 ],
   alphaCSR[ 210 ][ 42 ],
   alphaCSR[ 210 ][ 43 ],
   alphaCSR[ 210 ][ 44 ],
   alphaCSR[ 210 ][ 45 ],
   alphaCSR[ 210 ][ 46 ],
   alphaCSR[ 210 ][ 47 ],
   alphaCSR[ 210 ][ 48 ],
   alphaCSR[ 210 ][ 49 ],
   alphaCSR[ 210 ][ 50 ],
   alphaCSR[ 210 ][ 51 ],
   alphaCSR[ 210 ][ 52 ],
   alphaCSR[ 210 ][ 53 ],
   alphaCSR[ 210 ][ 54 ],
   alphaCSR[ 210 ][ 55 ],
   alphaCSR[ 210 ][ 56 ],
   alphaCSR[ 210 ][ 57 ],
   alphaCSR[ 210 ][ 58 ],
   alphaCSR[ 210 ][ 59 ],
   alphaCSR[ 210 ][ 60 ],
   alphaCSR[ 210 ][ 61 ],
   alphaCSR[ 210 ][ 62 ],
   alphaCSR[ 210 ][ 63 ],
   alphaCSR[ 210 ][ 64 ],
   alphaCSR[ 210 ][ 65 ],
   alphaCSR[ 210 ][ 66 ],
   alphaCSR[ 210 ][ 67 ],
   alphaCSR[ 210 ][ 68 ],
   alphaCSR[ 210 ][ 69 ],
   alphaCSR[ 210 ][ 70 ],
   alphaCSR[ 210 ][ 71 ],
   alphaCSR[ 210 ][ 72 ],
   alphaCSR[ 210 ][ 73 ],
   alphaCSR[ 210 ][ 74 ],
   alphaCSR[ 210 ][ 75 ],
   alphaCSR[ 210 ][ 76 ],
   alphaCSR[ 210 ][ 77 ],
   alphaCSR[ 210 ][ 78 ],
   alphaCSR[ 210 ][ 79 ],
   alphaCSR[ 210 ][ 80 ],
   alphaCSR[ 210 ][ 81 ],
   alphaCSR[ 210 ][ 82 ],
   alphaCSR[ 210 ][ 83 ],
   alphaCSR[ 210 ][ 84 ],
   alphaCSR[ 210 ][ 85 ],
   alphaCSR[ 210 ][ 86 ],
   alphaCSR[ 210 ][ 87 ],
   alphaCSR[ 210 ][ 88 ],
   alphaCSR[ 210 ][ 89 ],
   alphaCSR[ 210 ][ 90 ],
   alphaCSR[ 210 ][ 91 ],
   alphaCSR[ 210 ][ 92 ],
   alphaCSR[ 210 ][ 93 ],
   alphaCSR[ 210 ][ 94 ],
   alphaCSR[ 210 ][ 95 ],
   alphaCSR[ 210 ][ 96 ],
   alphaCSR[ 210 ][ 97 ],
   alphaCSR[ 210 ][ 98 ],
   alphaCSR[ 210 ][ 99 ],
   alphaCSR[ 210 ][ 100 ],
   alphaCSR[ 210 ][ 101 ],
   alphaCSR[ 210 ][ 102 ],
   alphaCSR[ 210 ][ 103 ],
   alphaCSR[ 210 ][ 104 ],
   alphaCSR[ 210 ][ 105 ],
   alphaCSR[ 210 ][ 106 ],
   alphaCSR[ 210 ][ 107 ],
   alphaCSR[ 210 ][ 108 ],
   alphaCSR[ 210 ][ 109 ],
   alphaCSR[ 210 ][ 110 ],
   alphaCSR[ 210 ][ 111 ],
   alphaCSR[ 210 ][ 112 ],
   alphaCSR[ 210 ][ 113 ],
   alphaCSR[ 210 ][ 114 ],
   alphaCSR[ 210 ][ 115 ],
   alphaCSR[ 210 ][ 116 ],
   alphaCSR[ 210 ][ 117 ],
   alphaCSR[ 210 ][ 118 ],
   alphaCSR[ 210 ][ 119 ],
   alphaCSR[ 210 ][ 120 ],
   alphaCSR[ 210 ][ 121 ],
   alphaCSR[ 210 ][ 122 ],
   alphaCSR[ 210 ][ 123 ],
   alphaCSR[ 210 ][ 124 ],
   alphaCSR[ 210 ][ 125 ],
   alphaCSR[ 210 ][ 126 ],
   alphaCSR[ 210 ][ 127 ],
   alphaCSR[ 210 ][ 128 ],
   alphaCSR[ 210 ][ 129 ],
   alphaCSR[ 210 ][ 130 ],
   alphaCSR[ 210 ][ 131 ],
   alphaCSR[ 210 ][ 132 ],
   alphaCSR[ 210 ][ 133 ],
   alphaCSR[ 210 ][ 134 ],
   alphaCSR[ 210 ][ 135 ],
   alphaCSR[ 210 ][ 136 ],
   alphaCSR[ 210 ][ 137 ],
   alphaCSR[ 210 ][ 138 ],
   alphaCSR[ 210 ][ 139 ],
   alphaCSR[ 210 ][ 140 ],
   alphaCSR[ 210 ][ 141 ],
   alphaCSR[ 210 ][ 142 ],
   alphaCSR[ 210 ][ 143 ],
   alphaCSR[ 210 ][ 144 ],
   alphaCSR[ 210 ][ 145 ],
   alphaCSR[ 210 ][ 146 ],
   alphaCSR[ 210 ][ 147 ],
   alphaCSR[ 210 ][ 148 ],
   alphaCSR[ 210 ][ 149 ],
   alphaCSR[ 210 ][ 150 ],
   alphaCSR[ 210 ][ 151 ],
   alphaCSR[ 210 ][ 152 ],
   alphaCSR[ 210 ][ 153 ],
   alphaCSR[ 210 ][ 154 ],
   alphaCSR[ 210 ][ 155 ],
   alphaCSR[ 210 ][ 156 ],
   alphaCSR[ 210 ][ 157 ],
   alphaCSR[ 210 ][ 158 ],
   alphaCSR[ 210 ][ 159 ],
   alphaCSR[ 210 ][ 160 ],
   alphaCSR[ 210 ][ 161 ],
   alphaCSR[ 210 ][ 162 ],
   alphaCSR[ 210 ][ 163 ],
   alphaCSR[ 210 ][ 164 ],
   alphaCSR[ 210 ][ 165 ],
   alphaCSR[ 210 ][ 166 ],
   alphaCSR[ 210 ][ 167 ],
   alphaCSR[ 210 ][ 168 ],
   alphaCSR[ 210 ][ 169 ],
   alphaCSR[ 210 ][ 170 ],
   alphaCSR[ 210 ][ 171 ],
   alphaCSR[ 210 ][ 172 ],
   alphaCSR[ 210 ][ 173 ],
   alphaCSR[ 210 ][ 174 ],
   alphaCSR[ 210 ][ 175 ],
   alphaCSR[ 210 ][ 176 ],
   alphaCSR[ 210 ][ 177 ],
   alphaCSR[ 210 ][ 178 ],
   alphaCSR[ 210 ][ 179 ],
   alphaCSR[ 210 ][ 180 ],
   alphaCSR[ 210 ][ 181 ],
   alphaCSR[ 210 ][ 182 ],
   alphaCSR[ 210 ][ 183 ],
   alphaCSR[ 210 ][ 184 ],
   alphaCSR[ 210 ][ 185 ],
   alphaCSR[ 210 ][ 186 ],
   alphaCSR[ 210 ][ 187 ],
   alphaCSR[ 210 ][ 188 ],
   alphaCSR[ 210 ][ 189 ],
   alphaCSR[ 210 ][ 190 ],
   alphaCSR[ 210 ][ 191 ],
   alphaCSR[ 210 ][ 192 ],
   alphaCSR[ 210 ][ 193 ],
   alphaCSR[ 210 ][ 194 ],
   alphaCSR[ 210 ][ 195 ],
   alphaCSR[ 210 ][ 196 ],
   alphaCSR[ 210 ][ 197 ],
   alphaCSR[ 210 ][ 198 ],
   alphaCSR[ 210 ][ 199 ],
   alphaCSR[ 210 ][ 200 ],
   alphaCSR[ 210 ][ 201 ],
   alphaCSR[ 210 ][ 202 ],
   alphaCSR[ 210 ][ 203 ],
   alphaCSR[ 210 ][ 204 ],
   alphaCSR[ 210 ][ 205 ],
   alphaCSR[ 210 ][ 206 ],
   alphaCSR[ 210 ][ 207 ],
   alphaCSR[ 210 ][ 208 ],
   alphaCSR[ 210 ][ 209 ],
   alphaCSR[ 210 ][ 210 ],
   alphaCSR[ 210 ][ 211 ],
   alphaCSR[ 210 ][ 212 ],
   alphaCSR[ 210 ][ 213 ],
   alphaCSR[ 210 ][ 214 ],
   alphaCSR[ 210 ][ 215 ],
   alphaCSR[ 210 ][ 216 ],
   alphaCSR[ 210 ][ 217 ],
   alphaCSR[ 210 ][ 218 ],
   alphaCSR[ 210 ][ 219 ],
   alphaCSR[ 210 ][ 220 ],
   alphaCSR[ 210 ][ 221 ],
   alphaCSR[ 210 ][ 222 ],
   alphaCSR[ 210 ][ 223 ],
   alphaCSR[ 210 ][ 224 ],
   alphaCSR[ 210 ][ 225 ],
   alphaCSR[ 210 ][ 226 ],
   alphaCSR[ 210 ][ 227 ],
   alphaCSR[ 210 ][ 228 ],
   alphaCSR[ 210 ][ 229 ],
   alphaCSR[ 210 ][ 230 ],
   alphaCSR[ 210 ][ 231 ],
   alphaCSR[ 210 ][ 232 ],
   alphaCSR[ 210 ][ 233 ],
   alphaCSR[ 210 ][ 234 ],
   alphaCSR[ 210 ][ 235 ],
   alphaCSR[ 210 ][ 236 ],
   alphaCSR[ 210 ][ 237 ],
   alphaCSR[ 210 ][ 238 ],
   alphaCSR[ 210 ][ 239 ],
   alphaCSR[ 210 ][ 240 ],
   alphaCSR[ 210 ][ 241 ],
   alphaCSR[ 210 ][ 242 ],
   alphaCSR[ 210 ][ 243 ],
   alphaCSR[ 210 ][ 244 ],
   alphaCSR[ 210 ][ 245 ],
   alphaCSR[ 210 ][ 246 ],
   alphaCSR[ 210 ][ 247 ],
   alphaCSR[ 210 ][ 248 ],
   alphaCSR[ 210 ][ 249 ],
   alphaCSR[ 210 ][ 250 ],
   alphaCSR[ 210 ][ 251 ],
   alphaCSR[ 210 ][ 252 ],
   alphaCSR[ 210 ][ 253 ],
   alphaCSR[ 210 ][ 254 ],
   alphaCSR[ 210 ][ 255 ],
   alphaCSR[ 210 ][ 256 ],
   alphaCSR[ 210 ][ 257 ],
   alphaCSR[ 210 ][ 258 ],
   alphaCSR[ 210 ][ 259 ],
   alphaCSR[ 210 ][ 260 ],
   alphaCSR[ 210 ][ 261 ],
   alphaCSR[ 210 ][ 262 ],
   alphaCSR[ 210 ][ 263 ],
   alphaCSR[ 210 ][ 264 ],
   alphaCSR[ 210 ][ 265 ],
   alphaCSR[ 210 ][ 266 ],
   alphaCSR[ 210 ][ 267 ],
   alphaCSR[ 210 ][ 268 ],
   alphaCSR[ 210 ][ 269 ],
   alphaCSR[ 210 ][ 270 ],
   alphaCSR[ 210 ][ 271 ],
   alphaCSR[ 210 ][ 272 ],
   alphaCSR[ 210 ][ 273 ],
   alphaCSR[ 210 ][ 274 ],
   alphaCSR[ 210 ][ 275 ],
   alphaCSR[ 210 ][ 276 ],
   alphaCSR[ 210 ][ 277 ],
   alphaCSR[ 210 ][ 278 ],
   alphaCSR[ 210 ][ 279 ],
   alphaCSR[ 210 ][ 280 ],
   alphaCSR[ 210 ][ 281 ],
   alphaCSR[ 210 ][ 282 ],
   alphaCSR[ 210 ][ 283 ],
   alphaCSR[ 210 ][ 284 ],
   alphaCSR[ 210 ][ 285 ],
   alphaCSR[ 210 ][ 286 ],
   alphaCSR[ 210 ][ 287 ],
   alphaCSR[ 210 ][ 288 ],
   alphaCSR[ 210 ][ 289 ],
   alphaCSR[ 210 ][ 290 ],
   alphaCSR[ 210 ][ 291 ],
   alphaCSR[ 210 ][ 292 ],
   alphaCSR[ 210 ][ 293 ],
   alphaCSR[ 210 ][ 294 ],
   alphaCSR[ 210 ][ 295 ],
   alphaCSR[ 210 ][ 296 ],
   alphaCSR[ 210 ][ 297 ],
   alphaCSR[ 210 ][ 298 ],
   alphaCSR[ 210 ][ 299 ],
   alphaCSR[ 210 ][ 300 ],
   alphaCSR[ 210 ][ 301 ],
   alphaCSR[ 210 ][ 302 ],
   alphaCSR[ 210 ][ 303 ],
   alphaCSR[ 210 ][ 304 ],
   alphaCSR[ 210 ][ 305 ],
   alphaCSR[ 210 ][ 306 ],
   alphaCSR[ 210 ][ 307 ],
   alphaCSR[ 210 ][ 308 ],
   alphaCSR[ 210 ][ 309 ],
   alphaCSR[ 210 ][ 310 ],
   alphaCSR[ 210 ][ 311 ],
   alphaCSR[ 210 ][ 312 ],
   alphaCSR[ 210 ][ 313 ],
   alphaCSR[ 210 ][ 314 ],
   alphaCSR[ 210 ][ 315 ],
   alphaCSR[ 210 ][ 316 ],
   alphaCSR[ 210 ][ 317 ],
   alphaCSR[ 210 ][ 318 ],
   alphaCSR[ 210 ][ 319 ],
   alphaCSR[ 210 ][ 320 ],
   alphaCSR[ 210 ][ 321 ],
   alphaCSR[ 210 ][ 322 ],
   alphaCSR[ 210 ][ 323 ],
   alphaCSR[ 210 ][ 324 ],
   alphaCSR[ 210 ][ 325 ],
   alphaCSR[ 210 ][ 326 ],
   alphaCSR[ 210 ][ 327 ],
   alphaCSR[ 210 ][ 328 ],
   alphaCSR[ 210 ][ 329 ],
   alphaCSR[ 210 ][ 330 ],
   alphaCSR[ 210 ][ 331 ],
   alphaCSR[ 210 ][ 332 ],
   alphaCSR[ 210 ][ 333 ],
   alphaCSR[ 210 ][ 334 ],
   alphaCSR[ 210 ][ 335 ],
   alphaCSR[ 210 ][ 336 ],
   alphaCSR[ 210 ][ 337 ],
   alphaCSR[ 210 ][ 338 ],
   alphaCSR[ 210 ][ 339 ],
   alphaCSR[ 210 ][ 340 ],
   alphaCSR[ 210 ][ 341 ],
   alphaCSR[ 210 ][ 342 ],
   alphaCSR[ 210 ][ 343 ],
   alphaCSR[ 210 ][ 344 ],
   alphaCSR[ 210 ][ 345 ],
   alphaCSR[ 210 ][ 346 ],
   alphaCSR[ 210 ][ 347 ],
   alphaCSR[ 210 ][ 348 ],
   alphaCSR[ 210 ][ 349 ],
   alphaCSR[ 210 ][ 350 ],
   alphaCSR[ 210 ][ 351 ],
   alphaCSR[ 210 ][ 352 ],
   alphaCSR[ 210 ][ 353 ],
   alphaCSR[ 210 ][ 354 ],
   alphaCSR[ 210 ][ 355 ],
   alphaCSR[ 210 ][ 356 ],
   alphaCSR[ 210 ][ 357 ],
   alphaCSR[ 210 ][ 358 ],
   alphaCSR[ 210 ][ 359 ],
   alphaCSR[ 210 ][ 360 ],
   alphaCSR[ 210 ][ 361 ],
   alphaCSR[ 210 ][ 362 ],
   alphaCSR[ 210 ][ 363 ],
   alphaCSR[ 210 ][ 364 ],
   alphaCSR[ 210 ][ 365 ],
   alphaCSR[ 210 ][ 366 ],
   alphaCSR[ 210 ][ 367 ],
   alphaCSR[ 210 ][ 368 ],
   alphaCSR[ 210 ][ 369 ],
   alphaCSR[ 210 ][ 370 ],
   alphaCSR[ 210 ][ 371 ],
   alphaCSR[ 210 ][ 372 ],
   alphaCSR[ 210 ][ 373 ],
   alphaCSR[ 210 ][ 374 ],
   alphaCSR[ 210 ][ 375 ],
   alphaCSR[ 210 ][ 376 ],
   alphaCSR[ 210 ][ 377 ],
   alphaCSR[ 210 ][ 378 ],
   alphaCSR[ 210 ][ 379 ],
   alphaCSR[ 210 ][ 380 ],
   alphaCSR[ 210 ][ 381 ],
   alphaCSR[ 210 ][ 382 ],
   alphaCSR[ 210 ][ 383 ],
   alphaCSR[ 211 ][ 0 ],
   alphaCSR[ 211 ][ 1 ],
   alphaCSR[ 211 ][ 2 ],
   alphaCSR[ 211 ][ 3 ],
   alphaCSR[ 211 ][ 4 ],
   alphaCSR[ 211 ][ 5 ],
   alphaCSR[ 211 ][ 6 ],
   alphaCSR[ 211 ][ 7 ],
   alphaCSR[ 211 ][ 8 ],
   alphaCSR[ 211 ][ 9 ],
   alphaCSR[ 211 ][ 10 ],
   alphaCSR[ 211 ][ 11 ],
   alphaCSR[ 211 ][ 12 ],
   alphaCSR[ 211 ][ 13 ],
   alphaCSR[ 211 ][ 14 ],
   alphaCSR[ 211 ][ 15 ],
   alphaCSR[ 211 ][ 16 ],
   alphaCSR[ 211 ][ 17 ],
   alphaCSR[ 211 ][ 18 ],
   alphaCSR[ 211 ][ 19 ],
   alphaCSR[ 211 ][ 20 ],
   alphaCSR[ 211 ][ 21 ],
   alphaCSR[ 211 ][ 22 ],
   alphaCSR[ 211 ][ 23 ],
   alphaCSR[ 211 ][ 24 ],
   alphaCSR[ 211 ][ 25 ],
   alphaCSR[ 211 ][ 26 ],
   alphaCSR[ 211 ][ 27 ],
   alphaCSR[ 211 ][ 28 ],
   alphaCSR[ 211 ][ 29 ],
   alphaCSR[ 211 ][ 30 ],
   alphaCSR[ 211 ][ 31 ],
   alphaCSR[ 211 ][ 32 ],
   alphaCSR[ 211 ][ 33 ],
   alphaCSR[ 211 ][ 34 ],
   alphaCSR[ 211 ][ 35 ],
   alphaCSR[ 211 ][ 36 ],
   alphaCSR[ 211 ][ 37 ],
   alphaCSR[ 211 ][ 38 ],
   alphaCSR[ 211 ][ 39 ],
   alphaCSR[ 211 ][ 40 ],
   alphaCSR[ 211 ][ 41 ],
   alphaCSR[ 211 ][ 42 ],
   alphaCSR[ 211 ][ 43 ],
   alphaCSR[ 211 ][ 44 ],
   alphaCSR[ 211 ][ 45 ],
   alphaCSR[ 211 ][ 46 ],
   alphaCSR[ 211 ][ 47 ],
   alphaCSR[ 211 ][ 48 ],
   alphaCSR[ 211 ][ 49 ],
   alphaCSR[ 211 ][ 50 ],
   alphaCSR[ 211 ][ 51 ],
   alphaCSR[ 211 ][ 52 ],
   alphaCSR[ 211 ][ 53 ],
   alphaCSR[ 211 ][ 54 ],
   alphaCSR[ 211 ][ 55 ],
   alphaCSR[ 211 ][ 56 ],
   alphaCSR[ 211 ][ 57 ],
   alphaCSR[ 211 ][ 58 ],
   alphaCSR[ 211 ][ 59 ],
   alphaCSR[ 211 ][ 60 ],
   alphaCSR[ 211 ][ 61 ],
   alphaCSR[ 211 ][ 62 ],
   alphaCSR[ 211 ][ 63 ],
   alphaCSR[ 211 ][ 64 ],
   alphaCSR[ 211 ][ 65 ],
   alphaCSR[ 211 ][ 66 ],
   alphaCSR[ 211 ][ 67 ],
   alphaCSR[ 211 ][ 68 ],
   alphaCSR[ 211 ][ 69 ],
   alphaCSR[ 211 ][ 70 ],
   alphaCSR[ 211 ][ 71 ],
   alphaCSR[ 211 ][ 72 ],
   alphaCSR[ 211 ][ 73 ],
   alphaCSR[ 211 ][ 74 ],
   alphaCSR[ 211 ][ 75 ],
   alphaCSR[ 211 ][ 76 ],
   alphaCSR[ 211 ][ 77 ],
   alphaCSR[ 211 ][ 78 ],
   alphaCSR[ 211 ][ 79 ],
   alphaCSR[ 211 ][ 80 ],
   alphaCSR[ 211 ][ 81 ],
   alphaCSR[ 211 ][ 82 ],
   alphaCSR[ 211 ][ 83 ],
   alphaCSR[ 211 ][ 84 ],
   alphaCSR[ 211 ][ 85 ],
   alphaCSR[ 211 ][ 86 ],
   alphaCSR[ 211 ][ 87 ],
   alphaCSR[ 211 ][ 88 ],
   alphaCSR[ 211 ][ 89 ],
   alphaCSR[ 211 ][ 90 ],
   alphaCSR[ 211 ][ 91 ],
   alphaCSR[ 211 ][ 92 ],
   alphaCSR[ 211 ][ 93 ],
   alphaCSR[ 211 ][ 94 ],
   alphaCSR[ 211 ][ 95 ],
   alphaCSR[ 211 ][ 96 ],
   alphaCSR[ 211 ][ 97 ],
   alphaCSR[ 211 ][ 98 ],
   alphaCSR[ 211 ][ 99 ],
   alphaCSR[ 211 ][ 100 ],
   alphaCSR[ 211 ][ 101 ],
   alphaCSR[ 211 ][ 102 ],
   alphaCSR[ 211 ][ 103 ],
   alphaCSR[ 211 ][ 104 ],
   alphaCSR[ 211 ][ 105 ],
   alphaCSR[ 211 ][ 106 ],
   alphaCSR[ 211 ][ 107 ],
   alphaCSR[ 211 ][ 108 ],
   alphaCSR[ 211 ][ 109 ],
   alphaCSR[ 211 ][ 110 ],
   alphaCSR[ 211 ][ 111 ],
   alphaCSR[ 211 ][ 112 ],
   alphaCSR[ 211 ][ 113 ],
   alphaCSR[ 211 ][ 114 ],
   alphaCSR[ 211 ][ 115 ],
   alphaCSR[ 211 ][ 116 ],
   alphaCSR[ 211 ][ 117 ],
   alphaCSR[ 211 ][ 118 ],
   alphaCSR[ 211 ][ 119 ],
   alphaCSR[ 211 ][ 120 ],
   alphaCSR[ 211 ][ 121 ],
   alphaCSR[ 211 ][ 122 ],
   alphaCSR[ 211 ][ 123 ],
   alphaCSR[ 211 ][ 124 ],
   alphaCSR[ 211 ][ 125 ],
   alphaCSR[ 211 ][ 126 ],
   alphaCSR[ 211 ][ 127 ],
   alphaCSR[ 211 ][ 128 ],
   alphaCSR[ 211 ][ 129 ],
   alphaCSR[ 211 ][ 130 ],
   alphaCSR[ 211 ][ 131 ],
   alphaCSR[ 211 ][ 132 ],
   alphaCSR[ 211 ][ 133 ],
   alphaCSR[ 211 ][ 134 ],
   alphaCSR[ 211 ][ 135 ],
   alphaCSR[ 211 ][ 136 ],
   alphaCSR[ 211 ][ 137 ],
   alphaCSR[ 211 ][ 138 ],
   alphaCSR[ 211 ][ 139 ],
   alphaCSR[ 211 ][ 140 ],
   alphaCSR[ 211 ][ 141 ],
   alphaCSR[ 211 ][ 142 ],
   alphaCSR[ 211 ][ 143 ],
   alphaCSR[ 211 ][ 144 ],
   alphaCSR[ 211 ][ 145 ],
   alphaCSR[ 211 ][ 146 ],
   alphaCSR[ 211 ][ 147 ],
   alphaCSR[ 211 ][ 148 ],
   alphaCSR[ 211 ][ 149 ],
   alphaCSR[ 211 ][ 150 ],
   alphaCSR[ 211 ][ 151 ],
   alphaCSR[ 211 ][ 152 ],
   alphaCSR[ 211 ][ 153 ],
   alphaCSR[ 211 ][ 154 ],
   alphaCSR[ 211 ][ 155 ],
   alphaCSR[ 211 ][ 156 ],
   alphaCSR[ 211 ][ 157 ],
   alphaCSR[ 211 ][ 158 ],
   alphaCSR[ 211 ][ 159 ],
   alphaCSR[ 211 ][ 160 ],
   alphaCSR[ 211 ][ 161 ],
   alphaCSR[ 211 ][ 162 ],
   alphaCSR[ 211 ][ 163 ],
   alphaCSR[ 211 ][ 164 ],
   alphaCSR[ 211 ][ 165 ],
   alphaCSR[ 211 ][ 166 ],
   alphaCSR[ 211 ][ 167 ],
   alphaCSR[ 211 ][ 168 ],
   alphaCSR[ 211 ][ 169 ],
   alphaCSR[ 211 ][ 170 ],
   alphaCSR[ 211 ][ 171 ],
   alphaCSR[ 211 ][ 172 ],
   alphaCSR[ 211 ][ 173 ],
   alphaCSR[ 211 ][ 174 ],
   alphaCSR[ 211 ][ 175 ],
   alphaCSR[ 211 ][ 176 ],
   alphaCSR[ 211 ][ 177 ],
   alphaCSR[ 211 ][ 178 ],
   alphaCSR[ 211 ][ 179 ],
   alphaCSR[ 211 ][ 180 ],
   alphaCSR[ 211 ][ 181 ],
   alphaCSR[ 211 ][ 182 ],
   alphaCSR[ 211 ][ 183 ],
   alphaCSR[ 211 ][ 184 ],
   alphaCSR[ 211 ][ 185 ],
   alphaCSR[ 211 ][ 186 ],
   alphaCSR[ 211 ][ 187 ],
   alphaCSR[ 211 ][ 188 ],
   alphaCSR[ 211 ][ 189 ],
   alphaCSR[ 211 ][ 190 ],
   alphaCSR[ 211 ][ 191 ],
   alphaCSR[ 211 ][ 192 ],
   alphaCSR[ 211 ][ 193 ],
   alphaCSR[ 211 ][ 194 ],
   alphaCSR[ 211 ][ 195 ],
   alphaCSR[ 211 ][ 196 ],
   alphaCSR[ 211 ][ 197 ],
   alphaCSR[ 211 ][ 198 ],
   alphaCSR[ 211 ][ 199 ],
   alphaCSR[ 211 ][ 200 ],
   alphaCSR[ 211 ][ 201 ],
   alphaCSR[ 211 ][ 202 ],
   alphaCSR[ 211 ][ 203 ],
   alphaCSR[ 211 ][ 204 ],
   alphaCSR[ 211 ][ 205 ],
   alphaCSR[ 211 ][ 206 ],
   alphaCSR[ 211 ][ 207 ],
   alphaCSR[ 211 ][ 208 ],
   alphaCSR[ 211 ][ 209 ],
   alphaCSR[ 211 ][ 210 ],
   alphaCSR[ 211 ][ 211 ],
   alphaCSR[ 211 ][ 212 ],
   alphaCSR[ 211 ][ 213 ],
   alphaCSR[ 211 ][ 214 ],
   alphaCSR[ 211 ][ 215 ],
   alphaCSR[ 211 ][ 216 ],
   alphaCSR[ 211 ][ 217 ],
   alphaCSR[ 211 ][ 218 ],
   alphaCSR[ 211 ][ 219 ],
   alphaCSR[ 211 ][ 220 ],
   alphaCSR[ 211 ][ 221 ],
   alphaCSR[ 211 ][ 222 ],
   alphaCSR[ 211 ][ 223 ],
   alphaCSR[ 211 ][ 224 ],
   alphaCSR[ 211 ][ 225 ],
   alphaCSR[ 211 ][ 226 ],
   alphaCSR[ 211 ][ 227 ],
   alphaCSR[ 211 ][ 228 ],
   alphaCSR[ 211 ][ 229 ],
   alphaCSR[ 211 ][ 230 ],
   alphaCSR[ 211 ][ 231 ],
   alphaCSR[ 211 ][ 232 ],
   alphaCSR[ 211 ][ 233 ],
   alphaCSR[ 211 ][ 234 ],
   alphaCSR[ 211 ][ 235 ],
   alphaCSR[ 211 ][ 236 ],
   alphaCSR[ 211 ][ 237 ],
   alphaCSR[ 211 ][ 238 ],
   alphaCSR[ 211 ][ 239 ],
   alphaCSR[ 211 ][ 240 ],
   alphaCSR[ 211 ][ 241 ],
   alphaCSR[ 211 ][ 242 ],
   alphaCSR[ 211 ][ 243 ],
   alphaCSR[ 211 ][ 244 ],
   alphaCSR[ 211 ][ 245 ],
   alphaCSR[ 211 ][ 246 ],
   alphaCSR[ 211 ][ 247 ],
   alphaCSR[ 211 ][ 248 ],
   alphaCSR[ 211 ][ 249 ],
   alphaCSR[ 211 ][ 250 ],
   alphaCSR[ 211 ][ 251 ],
   alphaCSR[ 211 ][ 252 ],
   alphaCSR[ 211 ][ 253 ],
   alphaCSR[ 211 ][ 254 ],
   alphaCSR[ 211 ][ 255 ],
   alphaCSR[ 211 ][ 256 ],
   alphaCSR[ 211 ][ 257 ],
   alphaCSR[ 211 ][ 258 ],
   alphaCSR[ 211 ][ 259 ],
   alphaCSR[ 211 ][ 260 ],
   alphaCSR[ 211 ][ 261 ],
   alphaCSR[ 211 ][ 262 ],
   alphaCSR[ 211 ][ 263 ],
   alphaCSR[ 211 ][ 264 ],
   alphaCSR[ 211 ][ 265 ],
   alphaCSR[ 211 ][ 266 ],
   alphaCSR[ 211 ][ 267 ],
   alphaCSR[ 211 ][ 268 ],
   alphaCSR[ 211 ][ 269 ],
   alphaCSR[ 211 ][ 270 ],
   alphaCSR[ 211 ][ 271 ],
   alphaCSR[ 211 ][ 272 ],
   alphaCSR[ 211 ][ 273 ],
   alphaCSR[ 211 ][ 274 ],
   alphaCSR[ 211 ][ 275 ],
   alphaCSR[ 211 ][ 276 ],
   alphaCSR[ 211 ][ 277 ],
   alphaCSR[ 211 ][ 278 ],
   alphaCSR[ 211 ][ 279 ],
   alphaCSR[ 211 ][ 280 ],
   alphaCSR[ 211 ][ 281 ],
   alphaCSR[ 211 ][ 282 ],
   alphaCSR[ 211 ][ 283 ],
   alphaCSR[ 211 ][ 284 ],
   alphaCSR[ 211 ][ 285 ],
   alphaCSR[ 211 ][ 286 ],
   alphaCSR[ 211 ][ 287 ],
   alphaCSR[ 211 ][ 288 ],
   alphaCSR[ 211 ][ 289 ],
   alphaCSR[ 211 ][ 290 ],
   alphaCSR[ 211 ][ 291 ],
   alphaCSR[ 211 ][ 292 ],
   alphaCSR[ 211 ][ 293 ],
   alphaCSR[ 211 ][ 294 ],
   alphaCSR[ 211 ][ 295 ],
   alphaCSR[ 211 ][ 296 ],
   alphaCSR[ 211 ][ 297 ],
   alphaCSR[ 211 ][ 298 ],
   alphaCSR[ 211 ][ 299 ],
   alphaCSR[ 211 ][ 300 ],
   alphaCSR[ 211 ][ 301 ],
   alphaCSR[ 211 ][ 302 ],
   alphaCSR[ 211 ][ 303 ],
   alphaCSR[ 211 ][ 304 ],
   alphaCSR[ 211 ][ 305 ],
   alphaCSR[ 211 ][ 306 ],
   alphaCSR[ 211 ][ 307 ],
   alphaCSR[ 211 ][ 308 ],
   alphaCSR[ 211 ][ 309 ],
   alphaCSR[ 211 ][ 310 ],
   alphaCSR[ 211 ][ 311 ],
   alphaCSR[ 211 ][ 312 ],
   alphaCSR[ 211 ][ 313 ],
   alphaCSR[ 211 ][ 314 ],
   alphaCSR[ 211 ][ 315 ],
   alphaCSR[ 211 ][ 316 ],
   alphaCSR[ 211 ][ 317 ],
   alphaCSR[ 211 ][ 318 ],
   alphaCSR[ 211 ][ 319 ],
   alphaCSR[ 211 ][ 320 ],
   alphaCSR[ 211 ][ 321 ],
   alphaCSR[ 211 ][ 322 ],
   alphaCSR[ 211 ][ 323 ],
   alphaCSR[ 211 ][ 324 ],
   alphaCSR[ 211 ][ 325 ],
   alphaCSR[ 211 ][ 326 ],
   alphaCSR[ 211 ][ 327 ],
   alphaCSR[ 211 ][ 328 ],
   alphaCSR[ 211 ][ 329 ],
   alphaCSR[ 211 ][ 330 ],
   alphaCSR[ 211 ][ 331 ],
   alphaCSR[ 211 ][ 332 ],
   alphaCSR[ 211 ][ 333 ],
   alphaCSR[ 211 ][ 334 ],
   alphaCSR[ 211 ][ 335 ],
   alphaCSR[ 211 ][ 336 ],
   alphaCSR[ 211 ][ 337 ],
   alphaCSR[ 211 ][ 338 ],
   alphaCSR[ 211 ][ 339 ],
   alphaCSR[ 211 ][ 340 ],
   alphaCSR[ 211 ][ 341 ],
   alphaCSR[ 211 ][ 342 ],
   alphaCSR[ 211 ][ 343 ],
   alphaCSR[ 211 ][ 344 ],
   alphaCSR[ 211 ][ 345 ],
   alphaCSR[ 211 ][ 346 ],
   alphaCSR[ 211 ][ 347 ],
   alphaCSR[ 211 ][ 348 ],
   alphaCSR[ 211 ][ 349 ],
   alphaCSR[ 211 ][ 350 ],
   alphaCSR[ 211 ][ 351 ],
   alphaCSR[ 211 ][ 352 ],
   alphaCSR[ 211 ][ 353 ],
   alphaCSR[ 211 ][ 354 ],
   alphaCSR[ 211 ][ 355 ],
   alphaCSR[ 211 ][ 356 ],
   alphaCSR[ 211 ][ 357 ],
   alphaCSR[ 211 ][ 358 ],
   alphaCSR[ 211 ][ 359 ],
   alphaCSR[ 211 ][ 360 ],
   alphaCSR[ 211 ][ 361 ],
   alphaCSR[ 211 ][ 362 ],
   alphaCSR[ 211 ][ 363 ],
   alphaCSR[ 211 ][ 364 ],
   alphaCSR[ 211 ][ 365 ],
   alphaCSR[ 211 ][ 366 ],
   alphaCSR[ 211 ][ 367 ],
   alphaCSR[ 211 ][ 368 ],
   alphaCSR[ 211 ][ 369 ],
   alphaCSR[ 211 ][ 370 ],
   alphaCSR[ 211 ][ 371 ],
   alphaCSR[ 211 ][ 372 ],
   alphaCSR[ 211 ][ 373 ],
   alphaCSR[ 211 ][ 374 ],
   alphaCSR[ 211 ][ 375 ],
   alphaCSR[ 211 ][ 376 ],
   alphaCSR[ 211 ][ 377 ],
   alphaCSR[ 211 ][ 378 ],
   alphaCSR[ 211 ][ 379 ],
   alphaCSR[ 211 ][ 380 ],
   alphaCSR[ 211 ][ 381 ],
   alphaCSR[ 211 ][ 382 ],
   alphaCSR[ 211 ][ 383 ],
   alphaCSR[ 212 ][ 0 ],
   alphaCSR[ 212 ][ 1 ],
   alphaCSR[ 212 ][ 2 ],
   alphaCSR[ 212 ][ 3 ],
   alphaCSR[ 212 ][ 4 ],
   alphaCSR[ 212 ][ 5 ],
   alphaCSR[ 212 ][ 6 ],
   alphaCSR[ 212 ][ 7 ],
   alphaCSR[ 212 ][ 8 ],
   alphaCSR[ 212 ][ 9 ],
   alphaCSR[ 212 ][ 10 ],
   alphaCSR[ 212 ][ 11 ],
   alphaCSR[ 212 ][ 12 ],
   alphaCSR[ 212 ][ 13 ],
   alphaCSR[ 212 ][ 14 ],
   alphaCSR[ 212 ][ 15 ],
   alphaCSR[ 212 ][ 16 ],
   alphaCSR[ 212 ][ 17 ],
   alphaCSR[ 212 ][ 18 ],
   alphaCSR[ 212 ][ 19 ],
   alphaCSR[ 212 ][ 20 ],
   alphaCSR[ 212 ][ 21 ],
   alphaCSR[ 212 ][ 22 ],
   alphaCSR[ 212 ][ 23 ],
   alphaCSR[ 212 ][ 24 ],
   alphaCSR[ 212 ][ 25 ],
   alphaCSR[ 212 ][ 26 ],
   alphaCSR[ 212 ][ 27 ],
   alphaCSR[ 212 ][ 28 ],
   alphaCSR[ 212 ][ 29 ],
   alphaCSR[ 212 ][ 30 ],
   alphaCSR[ 212 ][ 31 ],
   alphaCSR[ 212 ][ 32 ],
   alphaCSR[ 212 ][ 33 ],
   alphaCSR[ 212 ][ 34 ],
   alphaCSR[ 212 ][ 35 ],
   alphaCSR[ 212 ][ 36 ],
   alphaCSR[ 212 ][ 37 ],
   alphaCSR[ 212 ][ 38 ],
   alphaCSR[ 212 ][ 39 ],
   alphaCSR[ 212 ][ 40 ],
   alphaCSR[ 212 ][ 41 ],
   alphaCSR[ 212 ][ 42 ],
   alphaCSR[ 212 ][ 43 ],
   alphaCSR[ 212 ][ 44 ],
   alphaCSR[ 212 ][ 45 ],
   alphaCSR[ 212 ][ 46 ],
   alphaCSR[ 212 ][ 47 ],
   alphaCSR[ 212 ][ 48 ],
   alphaCSR[ 212 ][ 49 ],
   alphaCSR[ 212 ][ 50 ],
   alphaCSR[ 212 ][ 51 ],
   alphaCSR[ 212 ][ 52 ],
   alphaCSR[ 212 ][ 53 ],
   alphaCSR[ 212 ][ 54 ],
   alphaCSR[ 212 ][ 55 ],
   alphaCSR[ 212 ][ 56 ],
   alphaCSR[ 212 ][ 57 ],
   alphaCSR[ 212 ][ 58 ],
   alphaCSR[ 212 ][ 59 ],
   alphaCSR[ 212 ][ 60 ],
   alphaCSR[ 212 ][ 61 ],
   alphaCSR[ 212 ][ 62 ],
   alphaCSR[ 212 ][ 63 ],
   alphaCSR[ 212 ][ 64 ],
   alphaCSR[ 212 ][ 65 ],
   alphaCSR[ 212 ][ 66 ],
   alphaCSR[ 212 ][ 67 ],
   alphaCSR[ 212 ][ 68 ],
   alphaCSR[ 212 ][ 69 ],
   alphaCSR[ 212 ][ 70 ],
   alphaCSR[ 212 ][ 71 ],
   alphaCSR[ 212 ][ 72 ],
   alphaCSR[ 212 ][ 73 ],
   alphaCSR[ 212 ][ 74 ],
   alphaCSR[ 212 ][ 75 ],
   alphaCSR[ 212 ][ 76 ],
   alphaCSR[ 212 ][ 77 ],
   alphaCSR[ 212 ][ 78 ],
   alphaCSR[ 212 ][ 79 ],
   alphaCSR[ 212 ][ 80 ],
   alphaCSR[ 212 ][ 81 ],
   alphaCSR[ 212 ][ 82 ],
   alphaCSR[ 212 ][ 83 ],
   alphaCSR[ 212 ][ 84 ],
   alphaCSR[ 212 ][ 85 ],
   alphaCSR[ 212 ][ 86 ],
   alphaCSR[ 212 ][ 87 ],
   alphaCSR[ 212 ][ 88 ],
   alphaCSR[ 212 ][ 89 ],
   alphaCSR[ 212 ][ 90 ],
   alphaCSR[ 212 ][ 91 ],
   alphaCSR[ 212 ][ 92 ],
   alphaCSR[ 212 ][ 93 ],
   alphaCSR[ 212 ][ 94 ],
   alphaCSR[ 212 ][ 95 ],
   alphaCSR[ 212 ][ 96 ],
   alphaCSR[ 212 ][ 97 ],
   alphaCSR[ 212 ][ 98 ],
   alphaCSR[ 212 ][ 99 ],
   alphaCSR[ 212 ][ 100 ],
   alphaCSR[ 212 ][ 101 ],
   alphaCSR[ 212 ][ 102 ],
   alphaCSR[ 212 ][ 103 ],
   alphaCSR[ 212 ][ 104 ],
   alphaCSR[ 212 ][ 105 ],
   alphaCSR[ 212 ][ 106 ],
   alphaCSR[ 212 ][ 107 ],
   alphaCSR[ 212 ][ 108 ],
   alphaCSR[ 212 ][ 109 ],
   alphaCSR[ 212 ][ 110 ],
   alphaCSR[ 212 ][ 111 ],
   alphaCSR[ 212 ][ 112 ],
   alphaCSR[ 212 ][ 113 ],
   alphaCSR[ 212 ][ 114 ],
   alphaCSR[ 212 ][ 115 ],
   alphaCSR[ 212 ][ 116 ],
   alphaCSR[ 212 ][ 117 ],
   alphaCSR[ 212 ][ 118 ],
   alphaCSR[ 212 ][ 119 ],
   alphaCSR[ 212 ][ 120 ],
   alphaCSR[ 212 ][ 121 ],
   alphaCSR[ 212 ][ 122 ],
   alphaCSR[ 212 ][ 123 ],
   alphaCSR[ 212 ][ 124 ],
   alphaCSR[ 212 ][ 125 ],
   alphaCSR[ 212 ][ 126 ],
   alphaCSR[ 212 ][ 127 ],
   alphaCSR[ 212 ][ 128 ],
   alphaCSR[ 212 ][ 129 ],
   alphaCSR[ 212 ][ 130 ],
   alphaCSR[ 212 ][ 131 ],
   alphaCSR[ 212 ][ 132 ],
   alphaCSR[ 212 ][ 133 ],
   alphaCSR[ 212 ][ 134 ],
   alphaCSR[ 212 ][ 135 ],
   alphaCSR[ 212 ][ 136 ],
   alphaCSR[ 212 ][ 137 ],
   alphaCSR[ 212 ][ 138 ],
   alphaCSR[ 212 ][ 139 ],
   alphaCSR[ 212 ][ 140 ],
   alphaCSR[ 212 ][ 141 ],
   alphaCSR[ 212 ][ 142 ],
   alphaCSR[ 212 ][ 143 ],
   alphaCSR[ 212 ][ 144 ],
   alphaCSR[ 212 ][ 145 ],
   alphaCSR[ 212 ][ 146 ],
   alphaCSR[ 212 ][ 147 ],
   alphaCSR[ 212 ][ 148 ],
   alphaCSR[ 212 ][ 149 ],
   alphaCSR[ 212 ][ 150 ],
   alphaCSR[ 212 ][ 151 ],
   alphaCSR[ 212 ][ 152 ],
   alphaCSR[ 212 ][ 153 ],
   alphaCSR[ 212 ][ 154 ],
   alphaCSR[ 212 ][ 155 ],
   alphaCSR[ 212 ][ 156 ],
   alphaCSR[ 212 ][ 157 ],
   alphaCSR[ 212 ][ 158 ],
   alphaCSR[ 212 ][ 159 ],
   alphaCSR[ 212 ][ 160 ],
   alphaCSR[ 212 ][ 161 ],
   alphaCSR[ 212 ][ 162 ],
   alphaCSR[ 212 ][ 163 ],
   alphaCSR[ 212 ][ 164 ],
   alphaCSR[ 212 ][ 165 ],
   alphaCSR[ 212 ][ 166 ],
   alphaCSR[ 212 ][ 167 ],
   alphaCSR[ 212 ][ 168 ],
   alphaCSR[ 212 ][ 169 ],
   alphaCSR[ 212 ][ 170 ],
   alphaCSR[ 212 ][ 171 ],
   alphaCSR[ 212 ][ 172 ],
   alphaCSR[ 212 ][ 173 ],
   alphaCSR[ 212 ][ 174 ],
   alphaCSR[ 212 ][ 175 ],
   alphaCSR[ 212 ][ 176 ],
   alphaCSR[ 212 ][ 177 ],
   alphaCSR[ 212 ][ 178 ],
   alphaCSR[ 212 ][ 179 ],
   alphaCSR[ 212 ][ 180 ],
   alphaCSR[ 212 ][ 181 ],
   alphaCSR[ 212 ][ 182 ],
   alphaCSR[ 212 ][ 183 ],
   alphaCSR[ 212 ][ 184 ],
   alphaCSR[ 212 ][ 185 ],
   alphaCSR[ 212 ][ 186 ],
   alphaCSR[ 212 ][ 187 ],
   alphaCSR[ 212 ][ 188 ],
   alphaCSR[ 212 ][ 189 ],
   alphaCSR[ 212 ][ 190 ],
   alphaCSR[ 212 ][ 191 ],
   alphaCSR[ 212 ][ 192 ],
   alphaCSR[ 212 ][ 193 ],
   alphaCSR[ 212 ][ 194 ],
   alphaCSR[ 212 ][ 195 ],
   alphaCSR[ 212 ][ 196 ],
   alphaCSR[ 212 ][ 197 ],
   alphaCSR[ 212 ][ 198 ],
   alphaCSR[ 212 ][ 199 ],
   alphaCSR[ 212 ][ 200 ],
   alphaCSR[ 212 ][ 201 ],
   alphaCSR[ 212 ][ 202 ],
   alphaCSR[ 212 ][ 203 ],
   alphaCSR[ 212 ][ 204 ],
   alphaCSR[ 212 ][ 205 ],
   alphaCSR[ 212 ][ 206 ],
   alphaCSR[ 212 ][ 207 ],
   alphaCSR[ 212 ][ 208 ],
   alphaCSR[ 212 ][ 209 ],
   alphaCSR[ 212 ][ 210 ],
   alphaCSR[ 212 ][ 211 ],
   alphaCSR[ 212 ][ 212 ],
   alphaCSR[ 212 ][ 213 ],
   alphaCSR[ 212 ][ 214 ],
   alphaCSR[ 212 ][ 215 ],
   alphaCSR[ 212 ][ 216 ],
   alphaCSR[ 212 ][ 217 ],
   alphaCSR[ 212 ][ 218 ],
   alphaCSR[ 212 ][ 219 ],
   alphaCSR[ 212 ][ 220 ],
   alphaCSR[ 212 ][ 221 ],
   alphaCSR[ 212 ][ 222 ],
   alphaCSR[ 212 ][ 223 ],
   alphaCSR[ 212 ][ 224 ],
   alphaCSR[ 212 ][ 225 ],
   alphaCSR[ 212 ][ 226 ],
   alphaCSR[ 212 ][ 227 ],
   alphaCSR[ 212 ][ 228 ],
   alphaCSR[ 212 ][ 229 ],
   alphaCSR[ 212 ][ 230 ],
   alphaCSR[ 212 ][ 231 ],
   alphaCSR[ 212 ][ 232 ],
   alphaCSR[ 212 ][ 233 ],
   alphaCSR[ 212 ][ 234 ],
   alphaCSR[ 212 ][ 235 ],
   alphaCSR[ 212 ][ 236 ],
   alphaCSR[ 212 ][ 237 ],
   alphaCSR[ 212 ][ 238 ],
   alphaCSR[ 212 ][ 239 ],
   alphaCSR[ 212 ][ 240 ],
   alphaCSR[ 212 ][ 241 ],
   alphaCSR[ 212 ][ 242 ],
   alphaCSR[ 212 ][ 243 ],
   alphaCSR[ 212 ][ 244 ],
   alphaCSR[ 212 ][ 245 ],
   alphaCSR[ 212 ][ 246 ],
   alphaCSR[ 212 ][ 247 ],
   alphaCSR[ 212 ][ 248 ],
   alphaCSR[ 212 ][ 249 ],
   alphaCSR[ 212 ][ 250 ],
   alphaCSR[ 212 ][ 251 ],
   alphaCSR[ 212 ][ 252 ],
   alphaCSR[ 212 ][ 253 ],
   alphaCSR[ 212 ][ 254 ],
   alphaCSR[ 212 ][ 255 ],
   alphaCSR[ 212 ][ 256 ],
   alphaCSR[ 212 ][ 257 ],
   alphaCSR[ 212 ][ 258 ],
   alphaCSR[ 212 ][ 259 ],
   alphaCSR[ 212 ][ 260 ],
   alphaCSR[ 212 ][ 261 ],
   alphaCSR[ 212 ][ 262 ],
   alphaCSR[ 212 ][ 263 ],
   alphaCSR[ 212 ][ 264 ],
   alphaCSR[ 212 ][ 265 ],
   alphaCSR[ 212 ][ 266 ],
   alphaCSR[ 212 ][ 267 ],
   alphaCSR[ 212 ][ 268 ],
   alphaCSR[ 212 ][ 269 ],
   alphaCSR[ 212 ][ 270 ],
   alphaCSR[ 212 ][ 271 ],
   alphaCSR[ 212 ][ 272 ],
   alphaCSR[ 212 ][ 273 ],
   alphaCSR[ 212 ][ 274 ],
   alphaCSR[ 212 ][ 275 ],
   alphaCSR[ 212 ][ 276 ],
   alphaCSR[ 212 ][ 277 ],
   alphaCSR[ 212 ][ 278 ],
   alphaCSR[ 212 ][ 279 ],
   alphaCSR[ 212 ][ 280 ],
   alphaCSR[ 212 ][ 281 ],
   alphaCSR[ 212 ][ 282 ],
   alphaCSR[ 212 ][ 283 ],
   alphaCSR[ 212 ][ 284 ],
   alphaCSR[ 212 ][ 285 ],
   alphaCSR[ 212 ][ 286 ],
   alphaCSR[ 212 ][ 287 ],
   alphaCSR[ 212 ][ 288 ],
   alphaCSR[ 212 ][ 289 ],
   alphaCSR[ 212 ][ 290 ],
   alphaCSR[ 212 ][ 291 ],
   alphaCSR[ 212 ][ 292 ],
   alphaCSR[ 212 ][ 293 ],
   alphaCSR[ 212 ][ 294 ],
   alphaCSR[ 212 ][ 295 ],
   alphaCSR[ 212 ][ 296 ],
   alphaCSR[ 212 ][ 297 ],
   alphaCSR[ 212 ][ 298 ],
   alphaCSR[ 212 ][ 299 ],
   alphaCSR[ 212 ][ 300 ],
   alphaCSR[ 212 ][ 301 ],
   alphaCSR[ 212 ][ 302 ],
   alphaCSR[ 212 ][ 303 ],
   alphaCSR[ 212 ][ 304 ],
   alphaCSR[ 212 ][ 305 ],
   alphaCSR[ 212 ][ 306 ],
   alphaCSR[ 212 ][ 307 ],
   alphaCSR[ 212 ][ 308 ],
   alphaCSR[ 212 ][ 309 ],
   alphaCSR[ 212 ][ 310 ],
   alphaCSR[ 212 ][ 311 ],
   alphaCSR[ 212 ][ 312 ],
   alphaCSR[ 212 ][ 313 ],
   alphaCSR[ 212 ][ 314 ],
   alphaCSR[ 212 ][ 315 ],
   alphaCSR[ 212 ][ 316 ],
   alphaCSR[ 212 ][ 317 ],
   alphaCSR[ 212 ][ 318 ],
   alphaCSR[ 212 ][ 319 ],
   alphaCSR[ 212 ][ 320 ],
   alphaCSR[ 212 ][ 321 ],
   alphaCSR[ 212 ][ 322 ],
   alphaCSR[ 212 ][ 323 ],
   alphaCSR[ 212 ][ 324 ],
   alphaCSR[ 212 ][ 325 ],
   alphaCSR[ 212 ][ 326 ],
   alphaCSR[ 212 ][ 327 ],
   alphaCSR[ 212 ][ 328 ],
   alphaCSR[ 212 ][ 329 ],
   alphaCSR[ 212 ][ 330 ],
   alphaCSR[ 212 ][ 331 ],
   alphaCSR[ 212 ][ 332 ],
   alphaCSR[ 212 ][ 333 ],
   alphaCSR[ 212 ][ 334 ],
   alphaCSR[ 212 ][ 335 ],
   alphaCSR[ 212 ][ 336 ],
   alphaCSR[ 212 ][ 337 ],
   alphaCSR[ 212 ][ 338 ],
   alphaCSR[ 212 ][ 339 ],
   alphaCSR[ 212 ][ 340 ],
   alphaCSR[ 212 ][ 341 ],
   alphaCSR[ 212 ][ 342 ],
   alphaCSR[ 212 ][ 343 ],
   alphaCSR[ 212 ][ 344 ],
   alphaCSR[ 212 ][ 345 ],
   alphaCSR[ 212 ][ 346 ],
   alphaCSR[ 212 ][ 347 ],
   alphaCSR[ 212 ][ 348 ],
   alphaCSR[ 212 ][ 349 ],
   alphaCSR[ 212 ][ 350 ],
   alphaCSR[ 212 ][ 351 ],
   alphaCSR[ 212 ][ 352 ],
   alphaCSR[ 212 ][ 353 ],
   alphaCSR[ 212 ][ 354 ],
   alphaCSR[ 212 ][ 355 ],
   alphaCSR[ 212 ][ 356 ],
   alphaCSR[ 212 ][ 357 ],
   alphaCSR[ 212 ][ 358 ],
   alphaCSR[ 212 ][ 359 ],
   alphaCSR[ 212 ][ 360 ],
   alphaCSR[ 212 ][ 361 ],
   alphaCSR[ 212 ][ 362 ],
   alphaCSR[ 212 ][ 363 ],
   alphaCSR[ 212 ][ 364 ],
   alphaCSR[ 212 ][ 365 ],
   alphaCSR[ 212 ][ 366 ],
   alphaCSR[ 212 ][ 367 ],
   alphaCSR[ 212 ][ 368 ],
   alphaCSR[ 212 ][ 369 ],
   alphaCSR[ 212 ][ 370 ],
   alphaCSR[ 212 ][ 371 ],
   alphaCSR[ 212 ][ 372 ],
   alphaCSR[ 212 ][ 373 ],
   alphaCSR[ 212 ][ 374 ],
   alphaCSR[ 212 ][ 375 ],
   alphaCSR[ 212 ][ 376 ],
   alphaCSR[ 212 ][ 377 ],
   alphaCSR[ 212 ][ 378 ],
   alphaCSR[ 212 ][ 379 ],
   alphaCSR[ 212 ][ 380 ],
   alphaCSR[ 212 ][ 381 ],
   alphaCSR[ 212 ][ 382 ],
   alphaCSR[ 212 ][ 383 ],
   alphaCSR[ 213 ][ 0 ],
   alphaCSR[ 213 ][ 1 ],
   alphaCSR[ 213 ][ 2 ],
   alphaCSR[ 213 ][ 3 ],
   alphaCSR[ 213 ][ 4 ],
   alphaCSR[ 213 ][ 5 ],
   alphaCSR[ 213 ][ 6 ],
   alphaCSR[ 213 ][ 7 ],
   alphaCSR[ 213 ][ 8 ],
   alphaCSR[ 213 ][ 9 ],
   alphaCSR[ 213 ][ 10 ],
   alphaCSR[ 213 ][ 11 ],
   alphaCSR[ 213 ][ 12 ],
   alphaCSR[ 213 ][ 13 ],
   alphaCSR[ 213 ][ 14 ],
   alphaCSR[ 213 ][ 15 ],
   alphaCSR[ 213 ][ 16 ],
   alphaCSR[ 213 ][ 17 ],
   alphaCSR[ 213 ][ 18 ],
   alphaCSR[ 213 ][ 19 ],
   alphaCSR[ 213 ][ 20 ],
   alphaCSR[ 213 ][ 21 ],
   alphaCSR[ 213 ][ 22 ],
   alphaCSR[ 213 ][ 23 ],
   alphaCSR[ 213 ][ 24 ],
   alphaCSR[ 213 ][ 25 ],
   alphaCSR[ 213 ][ 26 ],
   alphaCSR[ 213 ][ 27 ],
   alphaCSR[ 213 ][ 28 ],
   alphaCSR[ 213 ][ 29 ],
   alphaCSR[ 213 ][ 30 ],
   alphaCSR[ 213 ][ 31 ],
   alphaCSR[ 213 ][ 32 ],
   alphaCSR[ 213 ][ 33 ],
   alphaCSR[ 213 ][ 34 ],
   alphaCSR[ 213 ][ 35 ],
   alphaCSR[ 213 ][ 36 ],
   alphaCSR[ 213 ][ 37 ],
   alphaCSR[ 213 ][ 38 ],
   alphaCSR[ 213 ][ 39 ],
   alphaCSR[ 213 ][ 40 ],
   alphaCSR[ 213 ][ 41 ],
   alphaCSR[ 213 ][ 42 ],
   alphaCSR[ 213 ][ 43 ],
   alphaCSR[ 213 ][ 44 ],
   alphaCSR[ 213 ][ 45 ],
   alphaCSR[ 213 ][ 46 ],
   alphaCSR[ 213 ][ 47 ],
   alphaCSR[ 213 ][ 48 ],
   alphaCSR[ 213 ][ 49 ],
   alphaCSR[ 213 ][ 50 ],
   alphaCSR[ 213 ][ 51 ],
   alphaCSR[ 213 ][ 52 ],
   alphaCSR[ 213 ][ 53 ],
   alphaCSR[ 213 ][ 54 ],
   alphaCSR[ 213 ][ 55 ],
   alphaCSR[ 213 ][ 56 ],
   alphaCSR[ 213 ][ 57 ],
   alphaCSR[ 213 ][ 58 ],
   alphaCSR[ 213 ][ 59 ],
   alphaCSR[ 213 ][ 60 ],
   alphaCSR[ 213 ][ 61 ],
   alphaCSR[ 213 ][ 62 ],
   alphaCSR[ 213 ][ 63 ],
   alphaCSR[ 213 ][ 64 ],
   alphaCSR[ 213 ][ 65 ],
   alphaCSR[ 213 ][ 66 ],
   alphaCSR[ 213 ][ 67 ],
   alphaCSR[ 213 ][ 68 ],
   alphaCSR[ 213 ][ 69 ],
   alphaCSR[ 213 ][ 70 ],
   alphaCSR[ 213 ][ 71 ],
   alphaCSR[ 213 ][ 72 ],
   alphaCSR[ 213 ][ 73 ],
   alphaCSR[ 213 ][ 74 ],
   alphaCSR[ 213 ][ 75 ],
   alphaCSR[ 213 ][ 76 ],
   alphaCSR[ 213 ][ 77 ],
   alphaCSR[ 213 ][ 78 ],
   alphaCSR[ 213 ][ 79 ],
   alphaCSR[ 213 ][ 80 ],
   alphaCSR[ 213 ][ 81 ],
   alphaCSR[ 213 ][ 82 ],
   alphaCSR[ 213 ][ 83 ],
   alphaCSR[ 213 ][ 84 ],
   alphaCSR[ 213 ][ 85 ],
   alphaCSR[ 213 ][ 86 ],
   alphaCSR[ 213 ][ 87 ],
   alphaCSR[ 213 ][ 88 ],
   alphaCSR[ 213 ][ 89 ],
   alphaCSR[ 213 ][ 90 ],
   alphaCSR[ 213 ][ 91 ],
   alphaCSR[ 213 ][ 92 ],
   alphaCSR[ 213 ][ 93 ],
   alphaCSR[ 213 ][ 94 ],
   alphaCSR[ 213 ][ 95 ],
   alphaCSR[ 213 ][ 96 ],
   alphaCSR[ 213 ][ 97 ],
   alphaCSR[ 213 ][ 98 ],
   alphaCSR[ 213 ][ 99 ],
   alphaCSR[ 213 ][ 100 ],
   alphaCSR[ 213 ][ 101 ],
   alphaCSR[ 213 ][ 102 ],
   alphaCSR[ 213 ][ 103 ],
   alphaCSR[ 213 ][ 104 ],
   alphaCSR[ 213 ][ 105 ],
   alphaCSR[ 213 ][ 106 ],
   alphaCSR[ 213 ][ 107 ],
   alphaCSR[ 213 ][ 108 ],
   alphaCSR[ 213 ][ 109 ],
   alphaCSR[ 213 ][ 110 ],
   alphaCSR[ 213 ][ 111 ],
   alphaCSR[ 213 ][ 112 ],
   alphaCSR[ 213 ][ 113 ],
   alphaCSR[ 213 ][ 114 ],
   alphaCSR[ 213 ][ 115 ],
   alphaCSR[ 213 ][ 116 ],
   alphaCSR[ 213 ][ 117 ],
   alphaCSR[ 213 ][ 118 ],
   alphaCSR[ 213 ][ 119 ],
   alphaCSR[ 213 ][ 120 ],
   alphaCSR[ 213 ][ 121 ],
   alphaCSR[ 213 ][ 122 ],
   alphaCSR[ 213 ][ 123 ],
   alphaCSR[ 213 ][ 124 ],
   alphaCSR[ 213 ][ 125 ],
   alphaCSR[ 213 ][ 126 ],
   alphaCSR[ 213 ][ 127 ],
   alphaCSR[ 213 ][ 128 ],
   alphaCSR[ 213 ][ 129 ],
   alphaCSR[ 213 ][ 130 ],
   alphaCSR[ 213 ][ 131 ],
   alphaCSR[ 213 ][ 132 ],
   alphaCSR[ 213 ][ 133 ],
   alphaCSR[ 213 ][ 134 ],
   alphaCSR[ 213 ][ 135 ],
   alphaCSR[ 213 ][ 136 ],
   alphaCSR[ 213 ][ 137 ],
   alphaCSR[ 213 ][ 138 ],
   alphaCSR[ 213 ][ 139 ],
   alphaCSR[ 213 ][ 140 ],
   alphaCSR[ 213 ][ 141 ],
   alphaCSR[ 213 ][ 142 ],
   alphaCSR[ 213 ][ 143 ],
   alphaCSR[ 213 ][ 144 ],
   alphaCSR[ 213 ][ 145 ],
   alphaCSR[ 213 ][ 146 ],
   alphaCSR[ 213 ][ 147 ],
   alphaCSR[ 213 ][ 148 ],
   alphaCSR[ 213 ][ 149 ],
   alphaCSR[ 213 ][ 150 ],
   alphaCSR[ 213 ][ 151 ],
   alphaCSR[ 213 ][ 152 ],
   alphaCSR[ 213 ][ 153 ],
   alphaCSR[ 213 ][ 154 ],
   alphaCSR[ 213 ][ 155 ],
   alphaCSR[ 213 ][ 156 ],
   alphaCSR[ 213 ][ 157 ],
   alphaCSR[ 213 ][ 158 ],
   alphaCSR[ 213 ][ 159 ],
   alphaCSR[ 213 ][ 160 ],
   alphaCSR[ 213 ][ 161 ],
   alphaCSR[ 213 ][ 162 ],
   alphaCSR[ 213 ][ 163 ],
   alphaCSR[ 213 ][ 164 ],
   alphaCSR[ 213 ][ 165 ],
   alphaCSR[ 213 ][ 166 ],
   alphaCSR[ 213 ][ 167 ],
   alphaCSR[ 213 ][ 168 ],
   alphaCSR[ 213 ][ 169 ],
   alphaCSR[ 213 ][ 170 ],
   alphaCSR[ 213 ][ 171 ],
   alphaCSR[ 213 ][ 172 ],
   alphaCSR[ 213 ][ 173 ],
   alphaCSR[ 213 ][ 174 ],
   alphaCSR[ 213 ][ 175 ],
   alphaCSR[ 213 ][ 176 ],
   alphaCSR[ 213 ][ 177 ],
   alphaCSR[ 213 ][ 178 ],
   alphaCSR[ 213 ][ 179 ],
   alphaCSR[ 213 ][ 180 ],
   alphaCSR[ 213 ][ 181 ],
   alphaCSR[ 213 ][ 182 ],
   alphaCSR[ 213 ][ 183 ],
   alphaCSR[ 213 ][ 184 ],
   alphaCSR[ 213 ][ 185 ],
   alphaCSR[ 213 ][ 186 ],
   alphaCSR[ 213 ][ 187 ],
   alphaCSR[ 213 ][ 188 ],
   alphaCSR[ 213 ][ 189 ],
   alphaCSR[ 213 ][ 190 ],
   alphaCSR[ 213 ][ 191 ],
   alphaCSR[ 213 ][ 192 ],
   alphaCSR[ 213 ][ 193 ],
   alphaCSR[ 213 ][ 194 ],
   alphaCSR[ 213 ][ 195 ],
   alphaCSR[ 213 ][ 196 ],
   alphaCSR[ 213 ][ 197 ],
   alphaCSR[ 213 ][ 198 ],
   alphaCSR[ 213 ][ 199 ],
   alphaCSR[ 213 ][ 200 ],
   alphaCSR[ 213 ][ 201 ],
   alphaCSR[ 213 ][ 202 ],
   alphaCSR[ 213 ][ 203 ],
   alphaCSR[ 213 ][ 204 ],
   alphaCSR[ 213 ][ 205 ],
   alphaCSR[ 213 ][ 206 ],
   alphaCSR[ 213 ][ 207 ],
   alphaCSR[ 213 ][ 208 ],
   alphaCSR[ 213 ][ 209 ],
   alphaCSR[ 213 ][ 210 ],
   alphaCSR[ 213 ][ 211 ],
   alphaCSR[ 213 ][ 212 ],
   alphaCSR[ 213 ][ 213 ],
   alphaCSR[ 213 ][ 214 ],
   alphaCSR[ 213 ][ 215 ],
   alphaCSR[ 213 ][ 216 ],
   alphaCSR[ 213 ][ 217 ],
   alphaCSR[ 213 ][ 218 ],
   alphaCSR[ 213 ][ 219 ],
   alphaCSR[ 213 ][ 220 ],
   alphaCSR[ 213 ][ 221 ],
   alphaCSR[ 213 ][ 222 ],
   alphaCSR[ 213 ][ 223 ],
   alphaCSR[ 213 ][ 224 ],
   alphaCSR[ 213 ][ 225 ],
   alphaCSR[ 213 ][ 226 ],
   alphaCSR[ 213 ][ 227 ],
   alphaCSR[ 213 ][ 228 ],
   alphaCSR[ 213 ][ 229 ],
   alphaCSR[ 213 ][ 230 ],
   alphaCSR[ 213 ][ 231 ],
   alphaCSR[ 213 ][ 232 ],
   alphaCSR[ 213 ][ 233 ],
   alphaCSR[ 213 ][ 234 ],
   alphaCSR[ 213 ][ 235 ],
   alphaCSR[ 213 ][ 236 ],
   alphaCSR[ 213 ][ 237 ],
   alphaCSR[ 213 ][ 238 ],
   alphaCSR[ 213 ][ 239 ],
   alphaCSR[ 213 ][ 240 ],
   alphaCSR[ 213 ][ 241 ],
   alphaCSR[ 213 ][ 242 ],
   alphaCSR[ 213 ][ 243 ],
   alphaCSR[ 213 ][ 244 ],
   alphaCSR[ 213 ][ 245 ],
   alphaCSR[ 213 ][ 246 ],
   alphaCSR[ 213 ][ 247 ],
   alphaCSR[ 213 ][ 248 ],
   alphaCSR[ 213 ][ 249 ],
   alphaCSR[ 213 ][ 250 ],
   alphaCSR[ 213 ][ 251 ],
   alphaCSR[ 213 ][ 252 ],
   alphaCSR[ 213 ][ 253 ],
   alphaCSR[ 213 ][ 254 ],
   alphaCSR[ 213 ][ 255 ],
   alphaCSR[ 213 ][ 256 ],
   alphaCSR[ 213 ][ 257 ],
   alphaCSR[ 213 ][ 258 ],
   alphaCSR[ 213 ][ 259 ],
   alphaCSR[ 213 ][ 260 ],
   alphaCSR[ 213 ][ 261 ],
   alphaCSR[ 213 ][ 262 ],
   alphaCSR[ 213 ][ 263 ],
   alphaCSR[ 213 ][ 264 ],
   alphaCSR[ 213 ][ 265 ],
   alphaCSR[ 213 ][ 266 ],
   alphaCSR[ 213 ][ 267 ],
   alphaCSR[ 213 ][ 268 ],
   alphaCSR[ 213 ][ 269 ],
   alphaCSR[ 213 ][ 270 ],
   alphaCSR[ 213 ][ 271 ],
   alphaCSR[ 213 ][ 272 ],
   alphaCSR[ 213 ][ 273 ],
   alphaCSR[ 213 ][ 274 ],
   alphaCSR[ 213 ][ 275 ],
   alphaCSR[ 213 ][ 276 ],
   alphaCSR[ 213 ][ 277 ],
   alphaCSR[ 213 ][ 278 ],
   alphaCSR[ 213 ][ 279 ],
   alphaCSR[ 213 ][ 280 ],
   alphaCSR[ 213 ][ 281 ],
   alphaCSR[ 213 ][ 282 ],
   alphaCSR[ 213 ][ 283 ],
   alphaCSR[ 213 ][ 284 ],
   alphaCSR[ 213 ][ 285 ],
   alphaCSR[ 213 ][ 286 ],
   alphaCSR[ 213 ][ 287 ],
   alphaCSR[ 213 ][ 288 ],
   alphaCSR[ 213 ][ 289 ],
   alphaCSR[ 213 ][ 290 ],
   alphaCSR[ 213 ][ 291 ],
   alphaCSR[ 213 ][ 292 ],
   alphaCSR[ 213 ][ 293 ],
   alphaCSR[ 213 ][ 294 ],
   alphaCSR[ 213 ][ 295 ],
   alphaCSR[ 213 ][ 296 ],
   alphaCSR[ 213 ][ 297 ],
   alphaCSR[ 213 ][ 298 ],
   alphaCSR[ 213 ][ 299 ],
   alphaCSR[ 213 ][ 300 ],
   alphaCSR[ 213 ][ 301 ],
   alphaCSR[ 213 ][ 302 ],
   alphaCSR[ 213 ][ 303 ],
   alphaCSR[ 213 ][ 304 ],
   alphaCSR[ 213 ][ 305 ],
   alphaCSR[ 213 ][ 306 ],
   alphaCSR[ 213 ][ 307 ],
   alphaCSR[ 213 ][ 308 ],
   alphaCSR[ 213 ][ 309 ],
   alphaCSR[ 213 ][ 310 ],
   alphaCSR[ 213 ][ 311 ],
   alphaCSR[ 213 ][ 312 ],
   alphaCSR[ 213 ][ 313 ],
   alphaCSR[ 213 ][ 314 ],
   alphaCSR[ 213 ][ 315 ],
   alphaCSR[ 213 ][ 316 ],
   alphaCSR[ 213 ][ 317 ],
   alphaCSR[ 213 ][ 318 ],
   alphaCSR[ 213 ][ 319 ],
   alphaCSR[ 213 ][ 320 ],
   alphaCSR[ 213 ][ 321 ],
   alphaCSR[ 213 ][ 322 ],
   alphaCSR[ 213 ][ 323 ],
   alphaCSR[ 213 ][ 324 ],
   alphaCSR[ 213 ][ 325 ],
   alphaCSR[ 213 ][ 326 ],
   alphaCSR[ 213 ][ 327 ],
   alphaCSR[ 213 ][ 328 ],
   alphaCSR[ 213 ][ 329 ],
   alphaCSR[ 213 ][ 330 ],
   alphaCSR[ 213 ][ 331 ],
   alphaCSR[ 213 ][ 332 ],
   alphaCSR[ 213 ][ 333 ],
   alphaCSR[ 213 ][ 334 ],
   alphaCSR[ 213 ][ 335 ],
   alphaCSR[ 213 ][ 336 ],
   alphaCSR[ 213 ][ 337 ],
   alphaCSR[ 213 ][ 338 ],
   alphaCSR[ 213 ][ 339 ],
   alphaCSR[ 213 ][ 340 ],
   alphaCSR[ 213 ][ 341 ],
   alphaCSR[ 213 ][ 342 ],
   alphaCSR[ 213 ][ 343 ],
   alphaCSR[ 213 ][ 344 ],
   alphaCSR[ 213 ][ 345 ],
   alphaCSR[ 213 ][ 346 ],
   alphaCSR[ 213 ][ 347 ],
   alphaCSR[ 213 ][ 348 ],
   alphaCSR[ 213 ][ 349 ],
   alphaCSR[ 213 ][ 350 ],
   alphaCSR[ 213 ][ 351 ],
   alphaCSR[ 213 ][ 352 ],
   alphaCSR[ 213 ][ 353 ],
   alphaCSR[ 213 ][ 354 ],
   alphaCSR[ 213 ][ 355 ],
   alphaCSR[ 213 ][ 356 ],
   alphaCSR[ 213 ][ 357 ],
   alphaCSR[ 213 ][ 358 ],
   alphaCSR[ 213 ][ 359 ],
   alphaCSR[ 213 ][ 360 ],
   alphaCSR[ 213 ][ 361 ],
   alphaCSR[ 213 ][ 362 ],
   alphaCSR[ 213 ][ 363 ],
   alphaCSR[ 213 ][ 364 ],
   alphaCSR[ 213 ][ 365 ],
   alphaCSR[ 213 ][ 366 ],
   alphaCSR[ 213 ][ 367 ],
   alphaCSR[ 213 ][ 368 ],
   alphaCSR[ 213 ][ 369 ],
   alphaCSR[ 213 ][ 370 ],
   alphaCSR[ 213 ][ 371 ],
   alphaCSR[ 213 ][ 372 ],
   alphaCSR[ 213 ][ 373 ],
   alphaCSR[ 213 ][ 374 ],
   alphaCSR[ 213 ][ 375 ],
   alphaCSR[ 213 ][ 376 ],
   alphaCSR[ 213 ][ 377 ],
   alphaCSR[ 213 ][ 378 ],
   alphaCSR[ 213 ][ 379 ],
   alphaCSR[ 213 ][ 380 ],
   alphaCSR[ 213 ][ 381 ],
   alphaCSR[ 213 ][ 382 ],
   alphaCSR[ 213 ][ 383 ],
   alphaCSR[ 214 ][ 0 ],
   alphaCSR[ 214 ][ 1 ],
   alphaCSR[ 214 ][ 2 ],
   alphaCSR[ 214 ][ 3 ],
   alphaCSR[ 214 ][ 4 ],
   alphaCSR[ 214 ][ 5 ],
   alphaCSR[ 214 ][ 6 ],
   alphaCSR[ 214 ][ 7 ],
   alphaCSR[ 214 ][ 8 ],
   alphaCSR[ 214 ][ 9 ],
   alphaCSR[ 214 ][ 10 ],
   alphaCSR[ 214 ][ 11 ],
   alphaCSR[ 214 ][ 12 ],
   alphaCSR[ 214 ][ 13 ],
   alphaCSR[ 214 ][ 14 ],
   alphaCSR[ 214 ][ 15 ],
   alphaCSR[ 214 ][ 16 ],
   alphaCSR[ 214 ][ 17 ],
   alphaCSR[ 214 ][ 18 ],
   alphaCSR[ 214 ][ 19 ],
   alphaCSR[ 214 ][ 20 ],
   alphaCSR[ 214 ][ 21 ],
   alphaCSR[ 214 ][ 22 ],
   alphaCSR[ 214 ][ 23 ],
   alphaCSR[ 214 ][ 24 ],
   alphaCSR[ 214 ][ 25 ],
   alphaCSR[ 214 ][ 26 ],
   alphaCSR[ 214 ][ 27 ],
   alphaCSR[ 214 ][ 28 ],
   alphaCSR[ 214 ][ 29 ],
   alphaCSR[ 214 ][ 30 ],
   alphaCSR[ 214 ][ 31 ],
   alphaCSR[ 214 ][ 32 ],
   alphaCSR[ 214 ][ 33 ],
   alphaCSR[ 214 ][ 34 ],
   alphaCSR[ 214 ][ 35 ],
   alphaCSR[ 214 ][ 36 ],
   alphaCSR[ 214 ][ 37 ],
   alphaCSR[ 214 ][ 38 ],
   alphaCSR[ 214 ][ 39 ],
   alphaCSR[ 214 ][ 40 ],
   alphaCSR[ 214 ][ 41 ],
   alphaCSR[ 214 ][ 42 ],
   alphaCSR[ 214 ][ 43 ],
   alphaCSR[ 214 ][ 44 ],
   alphaCSR[ 214 ][ 45 ],
   alphaCSR[ 214 ][ 46 ],
   alphaCSR[ 214 ][ 47 ],
   alphaCSR[ 214 ][ 48 ],
   alphaCSR[ 214 ][ 49 ],
   alphaCSR[ 214 ][ 50 ],
   alphaCSR[ 214 ][ 51 ],
   alphaCSR[ 214 ][ 52 ],
   alphaCSR[ 214 ][ 53 ],
   alphaCSR[ 214 ][ 54 ],
   alphaCSR[ 214 ][ 55 ],
   alphaCSR[ 214 ][ 56 ],
   alphaCSR[ 214 ][ 57 ],
   alphaCSR[ 214 ][ 58 ],
   alphaCSR[ 214 ][ 59 ],
   alphaCSR[ 214 ][ 60 ],
   alphaCSR[ 214 ][ 61 ],
   alphaCSR[ 214 ][ 62 ],
   alphaCSR[ 214 ][ 63 ],
   alphaCSR[ 214 ][ 64 ],
   alphaCSR[ 214 ][ 65 ],
   alphaCSR[ 214 ][ 66 ],
   alphaCSR[ 214 ][ 67 ],
   alphaCSR[ 214 ][ 68 ],
   alphaCSR[ 214 ][ 69 ],
   alphaCSR[ 214 ][ 70 ],
   alphaCSR[ 214 ][ 71 ],
   alphaCSR[ 214 ][ 72 ],
   alphaCSR[ 214 ][ 73 ],
   alphaCSR[ 214 ][ 74 ],
   alphaCSR[ 214 ][ 75 ],
   alphaCSR[ 214 ][ 76 ],
   alphaCSR[ 214 ][ 77 ],
   alphaCSR[ 214 ][ 78 ],
   alphaCSR[ 214 ][ 79 ],
   alphaCSR[ 214 ][ 80 ],
   alphaCSR[ 214 ][ 81 ],
   alphaCSR[ 214 ][ 82 ],
   alphaCSR[ 214 ][ 83 ],
   alphaCSR[ 214 ][ 84 ],
   alphaCSR[ 214 ][ 85 ],
   alphaCSR[ 214 ][ 86 ],
   alphaCSR[ 214 ][ 87 ],
   alphaCSR[ 214 ][ 88 ],
   alphaCSR[ 214 ][ 89 ],
   alphaCSR[ 214 ][ 90 ],
   alphaCSR[ 214 ][ 91 ],
   alphaCSR[ 214 ][ 92 ],
   alphaCSR[ 214 ][ 93 ],
   alphaCSR[ 214 ][ 94 ],
   alphaCSR[ 214 ][ 95 ],
   alphaCSR[ 214 ][ 96 ],
   alphaCSR[ 214 ][ 97 ],
   alphaCSR[ 214 ][ 98 ],
   alphaCSR[ 214 ][ 99 ],
   alphaCSR[ 214 ][ 100 ],
   alphaCSR[ 214 ][ 101 ],
   alphaCSR[ 214 ][ 102 ],
   alphaCSR[ 214 ][ 103 ],
   alphaCSR[ 214 ][ 104 ],
   alphaCSR[ 214 ][ 105 ],
   alphaCSR[ 214 ][ 106 ],
   alphaCSR[ 214 ][ 107 ],
   alphaCSR[ 214 ][ 108 ],
   alphaCSR[ 214 ][ 109 ],
   alphaCSR[ 214 ][ 110 ],
   alphaCSR[ 214 ][ 111 ],
   alphaCSR[ 214 ][ 112 ],
   alphaCSR[ 214 ][ 113 ],
   alphaCSR[ 214 ][ 114 ],
   alphaCSR[ 214 ][ 115 ],
   alphaCSR[ 214 ][ 116 ],
   alphaCSR[ 214 ][ 117 ],
   alphaCSR[ 214 ][ 118 ],
   alphaCSR[ 214 ][ 119 ],
   alphaCSR[ 214 ][ 120 ],
   alphaCSR[ 214 ][ 121 ],
   alphaCSR[ 214 ][ 122 ],
   alphaCSR[ 214 ][ 123 ],
   alphaCSR[ 214 ][ 124 ],
   alphaCSR[ 214 ][ 125 ],
   alphaCSR[ 214 ][ 126 ],
   alphaCSR[ 214 ][ 127 ],
   alphaCSR[ 214 ][ 128 ],
   alphaCSR[ 214 ][ 129 ],
   alphaCSR[ 214 ][ 130 ],
   alphaCSR[ 214 ][ 131 ],
   alphaCSR[ 214 ][ 132 ],
   alphaCSR[ 214 ][ 133 ],
   alphaCSR[ 214 ][ 134 ],
   alphaCSR[ 214 ][ 135 ],
   alphaCSR[ 214 ][ 136 ],
   alphaCSR[ 214 ][ 137 ],
   alphaCSR[ 214 ][ 138 ],
   alphaCSR[ 214 ][ 139 ],
   alphaCSR[ 214 ][ 140 ],
   alphaCSR[ 214 ][ 141 ],
   alphaCSR[ 214 ][ 142 ],
   alphaCSR[ 214 ][ 143 ],
   alphaCSR[ 214 ][ 144 ],
   alphaCSR[ 214 ][ 145 ],
   alphaCSR[ 214 ][ 146 ],
   alphaCSR[ 214 ][ 147 ],
   alphaCSR[ 214 ][ 148 ],
   alphaCSR[ 214 ][ 149 ],
   alphaCSR[ 214 ][ 150 ],
   alphaCSR[ 214 ][ 151 ],
   alphaCSR[ 214 ][ 152 ],
   alphaCSR[ 214 ][ 153 ],
   alphaCSR[ 214 ][ 154 ],
   alphaCSR[ 214 ][ 155 ],
   alphaCSR[ 214 ][ 156 ],
   alphaCSR[ 214 ][ 157 ],
   alphaCSR[ 214 ][ 158 ],
   alphaCSR[ 214 ][ 159 ],
   alphaCSR[ 214 ][ 160 ],
   alphaCSR[ 214 ][ 161 ],
   alphaCSR[ 214 ][ 162 ],
   alphaCSR[ 214 ][ 163 ],
   alphaCSR[ 214 ][ 164 ],
   alphaCSR[ 214 ][ 165 ],
   alphaCSR[ 214 ][ 166 ],
   alphaCSR[ 214 ][ 167 ],
   alphaCSR[ 214 ][ 168 ],
   alphaCSR[ 214 ][ 169 ],
   alphaCSR[ 214 ][ 170 ],
   alphaCSR[ 214 ][ 171 ],
   alphaCSR[ 214 ][ 172 ],
   alphaCSR[ 214 ][ 173 ],
   alphaCSR[ 214 ][ 174 ],
   alphaCSR[ 214 ][ 175 ],
   alphaCSR[ 214 ][ 176 ],
   alphaCSR[ 214 ][ 177 ],
   alphaCSR[ 214 ][ 178 ],
   alphaCSR[ 214 ][ 179 ],
   alphaCSR[ 214 ][ 180 ],
   alphaCSR[ 214 ][ 181 ],
   alphaCSR[ 214 ][ 182 ],
   alphaCSR[ 214 ][ 183 ],
   alphaCSR[ 214 ][ 184 ],
   alphaCSR[ 214 ][ 185 ],
   alphaCSR[ 214 ][ 186 ],
   alphaCSR[ 214 ][ 187 ],
   alphaCSR[ 214 ][ 188 ],
   alphaCSR[ 214 ][ 189 ],
   alphaCSR[ 214 ][ 190 ],
   alphaCSR[ 214 ][ 191 ],
   alphaCSR[ 214 ][ 192 ],
   alphaCSR[ 214 ][ 193 ],
   alphaCSR[ 214 ][ 194 ],
   alphaCSR[ 214 ][ 195 ],
   alphaCSR[ 214 ][ 196 ],
   alphaCSR[ 214 ][ 197 ],
   alphaCSR[ 214 ][ 198 ],
   alphaCSR[ 214 ][ 199 ],
   alphaCSR[ 214 ][ 200 ],
   alphaCSR[ 214 ][ 201 ],
   alphaCSR[ 214 ][ 202 ],
   alphaCSR[ 214 ][ 203 ],
   alphaCSR[ 214 ][ 204 ],
   alphaCSR[ 214 ][ 205 ],
   alphaCSR[ 214 ][ 206 ],
   alphaCSR[ 214 ][ 207 ],
   alphaCSR[ 214 ][ 208 ],
   alphaCSR[ 214 ][ 209 ],
   alphaCSR[ 214 ][ 210 ],
   alphaCSR[ 214 ][ 211 ],
   alphaCSR[ 214 ][ 212 ],
   alphaCSR[ 214 ][ 213 ],
   alphaCSR[ 214 ][ 214 ],
   alphaCSR[ 214 ][ 215 ],
   alphaCSR[ 214 ][ 216 ],
   alphaCSR[ 214 ][ 217 ],
   alphaCSR[ 214 ][ 218 ],
   alphaCSR[ 214 ][ 219 ],
   alphaCSR[ 214 ][ 220 ],
   alphaCSR[ 214 ][ 221 ],
   alphaCSR[ 214 ][ 222 ],
   alphaCSR[ 214 ][ 223 ],
   alphaCSR[ 214 ][ 224 ],
   alphaCSR[ 214 ][ 225 ],
   alphaCSR[ 214 ][ 226 ],
   alphaCSR[ 214 ][ 227 ],
   alphaCSR[ 214 ][ 228 ],
   alphaCSR[ 214 ][ 229 ],
   alphaCSR[ 214 ][ 230 ],
   alphaCSR[ 214 ][ 231 ],
   alphaCSR[ 214 ][ 232 ],
   alphaCSR[ 214 ][ 233 ],
   alphaCSR[ 214 ][ 234 ],
   alphaCSR[ 214 ][ 235 ],
   alphaCSR[ 214 ][ 236 ],
   alphaCSR[ 214 ][ 237 ],
   alphaCSR[ 214 ][ 238 ],
   alphaCSR[ 214 ][ 239 ],
   alphaCSR[ 214 ][ 240 ],
   alphaCSR[ 214 ][ 241 ],
   alphaCSR[ 214 ][ 242 ],
   alphaCSR[ 214 ][ 243 ],
   alphaCSR[ 214 ][ 244 ],
   alphaCSR[ 214 ][ 245 ],
   alphaCSR[ 214 ][ 246 ],
   alphaCSR[ 214 ][ 247 ],
   alphaCSR[ 214 ][ 248 ],
   alphaCSR[ 214 ][ 249 ],
   alphaCSR[ 214 ][ 250 ],
   alphaCSR[ 214 ][ 251 ],
   alphaCSR[ 214 ][ 252 ],
   alphaCSR[ 214 ][ 253 ],
   alphaCSR[ 214 ][ 254 ],
   alphaCSR[ 214 ][ 255 ],
   alphaCSR[ 214 ][ 256 ],
   alphaCSR[ 214 ][ 257 ],
   alphaCSR[ 214 ][ 258 ],
   alphaCSR[ 214 ][ 259 ],
   alphaCSR[ 214 ][ 260 ],
   alphaCSR[ 214 ][ 261 ],
   alphaCSR[ 214 ][ 262 ],
   alphaCSR[ 214 ][ 263 ],
   alphaCSR[ 214 ][ 264 ],
   alphaCSR[ 214 ][ 265 ],
   alphaCSR[ 214 ][ 266 ],
   alphaCSR[ 214 ][ 267 ],
   alphaCSR[ 214 ][ 268 ],
   alphaCSR[ 214 ][ 269 ],
   alphaCSR[ 214 ][ 270 ],
   alphaCSR[ 214 ][ 271 ],
   alphaCSR[ 214 ][ 272 ],
   alphaCSR[ 214 ][ 273 ],
   alphaCSR[ 214 ][ 274 ],
   alphaCSR[ 214 ][ 275 ],
   alphaCSR[ 214 ][ 276 ],
   alphaCSR[ 214 ][ 277 ],
   alphaCSR[ 214 ][ 278 ],
   alphaCSR[ 214 ][ 279 ],
   alphaCSR[ 214 ][ 280 ],
   alphaCSR[ 214 ][ 281 ],
   alphaCSR[ 214 ][ 282 ],
   alphaCSR[ 214 ][ 283 ],
   alphaCSR[ 214 ][ 284 ],
   alphaCSR[ 214 ][ 285 ],
   alphaCSR[ 214 ][ 286 ],
   alphaCSR[ 214 ][ 287 ],
   alphaCSR[ 214 ][ 288 ],
   alphaCSR[ 214 ][ 289 ],
   alphaCSR[ 214 ][ 290 ],
   alphaCSR[ 214 ][ 291 ],
   alphaCSR[ 214 ][ 292 ],
   alphaCSR[ 214 ][ 293 ],
   alphaCSR[ 214 ][ 294 ],
   alphaCSR[ 214 ][ 295 ],
   alphaCSR[ 214 ][ 296 ],
   alphaCSR[ 214 ][ 297 ],
   alphaCSR[ 214 ][ 298 ],
   alphaCSR[ 214 ][ 299 ],
   alphaCSR[ 214 ][ 300 ],
   alphaCSR[ 214 ][ 301 ],
   alphaCSR[ 214 ][ 302 ],
   alphaCSR[ 214 ][ 303 ],
   alphaCSR[ 214 ][ 304 ],
   alphaCSR[ 214 ][ 305 ],
   alphaCSR[ 214 ][ 306 ],
   alphaCSR[ 214 ][ 307 ],
   alphaCSR[ 214 ][ 308 ],
   alphaCSR[ 214 ][ 309 ],
   alphaCSR[ 214 ][ 310 ],
   alphaCSR[ 214 ][ 311 ],
   alphaCSR[ 214 ][ 312 ],
   alphaCSR[ 214 ][ 313 ],
   alphaCSR[ 214 ][ 314 ],
   alphaCSR[ 214 ][ 315 ],
   alphaCSR[ 214 ][ 316 ],
   alphaCSR[ 214 ][ 317 ],
   alphaCSR[ 214 ][ 318 ],
   alphaCSR[ 214 ][ 319 ],
   alphaCSR[ 214 ][ 320 ],
   alphaCSR[ 214 ][ 321 ],
   alphaCSR[ 214 ][ 322 ],
   alphaCSR[ 214 ][ 323 ],
   alphaCSR[ 214 ][ 324 ],
   alphaCSR[ 214 ][ 325 ],
   alphaCSR[ 214 ][ 326 ],
   alphaCSR[ 214 ][ 327 ],
   alphaCSR[ 214 ][ 328 ],
   alphaCSR[ 214 ][ 329 ],
   alphaCSR[ 214 ][ 330 ],
   alphaCSR[ 214 ][ 331 ],
   alphaCSR[ 214 ][ 332 ],
   alphaCSR[ 214 ][ 333 ],
   alphaCSR[ 214 ][ 334 ],
   alphaCSR[ 214 ][ 335 ],
   alphaCSR[ 214 ][ 336 ],
   alphaCSR[ 214 ][ 337 ],
   alphaCSR[ 214 ][ 338 ],
   alphaCSR[ 214 ][ 339 ],
   alphaCSR[ 214 ][ 340 ],
   alphaCSR[ 214 ][ 341 ],
   alphaCSR[ 214 ][ 342 ],
   alphaCSR[ 214 ][ 343 ],
   alphaCSR[ 214 ][ 344 ],
   alphaCSR[ 214 ][ 345 ],
   alphaCSR[ 214 ][ 346 ],
   alphaCSR[ 214 ][ 347 ],
   alphaCSR[ 214 ][ 348 ],
   alphaCSR[ 214 ][ 349 ],
   alphaCSR[ 214 ][ 350 ],
   alphaCSR[ 214 ][ 351 ],
   alphaCSR[ 214 ][ 352 ],
   alphaCSR[ 214 ][ 353 ],
   alphaCSR[ 214 ][ 354 ],
   alphaCSR[ 214 ][ 355 ],
   alphaCSR[ 214 ][ 356 ],
   alphaCSR[ 214 ][ 357 ],
   alphaCSR[ 214 ][ 358 ],
   alphaCSR[ 214 ][ 359 ],
   alphaCSR[ 214 ][ 360 ],
   alphaCSR[ 214 ][ 361 ],
   alphaCSR[ 214 ][ 362 ],
   alphaCSR[ 214 ][ 363 ],
   alphaCSR[ 214 ][ 364 ],
   alphaCSR[ 214 ][ 365 ],
   alphaCSR[ 214 ][ 366 ],
   alphaCSR[ 214 ][ 367 ],
   alphaCSR[ 214 ][ 368 ],
   alphaCSR[ 214 ][ 369 ],
   alphaCSR[ 214 ][ 370 ],
   alphaCSR[ 214 ][ 371 ],
   alphaCSR[ 214 ][ 372 ],
   alphaCSR[ 214 ][ 373 ],
   alphaCSR[ 214 ][ 374 ],
   alphaCSR[ 214 ][ 375 ],
   alphaCSR[ 214 ][ 376 ],
   alphaCSR[ 214 ][ 377 ],
   alphaCSR[ 214 ][ 378 ],
   alphaCSR[ 214 ][ 379 ],
   alphaCSR[ 214 ][ 380 ],
   alphaCSR[ 214 ][ 381 ],
   alphaCSR[ 214 ][ 382 ],
   alphaCSR[ 214 ][ 383 ],
   alphaCSR[ 215 ][ 0 ],
   alphaCSR[ 215 ][ 1 ],
   alphaCSR[ 215 ][ 2 ],
   alphaCSR[ 215 ][ 3 ],
   alphaCSR[ 215 ][ 4 ],
   alphaCSR[ 215 ][ 5 ],
   alphaCSR[ 215 ][ 6 ],
   alphaCSR[ 215 ][ 7 ],
   alphaCSR[ 215 ][ 8 ],
   alphaCSR[ 215 ][ 9 ],
   alphaCSR[ 215 ][ 10 ],
   alphaCSR[ 215 ][ 11 ],
   alphaCSR[ 215 ][ 12 ],
   alphaCSR[ 215 ][ 13 ],
   alphaCSR[ 215 ][ 14 ],
   alphaCSR[ 215 ][ 15 ],
   alphaCSR[ 215 ][ 16 ],
   alphaCSR[ 215 ][ 17 ],
   alphaCSR[ 215 ][ 18 ],
   alphaCSR[ 215 ][ 19 ],
   alphaCSR[ 215 ][ 20 ],
   alphaCSR[ 215 ][ 21 ],
   alphaCSR[ 215 ][ 22 ],
   alphaCSR[ 215 ][ 23 ],
   alphaCSR[ 215 ][ 24 ],
   alphaCSR[ 215 ][ 25 ],
   alphaCSR[ 215 ][ 26 ],
   alphaCSR[ 215 ][ 27 ],
   alphaCSR[ 215 ][ 28 ],
   alphaCSR[ 215 ][ 29 ],
   alphaCSR[ 215 ][ 30 ],
   alphaCSR[ 215 ][ 31 ],
   alphaCSR[ 215 ][ 32 ],
   alphaCSR[ 215 ][ 33 ],
   alphaCSR[ 215 ][ 34 ],
   alphaCSR[ 215 ][ 35 ],
   alphaCSR[ 215 ][ 36 ],
   alphaCSR[ 215 ][ 37 ],
   alphaCSR[ 215 ][ 38 ],
   alphaCSR[ 215 ][ 39 ],
   alphaCSR[ 215 ][ 40 ],
   alphaCSR[ 215 ][ 41 ],
   alphaCSR[ 215 ][ 42 ],
   alphaCSR[ 215 ][ 43 ],
   alphaCSR[ 215 ][ 44 ],
   alphaCSR[ 215 ][ 45 ],
   alphaCSR[ 215 ][ 46 ],
   alphaCSR[ 215 ][ 47 ],
   alphaCSR[ 215 ][ 48 ],
   alphaCSR[ 215 ][ 49 ],
   alphaCSR[ 215 ][ 50 ],
   alphaCSR[ 215 ][ 51 ],
   alphaCSR[ 215 ][ 52 ],
   alphaCSR[ 215 ][ 53 ],
   alphaCSR[ 215 ][ 54 ],
   alphaCSR[ 215 ][ 55 ],
   alphaCSR[ 215 ][ 56 ],
   alphaCSR[ 215 ][ 57 ],
   alphaCSR[ 215 ][ 58 ],
   alphaCSR[ 215 ][ 59 ],
   alphaCSR[ 215 ][ 60 ],
   alphaCSR[ 215 ][ 61 ],
   alphaCSR[ 215 ][ 62 ],
   alphaCSR[ 215 ][ 63 ],
   alphaCSR[ 215 ][ 64 ],
   alphaCSR[ 215 ][ 65 ],
   alphaCSR[ 215 ][ 66 ],
   alphaCSR[ 215 ][ 67 ],
   alphaCSR[ 215 ][ 68 ],
   alphaCSR[ 215 ][ 69 ],
   alphaCSR[ 215 ][ 70 ],
   alphaCSR[ 215 ][ 71 ],
   alphaCSR[ 215 ][ 72 ],
   alphaCSR[ 215 ][ 73 ],
   alphaCSR[ 215 ][ 74 ],
   alphaCSR[ 215 ][ 75 ],
   alphaCSR[ 215 ][ 76 ],
   alphaCSR[ 215 ][ 77 ],
   alphaCSR[ 215 ][ 78 ],
   alphaCSR[ 215 ][ 79 ],
   alphaCSR[ 215 ][ 80 ],
   alphaCSR[ 215 ][ 81 ],
   alphaCSR[ 215 ][ 82 ],
   alphaCSR[ 215 ][ 83 ],
   alphaCSR[ 215 ][ 84 ],
   alphaCSR[ 215 ][ 85 ],
   alphaCSR[ 215 ][ 86 ],
   alphaCSR[ 215 ][ 87 ],
   alphaCSR[ 215 ][ 88 ],
   alphaCSR[ 215 ][ 89 ],
   alphaCSR[ 215 ][ 90 ],
   alphaCSR[ 215 ][ 91 ],
   alphaCSR[ 215 ][ 92 ],
   alphaCSR[ 215 ][ 93 ],
   alphaCSR[ 215 ][ 94 ],
   alphaCSR[ 215 ][ 95 ],
   alphaCSR[ 215 ][ 96 ],
   alphaCSR[ 215 ][ 97 ],
   alphaCSR[ 215 ][ 98 ],
   alphaCSR[ 215 ][ 99 ],
   alphaCSR[ 215 ][ 100 ],
   alphaCSR[ 215 ][ 101 ],
   alphaCSR[ 215 ][ 102 ],
   alphaCSR[ 215 ][ 103 ],
   alphaCSR[ 215 ][ 104 ],
   alphaCSR[ 215 ][ 105 ],
   alphaCSR[ 215 ][ 106 ],
   alphaCSR[ 215 ][ 107 ],
   alphaCSR[ 215 ][ 108 ],
   alphaCSR[ 215 ][ 109 ],
   alphaCSR[ 215 ][ 110 ],
   alphaCSR[ 215 ][ 111 ],
   alphaCSR[ 215 ][ 112 ],
   alphaCSR[ 215 ][ 113 ],
   alphaCSR[ 215 ][ 114 ],
   alphaCSR[ 215 ][ 115 ],
   alphaCSR[ 215 ][ 116 ],
   alphaCSR[ 215 ][ 117 ],
   alphaCSR[ 215 ][ 118 ],
   alphaCSR[ 215 ][ 119 ],
   alphaCSR[ 215 ][ 120 ],
   alphaCSR[ 215 ][ 121 ],
   alphaCSR[ 215 ][ 122 ],
   alphaCSR[ 215 ][ 123 ],
   alphaCSR[ 215 ][ 124 ],
   alphaCSR[ 215 ][ 125 ],
   alphaCSR[ 215 ][ 126 ],
   alphaCSR[ 215 ][ 127 ],
   alphaCSR[ 215 ][ 128 ],
   alphaCSR[ 215 ][ 129 ],
   alphaCSR[ 215 ][ 130 ],
   alphaCSR[ 215 ][ 131 ],
   alphaCSR[ 215 ][ 132 ],
   alphaCSR[ 215 ][ 133 ],
   alphaCSR[ 215 ][ 134 ],
   alphaCSR[ 215 ][ 135 ],
   alphaCSR[ 215 ][ 136 ],
   alphaCSR[ 215 ][ 137 ],
   alphaCSR[ 215 ][ 138 ],
   alphaCSR[ 215 ][ 139 ],
   alphaCSR[ 215 ][ 140 ],
   alphaCSR[ 215 ][ 141 ],
   alphaCSR[ 215 ][ 142 ],
   alphaCSR[ 215 ][ 143 ],
   alphaCSR[ 215 ][ 144 ],
   alphaCSR[ 215 ][ 145 ],
   alphaCSR[ 215 ][ 146 ],
   alphaCSR[ 215 ][ 147 ],
   alphaCSR[ 215 ][ 148 ],
   alphaCSR[ 215 ][ 149 ],
   alphaCSR[ 215 ][ 150 ],
   alphaCSR[ 215 ][ 151 ],
   alphaCSR[ 215 ][ 152 ],
   alphaCSR[ 215 ][ 153 ],
   alphaCSR[ 215 ][ 154 ],
   alphaCSR[ 215 ][ 155 ],
   alphaCSR[ 215 ][ 156 ],
   alphaCSR[ 215 ][ 157 ],
   alphaCSR[ 215 ][ 158 ],
   alphaCSR[ 215 ][ 159 ],
   alphaCSR[ 215 ][ 160 ],
   alphaCSR[ 215 ][ 161 ],
   alphaCSR[ 215 ][ 162 ],
   alphaCSR[ 215 ][ 163 ],
   alphaCSR[ 215 ][ 164 ],
   alphaCSR[ 215 ][ 165 ],
   alphaCSR[ 215 ][ 166 ],
   alphaCSR[ 215 ][ 167 ],
   alphaCSR[ 215 ][ 168 ],
   alphaCSR[ 215 ][ 169 ],
   alphaCSR[ 215 ][ 170 ],
   alphaCSR[ 215 ][ 171 ],
   alphaCSR[ 215 ][ 172 ],
   alphaCSR[ 215 ][ 173 ],
   alphaCSR[ 215 ][ 174 ],
   alphaCSR[ 215 ][ 175 ],
   alphaCSR[ 215 ][ 176 ],
   alphaCSR[ 215 ][ 177 ],
   alphaCSR[ 215 ][ 178 ],
   alphaCSR[ 215 ][ 179 ],
   alphaCSR[ 215 ][ 180 ],
   alphaCSR[ 215 ][ 181 ],
   alphaCSR[ 215 ][ 182 ],
   alphaCSR[ 215 ][ 183 ],
   alphaCSR[ 215 ][ 184 ],
   alphaCSR[ 215 ][ 185 ],
   alphaCSR[ 215 ][ 186 ],
   alphaCSR[ 215 ][ 187 ],
   alphaCSR[ 215 ][ 188 ],
   alphaCSR[ 215 ][ 189 ],
   alphaCSR[ 215 ][ 190 ],
   alphaCSR[ 215 ][ 191 ],
   alphaCSR[ 215 ][ 192 ],
   alphaCSR[ 215 ][ 193 ],
   alphaCSR[ 215 ][ 194 ],
   alphaCSR[ 215 ][ 195 ],
   alphaCSR[ 215 ][ 196 ],
   alphaCSR[ 215 ][ 197 ],
   alphaCSR[ 215 ][ 198 ],
   alphaCSR[ 215 ][ 199 ],
   alphaCSR[ 215 ][ 200 ],
   alphaCSR[ 215 ][ 201 ],
   alphaCSR[ 215 ][ 202 ],
   alphaCSR[ 215 ][ 203 ],
   alphaCSR[ 215 ][ 204 ],
   alphaCSR[ 215 ][ 205 ],
   alphaCSR[ 215 ][ 206 ],
   alphaCSR[ 215 ][ 207 ],
   alphaCSR[ 215 ][ 208 ],
   alphaCSR[ 215 ][ 209 ],
   alphaCSR[ 215 ][ 210 ],
   alphaCSR[ 215 ][ 211 ],
   alphaCSR[ 215 ][ 212 ],
   alphaCSR[ 215 ][ 213 ],
   alphaCSR[ 215 ][ 214 ],
   alphaCSR[ 215 ][ 215 ],
   alphaCSR[ 215 ][ 216 ],
   alphaCSR[ 215 ][ 217 ],
   alphaCSR[ 215 ][ 218 ],
   alphaCSR[ 215 ][ 219 ],
   alphaCSR[ 215 ][ 220 ],
   alphaCSR[ 215 ][ 221 ],
   alphaCSR[ 215 ][ 222 ],
   alphaCSR[ 215 ][ 223 ],
   alphaCSR[ 215 ][ 224 ],
   alphaCSR[ 215 ][ 225 ],
   alphaCSR[ 215 ][ 226 ],
   alphaCSR[ 215 ][ 227 ],
   alphaCSR[ 215 ][ 228 ],
   alphaCSR[ 215 ][ 229 ],
   alphaCSR[ 215 ][ 230 ],
   alphaCSR[ 215 ][ 231 ],
   alphaCSR[ 215 ][ 232 ],
   alphaCSR[ 215 ][ 233 ],
   alphaCSR[ 215 ][ 234 ],
   alphaCSR[ 215 ][ 235 ],
   alphaCSR[ 215 ][ 236 ],
   alphaCSR[ 215 ][ 237 ],
   alphaCSR[ 215 ][ 238 ],
   alphaCSR[ 215 ][ 239 ],
   alphaCSR[ 215 ][ 240 ],
   alphaCSR[ 215 ][ 241 ],
   alphaCSR[ 215 ][ 242 ],
   alphaCSR[ 215 ][ 243 ],
   alphaCSR[ 215 ][ 244 ],
   alphaCSR[ 215 ][ 245 ],
   alphaCSR[ 215 ][ 246 ],
   alphaCSR[ 215 ][ 247 ],
   alphaCSR[ 215 ][ 248 ],
   alphaCSR[ 215 ][ 249 ],
   alphaCSR[ 215 ][ 250 ],
   alphaCSR[ 215 ][ 251 ],
   alphaCSR[ 215 ][ 252 ],
   alphaCSR[ 215 ][ 253 ],
   alphaCSR[ 215 ][ 254 ],
   alphaCSR[ 215 ][ 255 ],
   alphaCSR[ 215 ][ 256 ],
   alphaCSR[ 215 ][ 257 ],
   alphaCSR[ 215 ][ 258 ],
   alphaCSR[ 215 ][ 259 ],
   alphaCSR[ 215 ][ 260 ],
   alphaCSR[ 215 ][ 261 ],
   alphaCSR[ 215 ][ 262 ],
   alphaCSR[ 215 ][ 263 ],
   alphaCSR[ 215 ][ 264 ],
   alphaCSR[ 215 ][ 265 ],
   alphaCSR[ 215 ][ 266 ],
   alphaCSR[ 215 ][ 267 ],
   alphaCSR[ 215 ][ 268 ],
   alphaCSR[ 215 ][ 269 ],
   alphaCSR[ 215 ][ 270 ],
   alphaCSR[ 215 ][ 271 ],
   alphaCSR[ 215 ][ 272 ],
   alphaCSR[ 215 ][ 273 ],
   alphaCSR[ 215 ][ 274 ],
   alphaCSR[ 215 ][ 275 ],
   alphaCSR[ 215 ][ 276 ],
   alphaCSR[ 215 ][ 277 ],
   alphaCSR[ 215 ][ 278 ],
   alphaCSR[ 215 ][ 279 ],
   alphaCSR[ 215 ][ 280 ],
   alphaCSR[ 215 ][ 281 ],
   alphaCSR[ 215 ][ 282 ],
   alphaCSR[ 215 ][ 283 ],
   alphaCSR[ 215 ][ 284 ],
   alphaCSR[ 215 ][ 285 ],
   alphaCSR[ 215 ][ 286 ],
   alphaCSR[ 215 ][ 287 ],
   alphaCSR[ 215 ][ 288 ],
   alphaCSR[ 215 ][ 289 ],
   alphaCSR[ 215 ][ 290 ],
   alphaCSR[ 215 ][ 291 ],
   alphaCSR[ 215 ][ 292 ],
   alphaCSR[ 215 ][ 293 ],
   alphaCSR[ 215 ][ 294 ],
   alphaCSR[ 215 ][ 295 ],
   alphaCSR[ 215 ][ 296 ],
   alphaCSR[ 215 ][ 297 ],
   alphaCSR[ 215 ][ 298 ],
   alphaCSR[ 215 ][ 299 ],
   alphaCSR[ 215 ][ 300 ],
   alphaCSR[ 215 ][ 301 ],
   alphaCSR[ 215 ][ 302 ],
   alphaCSR[ 215 ][ 303 ],
   alphaCSR[ 215 ][ 304 ],
   alphaCSR[ 215 ][ 305 ],
   alphaCSR[ 215 ][ 306 ],
   alphaCSR[ 215 ][ 307 ],
   alphaCSR[ 215 ][ 308 ],
   alphaCSR[ 215 ][ 309 ],
   alphaCSR[ 215 ][ 310 ],
   alphaCSR[ 215 ][ 311 ],
   alphaCSR[ 215 ][ 312 ],
   alphaCSR[ 215 ][ 313 ],
   alphaCSR[ 215 ][ 314 ],
   alphaCSR[ 215 ][ 315 ],
   alphaCSR[ 215 ][ 316 ],
   alphaCSR[ 215 ][ 317 ],
   alphaCSR[ 215 ][ 318 ],
   alphaCSR[ 215 ][ 319 ],
   alphaCSR[ 215 ][ 320 ],
   alphaCSR[ 215 ][ 321 ],
   alphaCSR[ 215 ][ 322 ],
   alphaCSR[ 215 ][ 323 ],
   alphaCSR[ 215 ][ 324 ],
   alphaCSR[ 215 ][ 325 ],
   alphaCSR[ 215 ][ 326 ],
   alphaCSR[ 215 ][ 327 ],
   alphaCSR[ 215 ][ 328 ],
   alphaCSR[ 215 ][ 329 ],
   alphaCSR[ 215 ][ 330 ],
   alphaCSR[ 215 ][ 331 ],
   alphaCSR[ 215 ][ 332 ],
   alphaCSR[ 215 ][ 333 ],
   alphaCSR[ 215 ][ 334 ],
   alphaCSR[ 215 ][ 335 ],
   alphaCSR[ 215 ][ 336 ],
   alphaCSR[ 215 ][ 337 ],
   alphaCSR[ 215 ][ 338 ],
   alphaCSR[ 215 ][ 339 ],
   alphaCSR[ 215 ][ 340 ],
   alphaCSR[ 215 ][ 341 ],
   alphaCSR[ 215 ][ 342 ],
   alphaCSR[ 215 ][ 343 ],
   alphaCSR[ 215 ][ 344 ],
   alphaCSR[ 215 ][ 345 ],
   alphaCSR[ 215 ][ 346 ],
   alphaCSR[ 215 ][ 347 ],
   alphaCSR[ 215 ][ 348 ],
   alphaCSR[ 215 ][ 349 ],
   alphaCSR[ 215 ][ 350 ],
   alphaCSR[ 215 ][ 351 ],
   alphaCSR[ 215 ][ 352 ],
   alphaCSR[ 215 ][ 353 ],
   alphaCSR[ 215 ][ 354 ],
   alphaCSR[ 215 ][ 355 ],
   alphaCSR[ 215 ][ 356 ],
   alphaCSR[ 215 ][ 357 ],
   alphaCSR[ 215 ][ 358 ],
   alphaCSR[ 215 ][ 359 ],
   alphaCSR[ 215 ][ 360 ],
   alphaCSR[ 215 ][ 361 ],
   alphaCSR[ 215 ][ 362 ],
   alphaCSR[ 215 ][ 363 ],
   alphaCSR[ 215 ][ 364 ],
   alphaCSR[ 215 ][ 365 ],
   alphaCSR[ 215 ][ 366 ],
   alphaCSR[ 215 ][ 367 ],
   alphaCSR[ 215 ][ 368 ],
   alphaCSR[ 215 ][ 369 ],
   alphaCSR[ 215 ][ 370 ],
   alphaCSR[ 215 ][ 371 ],
   alphaCSR[ 215 ][ 372 ],
   alphaCSR[ 215 ][ 373 ],
   alphaCSR[ 215 ][ 374 ],
   alphaCSR[ 215 ][ 375 ],
   alphaCSR[ 215 ][ 376 ],
   alphaCSR[ 215 ][ 377 ],
   alphaCSR[ 215 ][ 378 ],
   alphaCSR[ 215 ][ 379 ],
   alphaCSR[ 215 ][ 380 ],
   alphaCSR[ 215 ][ 381 ],
   alphaCSR[ 215 ][ 382 ],
   alphaCSR[ 215 ][ 383 ],
   alphaCSR[ 216 ][ 0 ],
   alphaCSR[ 216 ][ 1 ],
   alphaCSR[ 216 ][ 2 ],
   alphaCSR[ 216 ][ 3 ],
   alphaCSR[ 216 ][ 4 ],
   alphaCSR[ 216 ][ 5 ],
   alphaCSR[ 216 ][ 6 ],
   alphaCSR[ 216 ][ 7 ],
   alphaCSR[ 216 ][ 8 ],
   alphaCSR[ 216 ][ 9 ],
   alphaCSR[ 216 ][ 10 ],
   alphaCSR[ 216 ][ 11 ],
   alphaCSR[ 216 ][ 12 ],
   alphaCSR[ 216 ][ 13 ],
   alphaCSR[ 216 ][ 14 ],
   alphaCSR[ 216 ][ 15 ],
   alphaCSR[ 216 ][ 16 ],
   alphaCSR[ 216 ][ 17 ],
   alphaCSR[ 216 ][ 18 ],
   alphaCSR[ 216 ][ 19 ],
   alphaCSR[ 216 ][ 20 ],
   alphaCSR[ 216 ][ 21 ],
   alphaCSR[ 216 ][ 22 ],
   alphaCSR[ 216 ][ 23 ],
   alphaCSR[ 216 ][ 24 ],
   alphaCSR[ 216 ][ 25 ],
   alphaCSR[ 216 ][ 26 ],
   alphaCSR[ 216 ][ 27 ],
   alphaCSR[ 216 ][ 28 ],
   alphaCSR[ 216 ][ 29 ],
   alphaCSR[ 216 ][ 30 ],
   alphaCSR[ 216 ][ 31 ],
   alphaCSR[ 216 ][ 32 ],
   alphaCSR[ 216 ][ 33 ],
   alphaCSR[ 216 ][ 34 ],
   alphaCSR[ 216 ][ 35 ],
   alphaCSR[ 216 ][ 36 ],
   alphaCSR[ 216 ][ 37 ],
   alphaCSR[ 216 ][ 38 ],
   alphaCSR[ 216 ][ 39 ],
   alphaCSR[ 216 ][ 40 ],
   alphaCSR[ 216 ][ 41 ],
   alphaCSR[ 216 ][ 42 ],
   alphaCSR[ 216 ][ 43 ],
   alphaCSR[ 216 ][ 44 ],
   alphaCSR[ 216 ][ 45 ],
   alphaCSR[ 216 ][ 46 ],
   alphaCSR[ 216 ][ 47 ],
   alphaCSR[ 216 ][ 48 ],
   alphaCSR[ 216 ][ 49 ],
   alphaCSR[ 216 ][ 50 ],
   alphaCSR[ 216 ][ 51 ],
   alphaCSR[ 216 ][ 52 ],
   alphaCSR[ 216 ][ 53 ],
   alphaCSR[ 216 ][ 54 ],
   alphaCSR[ 216 ][ 55 ],
   alphaCSR[ 216 ][ 56 ],
   alphaCSR[ 216 ][ 57 ],
   alphaCSR[ 216 ][ 58 ],
   alphaCSR[ 216 ][ 59 ],
   alphaCSR[ 216 ][ 60 ],
   alphaCSR[ 216 ][ 61 ],
   alphaCSR[ 216 ][ 62 ],
   alphaCSR[ 216 ][ 63 ],
   alphaCSR[ 216 ][ 64 ],
   alphaCSR[ 216 ][ 65 ],
   alphaCSR[ 216 ][ 66 ],
   alphaCSR[ 216 ][ 67 ],
   alphaCSR[ 216 ][ 68 ],
   alphaCSR[ 216 ][ 69 ],
   alphaCSR[ 216 ][ 70 ],
   alphaCSR[ 216 ][ 71 ],
   alphaCSR[ 216 ][ 72 ],
   alphaCSR[ 216 ][ 73 ],
   alphaCSR[ 216 ][ 74 ],
   alphaCSR[ 216 ][ 75 ],
   alphaCSR[ 216 ][ 76 ],
   alphaCSR[ 216 ][ 77 ],
   alphaCSR[ 216 ][ 78 ],
   alphaCSR[ 216 ][ 79 ],
   alphaCSR[ 216 ][ 80 ],
   alphaCSR[ 216 ][ 81 ],
   alphaCSR[ 216 ][ 82 ],
   alphaCSR[ 216 ][ 83 ],
   alphaCSR[ 216 ][ 84 ],
   alphaCSR[ 216 ][ 85 ],
   alphaCSR[ 216 ][ 86 ],
   alphaCSR[ 216 ][ 87 ],
   alphaCSR[ 216 ][ 88 ],
   alphaCSR[ 216 ][ 89 ],
   alphaCSR[ 216 ][ 90 ],
   alphaCSR[ 216 ][ 91 ],
   alphaCSR[ 216 ][ 92 ],
   alphaCSR[ 216 ][ 93 ],
   alphaCSR[ 216 ][ 94 ],
   alphaCSR[ 216 ][ 95 ],
   alphaCSR[ 216 ][ 96 ],
   alphaCSR[ 216 ][ 97 ],
   alphaCSR[ 216 ][ 98 ],
   alphaCSR[ 216 ][ 99 ],
   alphaCSR[ 216 ][ 100 ],
   alphaCSR[ 216 ][ 101 ],
   alphaCSR[ 216 ][ 102 ],
   alphaCSR[ 216 ][ 103 ],
   alphaCSR[ 216 ][ 104 ],
   alphaCSR[ 216 ][ 105 ],
   alphaCSR[ 216 ][ 106 ],
   alphaCSR[ 216 ][ 107 ],
   alphaCSR[ 216 ][ 108 ],
   alphaCSR[ 216 ][ 109 ],
   alphaCSR[ 216 ][ 110 ],
   alphaCSR[ 216 ][ 111 ],
   alphaCSR[ 216 ][ 112 ],
   alphaCSR[ 216 ][ 113 ],
   alphaCSR[ 216 ][ 114 ],
   alphaCSR[ 216 ][ 115 ],
   alphaCSR[ 216 ][ 116 ],
   alphaCSR[ 216 ][ 117 ],
   alphaCSR[ 216 ][ 118 ],
   alphaCSR[ 216 ][ 119 ],
   alphaCSR[ 216 ][ 120 ],
   alphaCSR[ 216 ][ 121 ],
   alphaCSR[ 216 ][ 122 ],
   alphaCSR[ 216 ][ 123 ],
   alphaCSR[ 216 ][ 124 ],
   alphaCSR[ 216 ][ 125 ],
   alphaCSR[ 216 ][ 126 ],
   alphaCSR[ 216 ][ 127 ],
   alphaCSR[ 216 ][ 128 ],
   alphaCSR[ 216 ][ 129 ],
   alphaCSR[ 216 ][ 130 ],
   alphaCSR[ 216 ][ 131 ],
   alphaCSR[ 216 ][ 132 ],
   alphaCSR[ 216 ][ 133 ],
   alphaCSR[ 216 ][ 134 ],
   alphaCSR[ 216 ][ 135 ],
   alphaCSR[ 216 ][ 136 ],
   alphaCSR[ 216 ][ 137 ],
   alphaCSR[ 216 ][ 138 ],
   alphaCSR[ 216 ][ 139 ],
   alphaCSR[ 216 ][ 140 ],
   alphaCSR[ 216 ][ 141 ],
   alphaCSR[ 216 ][ 142 ],
   alphaCSR[ 216 ][ 143 ],
   alphaCSR[ 216 ][ 144 ],
   alphaCSR[ 216 ][ 145 ],
   alphaCSR[ 216 ][ 146 ],
   alphaCSR[ 216 ][ 147 ],
   alphaCSR[ 216 ][ 148 ],
   alphaCSR[ 216 ][ 149 ],
   alphaCSR[ 216 ][ 150 ],
   alphaCSR[ 216 ][ 151 ],
   alphaCSR[ 216 ][ 152 ],
   alphaCSR[ 216 ][ 153 ],
   alphaCSR[ 216 ][ 154 ],
   alphaCSR[ 216 ][ 155 ],
   alphaCSR[ 216 ][ 156 ],
   alphaCSR[ 216 ][ 157 ],
   alphaCSR[ 216 ][ 158 ],
   alphaCSR[ 216 ][ 159 ],
   alphaCSR[ 216 ][ 160 ],
   alphaCSR[ 216 ][ 161 ],
   alphaCSR[ 216 ][ 162 ],
   alphaCSR[ 216 ][ 163 ],
   alphaCSR[ 216 ][ 164 ],
   alphaCSR[ 216 ][ 165 ],
   alphaCSR[ 216 ][ 166 ],
   alphaCSR[ 216 ][ 167 ],
   alphaCSR[ 216 ][ 168 ],
   alphaCSR[ 216 ][ 169 ],
   alphaCSR[ 216 ][ 170 ],
   alphaCSR[ 216 ][ 171 ],
   alphaCSR[ 216 ][ 172 ],
   alphaCSR[ 216 ][ 173 ],
   alphaCSR[ 216 ][ 174 ],
   alphaCSR[ 216 ][ 175 ],
   alphaCSR[ 216 ][ 176 ],
   alphaCSR[ 216 ][ 177 ],
   alphaCSR[ 216 ][ 178 ],
   alphaCSR[ 216 ][ 179 ],
   alphaCSR[ 216 ][ 180 ],
   alphaCSR[ 216 ][ 181 ],
   alphaCSR[ 216 ][ 182 ],
   alphaCSR[ 216 ][ 183 ],
   alphaCSR[ 216 ][ 184 ],
   alphaCSR[ 216 ][ 185 ],
   alphaCSR[ 216 ][ 186 ],
   alphaCSR[ 216 ][ 187 ],
   alphaCSR[ 216 ][ 188 ],
   alphaCSR[ 216 ][ 189 ],
   alphaCSR[ 216 ][ 190 ],
   alphaCSR[ 216 ][ 191 ],
   alphaCSR[ 216 ][ 192 ],
   alphaCSR[ 216 ][ 193 ],
   alphaCSR[ 216 ][ 194 ],
   alphaCSR[ 216 ][ 195 ],
   alphaCSR[ 216 ][ 196 ],
   alphaCSR[ 216 ][ 197 ],
   alphaCSR[ 216 ][ 198 ],
   alphaCSR[ 216 ][ 199 ],
   alphaCSR[ 216 ][ 200 ],
   alphaCSR[ 216 ][ 201 ],
   alphaCSR[ 216 ][ 202 ],
   alphaCSR[ 216 ][ 203 ],
   alphaCSR[ 216 ][ 204 ],
   alphaCSR[ 216 ][ 205 ],
   alphaCSR[ 216 ][ 206 ],
   alphaCSR[ 216 ][ 207 ],
   alphaCSR[ 216 ][ 208 ],
   alphaCSR[ 216 ][ 209 ],
   alphaCSR[ 216 ][ 210 ],
   alphaCSR[ 216 ][ 211 ],
   alphaCSR[ 216 ][ 212 ],
   alphaCSR[ 216 ][ 213 ],
   alphaCSR[ 216 ][ 214 ],
   alphaCSR[ 216 ][ 215 ],
   alphaCSR[ 216 ][ 216 ],
   alphaCSR[ 216 ][ 217 ],
   alphaCSR[ 216 ][ 218 ],
   alphaCSR[ 216 ][ 219 ],
   alphaCSR[ 216 ][ 220 ],
   alphaCSR[ 216 ][ 221 ],
   alphaCSR[ 216 ][ 222 ],
   alphaCSR[ 216 ][ 223 ],
   alphaCSR[ 216 ][ 224 ],
   alphaCSR[ 216 ][ 225 ],
   alphaCSR[ 216 ][ 226 ],
   alphaCSR[ 216 ][ 227 ],
   alphaCSR[ 216 ][ 228 ],
   alphaCSR[ 216 ][ 229 ],
   alphaCSR[ 216 ][ 230 ],
   alphaCSR[ 216 ][ 231 ],
   alphaCSR[ 216 ][ 232 ],
   alphaCSR[ 216 ][ 233 ],
   alphaCSR[ 216 ][ 234 ],
   alphaCSR[ 216 ][ 235 ],
   alphaCSR[ 216 ][ 236 ],
   alphaCSR[ 216 ][ 237 ],
   alphaCSR[ 216 ][ 238 ],
   alphaCSR[ 216 ][ 239 ],
   alphaCSR[ 216 ][ 240 ],
   alphaCSR[ 216 ][ 241 ],
   alphaCSR[ 216 ][ 242 ],
   alphaCSR[ 216 ][ 243 ],
   alphaCSR[ 216 ][ 244 ],
   alphaCSR[ 216 ][ 245 ],
   alphaCSR[ 216 ][ 246 ],
   alphaCSR[ 216 ][ 247 ],
   alphaCSR[ 216 ][ 248 ],
   alphaCSR[ 216 ][ 249 ],
   alphaCSR[ 216 ][ 250 ],
   alphaCSR[ 216 ][ 251 ],
   alphaCSR[ 216 ][ 252 ],
   alphaCSR[ 216 ][ 253 ],
   alphaCSR[ 216 ][ 254 ],
   alphaCSR[ 216 ][ 255 ],
   alphaCSR[ 216 ][ 256 ],
   alphaCSR[ 216 ][ 257 ],
   alphaCSR[ 216 ][ 258 ],
   alphaCSR[ 216 ][ 259 ],
   alphaCSR[ 216 ][ 260 ],
   alphaCSR[ 216 ][ 261 ],
   alphaCSR[ 216 ][ 262 ],
   alphaCSR[ 216 ][ 263 ],
   alphaCSR[ 216 ][ 264 ],
   alphaCSR[ 216 ][ 265 ],
   alphaCSR[ 216 ][ 266 ],
   alphaCSR[ 216 ][ 267 ],
   alphaCSR[ 216 ][ 268 ],
   alphaCSR[ 216 ][ 269 ],
   alphaCSR[ 216 ][ 270 ],
   alphaCSR[ 216 ][ 271 ],
   alphaCSR[ 216 ][ 272 ],
   alphaCSR[ 216 ][ 273 ],
   alphaCSR[ 216 ][ 274 ],
   alphaCSR[ 216 ][ 275 ],
   alphaCSR[ 216 ][ 276 ],
   alphaCSR[ 216 ][ 277 ],
   alphaCSR[ 216 ][ 278 ],
   alphaCSR[ 216 ][ 279 ],
   alphaCSR[ 216 ][ 280 ],
   alphaCSR[ 216 ][ 281 ],
   alphaCSR[ 216 ][ 282 ],
   alphaCSR[ 216 ][ 283 ],
   alphaCSR[ 216 ][ 284 ],
   alphaCSR[ 216 ][ 285 ],
   alphaCSR[ 216 ][ 286 ],
   alphaCSR[ 216 ][ 287 ],
   alphaCSR[ 216 ][ 288 ],
   alphaCSR[ 216 ][ 289 ],
   alphaCSR[ 216 ][ 290 ],
   alphaCSR[ 216 ][ 291 ],
   alphaCSR[ 216 ][ 292 ],
   alphaCSR[ 216 ][ 293 ],
   alphaCSR[ 216 ][ 294 ],
   alphaCSR[ 216 ][ 295 ],
   alphaCSR[ 216 ][ 296 ],
   alphaCSR[ 216 ][ 297 ],
   alphaCSR[ 216 ][ 298 ],
   alphaCSR[ 216 ][ 299 ],
   alphaCSR[ 216 ][ 300 ],
   alphaCSR[ 216 ][ 301 ],
   alphaCSR[ 216 ][ 302 ],
   alphaCSR[ 216 ][ 303 ],
   alphaCSR[ 216 ][ 304 ],
   alphaCSR[ 216 ][ 305 ],
   alphaCSR[ 216 ][ 306 ],
   alphaCSR[ 216 ][ 307 ],
   alphaCSR[ 216 ][ 308 ],
   alphaCSR[ 216 ][ 309 ],
   alphaCSR[ 216 ][ 310 ],
   alphaCSR[ 216 ][ 311 ],
   alphaCSR[ 216 ][ 312 ],
   alphaCSR[ 216 ][ 313 ],
   alphaCSR[ 216 ][ 314 ],
   alphaCSR[ 216 ][ 315 ],
   alphaCSR[ 216 ][ 316 ],
   alphaCSR[ 216 ][ 317 ],
   alphaCSR[ 216 ][ 318 ],
   alphaCSR[ 216 ][ 319 ],
   alphaCSR[ 216 ][ 320 ],
   alphaCSR[ 216 ][ 321 ],
   alphaCSR[ 216 ][ 322 ],
   alphaCSR[ 216 ][ 323 ],
   alphaCSR[ 216 ][ 324 ],
   alphaCSR[ 216 ][ 325 ],
   alphaCSR[ 216 ][ 326 ],
   alphaCSR[ 216 ][ 327 ],
   alphaCSR[ 216 ][ 328 ],
   alphaCSR[ 216 ][ 329 ],
   alphaCSR[ 216 ][ 330 ],
   alphaCSR[ 216 ][ 331 ],
   alphaCSR[ 216 ][ 332 ],
   alphaCSR[ 216 ][ 333 ],
   alphaCSR[ 216 ][ 334 ],
   alphaCSR[ 216 ][ 335 ],
   alphaCSR[ 216 ][ 336 ],
   alphaCSR[ 216 ][ 337 ],
   alphaCSR[ 216 ][ 338 ],
   alphaCSR[ 216 ][ 339 ],
   alphaCSR[ 216 ][ 340 ],
   alphaCSR[ 216 ][ 341 ],
   alphaCSR[ 216 ][ 342 ],
   alphaCSR[ 216 ][ 343 ],
   alphaCSR[ 216 ][ 344 ],
   alphaCSR[ 216 ][ 345 ],
   alphaCSR[ 216 ][ 346 ],
   alphaCSR[ 216 ][ 347 ],
   alphaCSR[ 216 ][ 348 ],
   alphaCSR[ 216 ][ 349 ],
   alphaCSR[ 216 ][ 350 ],
   alphaCSR[ 216 ][ 351 ],
   alphaCSR[ 216 ][ 352 ],
   alphaCSR[ 216 ][ 353 ],
   alphaCSR[ 216 ][ 354 ],
   alphaCSR[ 216 ][ 355 ],
   alphaCSR[ 216 ][ 356 ],
   alphaCSR[ 216 ][ 357 ],
   alphaCSR[ 216 ][ 358 ],
   alphaCSR[ 216 ][ 359 ],
   alphaCSR[ 216 ][ 360 ],
   alphaCSR[ 216 ][ 361 ],
   alphaCSR[ 216 ][ 362 ],
   alphaCSR[ 216 ][ 363 ],
   alphaCSR[ 216 ][ 364 ],
   alphaCSR[ 216 ][ 365 ],
   alphaCSR[ 216 ][ 366 ],
   alphaCSR[ 216 ][ 367 ],
   alphaCSR[ 216 ][ 368 ],
   alphaCSR[ 216 ][ 369 ],
   alphaCSR[ 216 ][ 370 ],
   alphaCSR[ 216 ][ 371 ],
   alphaCSR[ 216 ][ 372 ],
   alphaCSR[ 216 ][ 373 ],
   alphaCSR[ 216 ][ 374 ],
   alphaCSR[ 216 ][ 375 ],
   alphaCSR[ 216 ][ 376 ],
   alphaCSR[ 216 ][ 377 ],
   alphaCSR[ 216 ][ 378 ],
   alphaCSR[ 216 ][ 379 ],
   alphaCSR[ 216 ][ 380 ],
   alphaCSR[ 216 ][ 381 ],
   alphaCSR[ 216 ][ 382 ],
   alphaCSR[ 216 ][ 383 ],
   alphaCSR[ 217 ][ 0 ],
   alphaCSR[ 217 ][ 1 ],
   alphaCSR[ 217 ][ 2 ],
   alphaCSR[ 217 ][ 3 ],
   alphaCSR[ 217 ][ 4 ],
   alphaCSR[ 217 ][ 5 ],
   alphaCSR[ 217 ][ 6 ],
   alphaCSR[ 217 ][ 7 ],
   alphaCSR[ 217 ][ 8 ],
   alphaCSR[ 217 ][ 9 ],
   alphaCSR[ 217 ][ 10 ],
   alphaCSR[ 217 ][ 11 ],
   alphaCSR[ 217 ][ 12 ],
   alphaCSR[ 217 ][ 13 ],
   alphaCSR[ 217 ][ 14 ],
   alphaCSR[ 217 ][ 15 ],
   alphaCSR[ 217 ][ 16 ],
   alphaCSR[ 217 ][ 17 ],
   alphaCSR[ 217 ][ 18 ],
   alphaCSR[ 217 ][ 19 ],
   alphaCSR[ 217 ][ 20 ],
   alphaCSR[ 217 ][ 21 ],
   alphaCSR[ 217 ][ 22 ],
   alphaCSR[ 217 ][ 23 ],
   alphaCSR[ 217 ][ 24 ],
   alphaCSR[ 217 ][ 25 ],
   alphaCSR[ 217 ][ 26 ],
   alphaCSR[ 217 ][ 27 ],
   alphaCSR[ 217 ][ 28 ],
   alphaCSR[ 217 ][ 29 ],
   alphaCSR[ 217 ][ 30 ],
   alphaCSR[ 217 ][ 31 ],
   alphaCSR[ 217 ][ 32 ],
   alphaCSR[ 217 ][ 33 ],
   alphaCSR[ 217 ][ 34 ],
   alphaCSR[ 217 ][ 35 ],
   alphaCSR[ 217 ][ 36 ],
   alphaCSR[ 217 ][ 37 ],
   alphaCSR[ 217 ][ 38 ],
   alphaCSR[ 217 ][ 39 ],
   alphaCSR[ 217 ][ 40 ],
   alphaCSR[ 217 ][ 41 ],
   alphaCSR[ 217 ][ 42 ],
   alphaCSR[ 217 ][ 43 ],
   alphaCSR[ 217 ][ 44 ],
   alphaCSR[ 217 ][ 45 ],
   alphaCSR[ 217 ][ 46 ],
   alphaCSR[ 217 ][ 47 ],
   alphaCSR[ 217 ][ 48 ],
   alphaCSR[ 217 ][ 49 ],
   alphaCSR[ 217 ][ 50 ],
   alphaCSR[ 217 ][ 51 ],
   alphaCSR[ 217 ][ 52 ],
   alphaCSR[ 217 ][ 53 ],
   alphaCSR[ 217 ][ 54 ],
   alphaCSR[ 217 ][ 55 ],
   alphaCSR[ 217 ][ 56 ],
   alphaCSR[ 217 ][ 57 ],
   alphaCSR[ 217 ][ 58 ],
   alphaCSR[ 217 ][ 59 ],
   alphaCSR[ 217 ][ 60 ],
   alphaCSR[ 217 ][ 61 ],
   alphaCSR[ 217 ][ 62 ],
   alphaCSR[ 217 ][ 63 ],
   alphaCSR[ 217 ][ 64 ],
   alphaCSR[ 217 ][ 65 ],
   alphaCSR[ 217 ][ 66 ],
   alphaCSR[ 217 ][ 67 ],
   alphaCSR[ 217 ][ 68 ],
   alphaCSR[ 217 ][ 69 ],
   alphaCSR[ 217 ][ 70 ],
   alphaCSR[ 217 ][ 71 ],
   alphaCSR[ 217 ][ 72 ],
   alphaCSR[ 217 ][ 73 ],
   alphaCSR[ 217 ][ 74 ],
   alphaCSR[ 217 ][ 75 ],
   alphaCSR[ 217 ][ 76 ],
   alphaCSR[ 217 ][ 77 ],
   alphaCSR[ 217 ][ 78 ],
   alphaCSR[ 217 ][ 79 ],
   alphaCSR[ 217 ][ 80 ],
   alphaCSR[ 217 ][ 81 ],
   alphaCSR[ 217 ][ 82 ],
   alphaCSR[ 217 ][ 83 ],
   alphaCSR[ 217 ][ 84 ],
   alphaCSR[ 217 ][ 85 ],
   alphaCSR[ 217 ][ 86 ],
   alphaCSR[ 217 ][ 87 ],
   alphaCSR[ 217 ][ 88 ],
   alphaCSR[ 217 ][ 89 ],
   alphaCSR[ 217 ][ 90 ],
   alphaCSR[ 217 ][ 91 ],
   alphaCSR[ 217 ][ 92 ],
   alphaCSR[ 217 ][ 93 ],
   alphaCSR[ 217 ][ 94 ],
   alphaCSR[ 217 ][ 95 ],
   alphaCSR[ 217 ][ 96 ],
   alphaCSR[ 217 ][ 97 ],
   alphaCSR[ 217 ][ 98 ],
   alphaCSR[ 217 ][ 99 ],
   alphaCSR[ 217 ][ 100 ],
   alphaCSR[ 217 ][ 101 ],
   alphaCSR[ 217 ][ 102 ],
   alphaCSR[ 217 ][ 103 ],
   alphaCSR[ 217 ][ 104 ],
   alphaCSR[ 217 ][ 105 ],
   alphaCSR[ 217 ][ 106 ],
   alphaCSR[ 217 ][ 107 ],
   alphaCSR[ 217 ][ 108 ],
   alphaCSR[ 217 ][ 109 ],
   alphaCSR[ 217 ][ 110 ],
   alphaCSR[ 217 ][ 111 ],
   alphaCSR[ 217 ][ 112 ],
   alphaCSR[ 217 ][ 113 ],
   alphaCSR[ 217 ][ 114 ],
   alphaCSR[ 217 ][ 115 ],
   alphaCSR[ 217 ][ 116 ],
   alphaCSR[ 217 ][ 117 ],
   alphaCSR[ 217 ][ 118 ],
   alphaCSR[ 217 ][ 119 ],
   alphaCSR[ 217 ][ 120 ],
   alphaCSR[ 217 ][ 121 ],
   alphaCSR[ 217 ][ 122 ],
   alphaCSR[ 217 ][ 123 ],
   alphaCSR[ 217 ][ 124 ],
   alphaCSR[ 217 ][ 125 ],
   alphaCSR[ 217 ][ 126 ],
   alphaCSR[ 217 ][ 127 ],
   alphaCSR[ 217 ][ 128 ],
   alphaCSR[ 217 ][ 129 ],
   alphaCSR[ 217 ][ 130 ],
   alphaCSR[ 217 ][ 131 ],
   alphaCSR[ 217 ][ 132 ],
   alphaCSR[ 217 ][ 133 ],
   alphaCSR[ 217 ][ 134 ],
   alphaCSR[ 217 ][ 135 ],
   alphaCSR[ 217 ][ 136 ],
   alphaCSR[ 217 ][ 137 ],
   alphaCSR[ 217 ][ 138 ],
   alphaCSR[ 217 ][ 139 ],
   alphaCSR[ 217 ][ 140 ],
   alphaCSR[ 217 ][ 141 ],
   alphaCSR[ 217 ][ 142 ],
   alphaCSR[ 217 ][ 143 ],
   alphaCSR[ 217 ][ 144 ],
   alphaCSR[ 217 ][ 145 ],
   alphaCSR[ 217 ][ 146 ],
   alphaCSR[ 217 ][ 147 ],
   alphaCSR[ 217 ][ 148 ],
   alphaCSR[ 217 ][ 149 ],
   alphaCSR[ 217 ][ 150 ],
   alphaCSR[ 217 ][ 151 ],
   alphaCSR[ 217 ][ 152 ],
   alphaCSR[ 217 ][ 153 ],
   alphaCSR[ 217 ][ 154 ],
   alphaCSR[ 217 ][ 155 ],
   alphaCSR[ 217 ][ 156 ],
   alphaCSR[ 217 ][ 157 ],
   alphaCSR[ 217 ][ 158 ],
   alphaCSR[ 217 ][ 159 ],
   alphaCSR[ 217 ][ 160 ],
   alphaCSR[ 217 ][ 161 ],
   alphaCSR[ 217 ][ 162 ],
   alphaCSR[ 217 ][ 163 ],
   alphaCSR[ 217 ][ 164 ],
   alphaCSR[ 217 ][ 165 ],
   alphaCSR[ 217 ][ 166 ],
   alphaCSR[ 217 ][ 167 ],
   alphaCSR[ 217 ][ 168 ],
   alphaCSR[ 217 ][ 169 ],
   alphaCSR[ 217 ][ 170 ],
   alphaCSR[ 217 ][ 171 ],
   alphaCSR[ 217 ][ 172 ],
   alphaCSR[ 217 ][ 173 ],
   alphaCSR[ 217 ][ 174 ],
   alphaCSR[ 217 ][ 175 ],
   alphaCSR[ 217 ][ 176 ],
   alphaCSR[ 217 ][ 177 ],
   alphaCSR[ 217 ][ 178 ],
   alphaCSR[ 217 ][ 179 ],
   alphaCSR[ 217 ][ 180 ],
   alphaCSR[ 217 ][ 181 ],
   alphaCSR[ 217 ][ 182 ],
   alphaCSR[ 217 ][ 183 ],
   alphaCSR[ 217 ][ 184 ],
   alphaCSR[ 217 ][ 185 ],
   alphaCSR[ 217 ][ 186 ],
   alphaCSR[ 217 ][ 187 ],
   alphaCSR[ 217 ][ 188 ],
   alphaCSR[ 217 ][ 189 ],
   alphaCSR[ 217 ][ 190 ],
   alphaCSR[ 217 ][ 191 ],
   alphaCSR[ 217 ][ 192 ],
   alphaCSR[ 217 ][ 193 ],
   alphaCSR[ 217 ][ 194 ],
   alphaCSR[ 217 ][ 195 ],
   alphaCSR[ 217 ][ 196 ],
   alphaCSR[ 217 ][ 197 ],
   alphaCSR[ 217 ][ 198 ],
   alphaCSR[ 217 ][ 199 ],
   alphaCSR[ 217 ][ 200 ],
   alphaCSR[ 217 ][ 201 ],
   alphaCSR[ 217 ][ 202 ],
   alphaCSR[ 217 ][ 203 ],
   alphaCSR[ 217 ][ 204 ],
   alphaCSR[ 217 ][ 205 ],
   alphaCSR[ 217 ][ 206 ],
   alphaCSR[ 217 ][ 207 ],
   alphaCSR[ 217 ][ 208 ],
   alphaCSR[ 217 ][ 209 ],
   alphaCSR[ 217 ][ 210 ],
   alphaCSR[ 217 ][ 211 ],
   alphaCSR[ 217 ][ 212 ],
   alphaCSR[ 217 ][ 213 ],
   alphaCSR[ 217 ][ 214 ],
   alphaCSR[ 217 ][ 215 ],
   alphaCSR[ 217 ][ 216 ],
   alphaCSR[ 217 ][ 217 ],
   alphaCSR[ 217 ][ 218 ],
   alphaCSR[ 217 ][ 219 ],
   alphaCSR[ 217 ][ 220 ],
   alphaCSR[ 217 ][ 221 ],
   alphaCSR[ 217 ][ 222 ],
   alphaCSR[ 217 ][ 223 ],
   alphaCSR[ 217 ][ 224 ],
   alphaCSR[ 217 ][ 225 ],
   alphaCSR[ 217 ][ 226 ],
   alphaCSR[ 217 ][ 227 ],
   alphaCSR[ 217 ][ 228 ],
   alphaCSR[ 217 ][ 229 ],
   alphaCSR[ 217 ][ 230 ],
   alphaCSR[ 217 ][ 231 ],
   alphaCSR[ 217 ][ 232 ],
   alphaCSR[ 217 ][ 233 ],
   alphaCSR[ 217 ][ 234 ],
   alphaCSR[ 217 ][ 235 ],
   alphaCSR[ 217 ][ 236 ],
   alphaCSR[ 217 ][ 237 ],
   alphaCSR[ 217 ][ 238 ],
   alphaCSR[ 217 ][ 239 ],
   alphaCSR[ 217 ][ 240 ],
   alphaCSR[ 217 ][ 241 ],
   alphaCSR[ 217 ][ 242 ],
   alphaCSR[ 217 ][ 243 ],
   alphaCSR[ 217 ][ 244 ],
   alphaCSR[ 217 ][ 245 ],
   alphaCSR[ 217 ][ 246 ],
   alphaCSR[ 217 ][ 247 ],
   alphaCSR[ 217 ][ 248 ],
   alphaCSR[ 217 ][ 249 ],
   alphaCSR[ 217 ][ 250 ],
   alphaCSR[ 217 ][ 251 ],
   alphaCSR[ 217 ][ 252 ],
   alphaCSR[ 217 ][ 253 ],
   alphaCSR[ 217 ][ 254 ],
   alphaCSR[ 217 ][ 255 ],
   alphaCSR[ 217 ][ 256 ],
   alphaCSR[ 217 ][ 257 ],
   alphaCSR[ 217 ][ 258 ],
   alphaCSR[ 217 ][ 259 ],
   alphaCSR[ 217 ][ 260 ],
   alphaCSR[ 217 ][ 261 ],
   alphaCSR[ 217 ][ 262 ],
   alphaCSR[ 217 ][ 263 ],
   alphaCSR[ 217 ][ 264 ],
   alphaCSR[ 217 ][ 265 ],
   alphaCSR[ 217 ][ 266 ],
   alphaCSR[ 217 ][ 267 ],
   alphaCSR[ 217 ][ 268 ],
   alphaCSR[ 217 ][ 269 ],
   alphaCSR[ 217 ][ 270 ],
   alphaCSR[ 217 ][ 271 ],
   alphaCSR[ 217 ][ 272 ],
   alphaCSR[ 217 ][ 273 ],
   alphaCSR[ 217 ][ 274 ],
   alphaCSR[ 217 ][ 275 ],
   alphaCSR[ 217 ][ 276 ],
   alphaCSR[ 217 ][ 277 ],
   alphaCSR[ 217 ][ 278 ],
   alphaCSR[ 217 ][ 279 ],
   alphaCSR[ 217 ][ 280 ],
   alphaCSR[ 217 ][ 281 ],
   alphaCSR[ 217 ][ 282 ],
   alphaCSR[ 217 ][ 283 ],
   alphaCSR[ 217 ][ 284 ],
   alphaCSR[ 217 ][ 285 ],
   alphaCSR[ 217 ][ 286 ],
   alphaCSR[ 217 ][ 287 ],
   alphaCSR[ 217 ][ 288 ],
   alphaCSR[ 217 ][ 289 ],
   alphaCSR[ 217 ][ 290 ],
   alphaCSR[ 217 ][ 291 ],
   alphaCSR[ 217 ][ 292 ],
   alphaCSR[ 217 ][ 293 ],
   alphaCSR[ 217 ][ 294 ],
   alphaCSR[ 217 ][ 295 ],
   alphaCSR[ 217 ][ 296 ],
   alphaCSR[ 217 ][ 297 ],
   alphaCSR[ 217 ][ 298 ],
   alphaCSR[ 217 ][ 299 ],
   alphaCSR[ 217 ][ 300 ],
   alphaCSR[ 217 ][ 301 ],
   alphaCSR[ 217 ][ 302 ],
   alphaCSR[ 217 ][ 303 ],
   alphaCSR[ 217 ][ 304 ],
   alphaCSR[ 217 ][ 305 ],
   alphaCSR[ 217 ][ 306 ],
   alphaCSR[ 217 ][ 307 ],
   alphaCSR[ 217 ][ 308 ],
   alphaCSR[ 217 ][ 309 ],
   alphaCSR[ 217 ][ 310 ],
   alphaCSR[ 217 ][ 311 ],
   alphaCSR[ 217 ][ 312 ],
   alphaCSR[ 217 ][ 313 ],
   alphaCSR[ 217 ][ 314 ],
   alphaCSR[ 217 ][ 315 ],
   alphaCSR[ 217 ][ 316 ],
   alphaCSR[ 217 ][ 317 ],
   alphaCSR[ 217 ][ 318 ],
   alphaCSR[ 217 ][ 319 ],
   alphaCSR[ 217 ][ 320 ],
   alphaCSR[ 217 ][ 321 ],
   alphaCSR[ 217 ][ 322 ],
   alphaCSR[ 217 ][ 323 ],
   alphaCSR[ 217 ][ 324 ],
   alphaCSR[ 217 ][ 325 ],
   alphaCSR[ 217 ][ 326 ],
   alphaCSR[ 217 ][ 327 ],
   alphaCSR[ 217 ][ 328 ],
   alphaCSR[ 217 ][ 329 ],
   alphaCSR[ 217 ][ 330 ],
   alphaCSR[ 217 ][ 331 ],
   alphaCSR[ 217 ][ 332 ],
   alphaCSR[ 217 ][ 333 ],
   alphaCSR[ 217 ][ 334 ],
   alphaCSR[ 217 ][ 335 ],
   alphaCSR[ 217 ][ 336 ],
   alphaCSR[ 217 ][ 337 ],
   alphaCSR[ 217 ][ 338 ],
   alphaCSR[ 217 ][ 339 ],
   alphaCSR[ 217 ][ 340 ],
   alphaCSR[ 217 ][ 341 ],
   alphaCSR[ 217 ][ 342 ],
   alphaCSR[ 217 ][ 343 ],
   alphaCSR[ 217 ][ 344 ],
   alphaCSR[ 217 ][ 345 ],
   alphaCSR[ 217 ][ 346 ],
   alphaCSR[ 217 ][ 347 ],
   alphaCSR[ 217 ][ 348 ],
   alphaCSR[ 217 ][ 349 ],
   alphaCSR[ 217 ][ 350 ],
   alphaCSR[ 217 ][ 351 ],
   alphaCSR[ 217 ][ 352 ],
   alphaCSR[ 217 ][ 353 ],
   alphaCSR[ 217 ][ 354 ],
   alphaCSR[ 217 ][ 355 ],
   alphaCSR[ 217 ][ 356 ],
   alphaCSR[ 217 ][ 357 ],
   alphaCSR[ 217 ][ 358 ],
   alphaCSR[ 217 ][ 359 ],
   alphaCSR[ 217 ][ 360 ],
   alphaCSR[ 217 ][ 361 ],
   alphaCSR[ 217 ][ 362 ],
   alphaCSR[ 217 ][ 363 ],
   alphaCSR[ 217 ][ 364 ],
   alphaCSR[ 217 ][ 365 ],
   alphaCSR[ 217 ][ 366 ],
   alphaCSR[ 217 ][ 367 ],
   alphaCSR[ 217 ][ 368 ],
   alphaCSR[ 217 ][ 369 ],
   alphaCSR[ 217 ][ 370 ],
   alphaCSR[ 217 ][ 371 ],
   alphaCSR[ 217 ][ 372 ],
   alphaCSR[ 217 ][ 373 ],
   alphaCSR[ 217 ][ 374 ],
   alphaCSR[ 217 ][ 375 ],
   alphaCSR[ 217 ][ 376 ],
   alphaCSR[ 217 ][ 377 ],
   alphaCSR[ 217 ][ 378 ],
   alphaCSR[ 217 ][ 379 ],
   alphaCSR[ 217 ][ 380 ],
   alphaCSR[ 217 ][ 381 ],
   alphaCSR[ 217 ][ 382 ],
   alphaCSR[ 217 ][ 383 ],
   alphaCSR[ 218 ][ 0 ],
   alphaCSR[ 218 ][ 1 ],
   alphaCSR[ 218 ][ 2 ],
   alphaCSR[ 218 ][ 3 ],
   alphaCSR[ 218 ][ 4 ],
   alphaCSR[ 218 ][ 5 ],
   alphaCSR[ 218 ][ 6 ],
   alphaCSR[ 218 ][ 7 ],
   alphaCSR[ 218 ][ 8 ],
   alphaCSR[ 218 ][ 9 ],
   alphaCSR[ 218 ][ 10 ],
   alphaCSR[ 218 ][ 11 ],
   alphaCSR[ 218 ][ 12 ],
   alphaCSR[ 218 ][ 13 ],
   alphaCSR[ 218 ][ 14 ],
   alphaCSR[ 218 ][ 15 ],
   alphaCSR[ 218 ][ 16 ],
   alphaCSR[ 218 ][ 17 ],
   alphaCSR[ 218 ][ 18 ],
   alphaCSR[ 218 ][ 19 ],
   alphaCSR[ 218 ][ 20 ],
   alphaCSR[ 218 ][ 21 ],
   alphaCSR[ 218 ][ 22 ],
   alphaCSR[ 218 ][ 23 ],
   alphaCSR[ 218 ][ 24 ],
   alphaCSR[ 218 ][ 25 ],
   alphaCSR[ 218 ][ 26 ],
   alphaCSR[ 218 ][ 27 ],
   alphaCSR[ 218 ][ 28 ],
   alphaCSR[ 218 ][ 29 ],
   alphaCSR[ 218 ][ 30 ],
   alphaCSR[ 218 ][ 31 ],
   alphaCSR[ 218 ][ 32 ],
   alphaCSR[ 218 ][ 33 ],
   alphaCSR[ 218 ][ 34 ],
   alphaCSR[ 218 ][ 35 ],
   alphaCSR[ 218 ][ 36 ],
   alphaCSR[ 218 ][ 37 ],
   alphaCSR[ 218 ][ 38 ],
   alphaCSR[ 218 ][ 39 ],
   alphaCSR[ 218 ][ 40 ],
   alphaCSR[ 218 ][ 41 ],
   alphaCSR[ 218 ][ 42 ],
   alphaCSR[ 218 ][ 43 ],
   alphaCSR[ 218 ][ 44 ],
   alphaCSR[ 218 ][ 45 ],
   alphaCSR[ 218 ][ 46 ],
   alphaCSR[ 218 ][ 47 ],
   alphaCSR[ 218 ][ 48 ],
   alphaCSR[ 218 ][ 49 ],
   alphaCSR[ 218 ][ 50 ],
   alphaCSR[ 218 ][ 51 ],
   alphaCSR[ 218 ][ 52 ],
   alphaCSR[ 218 ][ 53 ],
   alphaCSR[ 218 ][ 54 ],
   alphaCSR[ 218 ][ 55 ],
   alphaCSR[ 218 ][ 56 ],
   alphaCSR[ 218 ][ 57 ],
   alphaCSR[ 218 ][ 58 ],
   alphaCSR[ 218 ][ 59 ],
   alphaCSR[ 218 ][ 60 ],
   alphaCSR[ 218 ][ 61 ],
   alphaCSR[ 218 ][ 62 ],
   alphaCSR[ 218 ][ 63 ],
   alphaCSR[ 218 ][ 64 ],
   alphaCSR[ 218 ][ 65 ],
   alphaCSR[ 218 ][ 66 ],
   alphaCSR[ 218 ][ 67 ],
   alphaCSR[ 218 ][ 68 ],
   alphaCSR[ 218 ][ 69 ],
   alphaCSR[ 218 ][ 70 ],
   alphaCSR[ 218 ][ 71 ],
   alphaCSR[ 218 ][ 72 ],
   alphaCSR[ 218 ][ 73 ],
   alphaCSR[ 218 ][ 74 ],
   alphaCSR[ 218 ][ 75 ],
   alphaCSR[ 218 ][ 76 ],
   alphaCSR[ 218 ][ 77 ],
   alphaCSR[ 218 ][ 78 ],
   alphaCSR[ 218 ][ 79 ],
   alphaCSR[ 218 ][ 80 ],
   alphaCSR[ 218 ][ 81 ],
   alphaCSR[ 218 ][ 82 ],
   alphaCSR[ 218 ][ 83 ],
   alphaCSR[ 218 ][ 84 ],
   alphaCSR[ 218 ][ 85 ],
   alphaCSR[ 218 ][ 86 ],
   alphaCSR[ 218 ][ 87 ],
   alphaCSR[ 218 ][ 88 ],
   alphaCSR[ 218 ][ 89 ],
   alphaCSR[ 218 ][ 90 ],
   alphaCSR[ 218 ][ 91 ],
   alphaCSR[ 218 ][ 92 ],
   alphaCSR[ 218 ][ 93 ],
   alphaCSR[ 218 ][ 94 ],
   alphaCSR[ 218 ][ 95 ],
   alphaCSR[ 218 ][ 96 ],
   alphaCSR[ 218 ][ 97 ],
   alphaCSR[ 218 ][ 98 ],
   alphaCSR[ 218 ][ 99 ],
   alphaCSR[ 218 ][ 100 ],
   alphaCSR[ 218 ][ 101 ],
   alphaCSR[ 218 ][ 102 ],
   alphaCSR[ 218 ][ 103 ],
   alphaCSR[ 218 ][ 104 ],
   alphaCSR[ 218 ][ 105 ],
   alphaCSR[ 218 ][ 106 ],
   alphaCSR[ 218 ][ 107 ],
   alphaCSR[ 218 ][ 108 ],
   alphaCSR[ 218 ][ 109 ],
   alphaCSR[ 218 ][ 110 ],
   alphaCSR[ 218 ][ 111 ],
   alphaCSR[ 218 ][ 112 ],
   alphaCSR[ 218 ][ 113 ],
   alphaCSR[ 218 ][ 114 ],
   alphaCSR[ 218 ][ 115 ],
   alphaCSR[ 218 ][ 116 ],
   alphaCSR[ 218 ][ 117 ],
   alphaCSR[ 218 ][ 118 ],
   alphaCSR[ 218 ][ 119 ],
   alphaCSR[ 218 ][ 120 ],
   alphaCSR[ 218 ][ 121 ],
   alphaCSR[ 218 ][ 122 ],
   alphaCSR[ 218 ][ 123 ],
   alphaCSR[ 218 ][ 124 ],
   alphaCSR[ 218 ][ 125 ],
   alphaCSR[ 218 ][ 126 ],
   alphaCSR[ 218 ][ 127 ],
   alphaCSR[ 218 ][ 128 ],
   alphaCSR[ 218 ][ 129 ],
   alphaCSR[ 218 ][ 130 ],
   alphaCSR[ 218 ][ 131 ],
   alphaCSR[ 218 ][ 132 ],
   alphaCSR[ 218 ][ 133 ],
   alphaCSR[ 218 ][ 134 ],
   alphaCSR[ 218 ][ 135 ],
   alphaCSR[ 218 ][ 136 ],
   alphaCSR[ 218 ][ 137 ],
   alphaCSR[ 218 ][ 138 ],
   alphaCSR[ 218 ][ 139 ],
   alphaCSR[ 218 ][ 140 ],
   alphaCSR[ 218 ][ 141 ],
   alphaCSR[ 218 ][ 142 ],
   alphaCSR[ 218 ][ 143 ],
   alphaCSR[ 218 ][ 144 ],
   alphaCSR[ 218 ][ 145 ],
   alphaCSR[ 218 ][ 146 ],
   alphaCSR[ 218 ][ 147 ],
   alphaCSR[ 218 ][ 148 ],
   alphaCSR[ 218 ][ 149 ],
   alphaCSR[ 218 ][ 150 ],
   alphaCSR[ 218 ][ 151 ],
   alphaCSR[ 218 ][ 152 ],
   alphaCSR[ 218 ][ 153 ],
   alphaCSR[ 218 ][ 154 ],
   alphaCSR[ 218 ][ 155 ],
   alphaCSR[ 218 ][ 156 ],
   alphaCSR[ 218 ][ 157 ],
   alphaCSR[ 218 ][ 158 ],
   alphaCSR[ 218 ][ 159 ],
   alphaCSR[ 218 ][ 160 ],
   alphaCSR[ 218 ][ 161 ],
   alphaCSR[ 218 ][ 162 ],
   alphaCSR[ 218 ][ 163 ],
   alphaCSR[ 218 ][ 164 ],
   alphaCSR[ 218 ][ 165 ],
   alphaCSR[ 218 ][ 166 ],
   alphaCSR[ 218 ][ 167 ],
   alphaCSR[ 218 ][ 168 ],
   alphaCSR[ 218 ][ 169 ],
   alphaCSR[ 218 ][ 170 ],
   alphaCSR[ 218 ][ 171 ],
   alphaCSR[ 218 ][ 172 ],
   alphaCSR[ 218 ][ 173 ],
   alphaCSR[ 218 ][ 174 ],
   alphaCSR[ 218 ][ 175 ],
   alphaCSR[ 218 ][ 176 ],
   alphaCSR[ 218 ][ 177 ],
   alphaCSR[ 218 ][ 178 ],
   alphaCSR[ 218 ][ 179 ],
   alphaCSR[ 218 ][ 180 ],
   alphaCSR[ 218 ][ 181 ],
   alphaCSR[ 218 ][ 182 ],
   alphaCSR[ 218 ][ 183 ],
   alphaCSR[ 218 ][ 184 ],
   alphaCSR[ 218 ][ 185 ],
   alphaCSR[ 218 ][ 186 ],
   alphaCSR[ 218 ][ 187 ],
   alphaCSR[ 218 ][ 188 ],
   alphaCSR[ 218 ][ 189 ],
   alphaCSR[ 218 ][ 190 ],
   alphaCSR[ 218 ][ 191 ],
   alphaCSR[ 218 ][ 192 ],
   alphaCSR[ 218 ][ 193 ],
   alphaCSR[ 218 ][ 194 ],
   alphaCSR[ 218 ][ 195 ],
   alphaCSR[ 218 ][ 196 ],
   alphaCSR[ 218 ][ 197 ],
   alphaCSR[ 218 ][ 198 ],
   alphaCSR[ 218 ][ 199 ],
   alphaCSR[ 218 ][ 200 ],
   alphaCSR[ 218 ][ 201 ],
   alphaCSR[ 218 ][ 202 ],
   alphaCSR[ 218 ][ 203 ],
   alphaCSR[ 218 ][ 204 ],
   alphaCSR[ 218 ][ 205 ],
   alphaCSR[ 218 ][ 206 ],
   alphaCSR[ 218 ][ 207 ],
   alphaCSR[ 218 ][ 208 ],
   alphaCSR[ 218 ][ 209 ],
   alphaCSR[ 218 ][ 210 ],
   alphaCSR[ 218 ][ 211 ],
   alphaCSR[ 218 ][ 212 ],
   alphaCSR[ 218 ][ 213 ],
   alphaCSR[ 218 ][ 214 ],
   alphaCSR[ 218 ][ 215 ],
   alphaCSR[ 218 ][ 216 ],
   alphaCSR[ 218 ][ 217 ],
   alphaCSR[ 218 ][ 218 ],
   alphaCSR[ 218 ][ 219 ],
   alphaCSR[ 218 ][ 220 ],
   alphaCSR[ 218 ][ 221 ],
   alphaCSR[ 218 ][ 222 ],
   alphaCSR[ 218 ][ 223 ],
   alphaCSR[ 218 ][ 224 ],
   alphaCSR[ 218 ][ 225 ],
   alphaCSR[ 218 ][ 226 ],
   alphaCSR[ 218 ][ 227 ],
   alphaCSR[ 218 ][ 228 ],
   alphaCSR[ 218 ][ 229 ],
   alphaCSR[ 218 ][ 230 ],
   alphaCSR[ 218 ][ 231 ],
   alphaCSR[ 218 ][ 232 ],
   alphaCSR[ 218 ][ 233 ],
   alphaCSR[ 218 ][ 234 ],
   alphaCSR[ 218 ][ 235 ],
   alphaCSR[ 218 ][ 236 ],
   alphaCSR[ 218 ][ 237 ],
   alphaCSR[ 218 ][ 238 ],
   alphaCSR[ 218 ][ 239 ],
   alphaCSR[ 218 ][ 240 ],
   alphaCSR[ 218 ][ 241 ],
   alphaCSR[ 218 ][ 242 ],
   alphaCSR[ 218 ][ 243 ],
   alphaCSR[ 218 ][ 244 ],
   alphaCSR[ 218 ][ 245 ],
   alphaCSR[ 218 ][ 246 ],
   alphaCSR[ 218 ][ 247 ],
   alphaCSR[ 218 ][ 248 ],
   alphaCSR[ 218 ][ 249 ],
   alphaCSR[ 218 ][ 250 ],
   alphaCSR[ 218 ][ 251 ],
   alphaCSR[ 218 ][ 252 ],
   alphaCSR[ 218 ][ 253 ],
   alphaCSR[ 218 ][ 254 ],
   alphaCSR[ 218 ][ 255 ],
   alphaCSR[ 218 ][ 256 ],
   alphaCSR[ 218 ][ 257 ],
   alphaCSR[ 218 ][ 258 ],
   alphaCSR[ 218 ][ 259 ],
   alphaCSR[ 218 ][ 260 ],
   alphaCSR[ 218 ][ 261 ],
   alphaCSR[ 218 ][ 262 ],
   alphaCSR[ 218 ][ 263 ],
   alphaCSR[ 218 ][ 264 ],
   alphaCSR[ 218 ][ 265 ],
   alphaCSR[ 218 ][ 266 ],
   alphaCSR[ 218 ][ 267 ],
   alphaCSR[ 218 ][ 268 ],
   alphaCSR[ 218 ][ 269 ],
   alphaCSR[ 218 ][ 270 ],
   alphaCSR[ 218 ][ 271 ],
   alphaCSR[ 218 ][ 272 ],
   alphaCSR[ 218 ][ 273 ],
   alphaCSR[ 218 ][ 274 ],
   alphaCSR[ 218 ][ 275 ],
   alphaCSR[ 218 ][ 276 ],
   alphaCSR[ 218 ][ 277 ],
   alphaCSR[ 218 ][ 278 ],
   alphaCSR[ 218 ][ 279 ],
   alphaCSR[ 218 ][ 280 ],
   alphaCSR[ 218 ][ 281 ],
   alphaCSR[ 218 ][ 282 ],
   alphaCSR[ 218 ][ 283 ],
   alphaCSR[ 218 ][ 284 ],
   alphaCSR[ 218 ][ 285 ],
   alphaCSR[ 218 ][ 286 ],
   alphaCSR[ 218 ][ 287 ],
   alphaCSR[ 218 ][ 288 ],
   alphaCSR[ 218 ][ 289 ],
   alphaCSR[ 218 ][ 290 ],
   alphaCSR[ 218 ][ 291 ],
   alphaCSR[ 218 ][ 292 ],
   alphaCSR[ 218 ][ 293 ],
   alphaCSR[ 218 ][ 294 ],
   alphaCSR[ 218 ][ 295 ],
   alphaCSR[ 218 ][ 296 ],
   alphaCSR[ 218 ][ 297 ],
   alphaCSR[ 218 ][ 298 ],
   alphaCSR[ 218 ][ 299 ],
   alphaCSR[ 218 ][ 300 ],
   alphaCSR[ 218 ][ 301 ],
   alphaCSR[ 218 ][ 302 ],
   alphaCSR[ 218 ][ 303 ],
   alphaCSR[ 218 ][ 304 ],
   alphaCSR[ 218 ][ 305 ],
   alphaCSR[ 218 ][ 306 ],
   alphaCSR[ 218 ][ 307 ],
   alphaCSR[ 218 ][ 308 ],
   alphaCSR[ 218 ][ 309 ],
   alphaCSR[ 218 ][ 310 ],
   alphaCSR[ 218 ][ 311 ],
   alphaCSR[ 218 ][ 312 ],
   alphaCSR[ 218 ][ 313 ],
   alphaCSR[ 218 ][ 314 ],
   alphaCSR[ 218 ][ 315 ],
   alphaCSR[ 218 ][ 316 ],
   alphaCSR[ 218 ][ 317 ],
   alphaCSR[ 218 ][ 318 ],
   alphaCSR[ 218 ][ 319 ],
   alphaCSR[ 218 ][ 320 ],
   alphaCSR[ 218 ][ 321 ],
   alphaCSR[ 218 ][ 322 ],
   alphaCSR[ 218 ][ 323 ],
   alphaCSR[ 218 ][ 324 ],
   alphaCSR[ 218 ][ 325 ],
   alphaCSR[ 218 ][ 326 ],
   alphaCSR[ 218 ][ 327 ],
   alphaCSR[ 218 ][ 328 ],
   alphaCSR[ 218 ][ 329 ],
   alphaCSR[ 218 ][ 330 ],
   alphaCSR[ 218 ][ 331 ],
   alphaCSR[ 218 ][ 332 ],
   alphaCSR[ 218 ][ 333 ],
   alphaCSR[ 218 ][ 334 ],
   alphaCSR[ 218 ][ 335 ],
   alphaCSR[ 218 ][ 336 ],
   alphaCSR[ 218 ][ 337 ],
   alphaCSR[ 218 ][ 338 ],
   alphaCSR[ 218 ][ 339 ],
   alphaCSR[ 218 ][ 340 ],
   alphaCSR[ 218 ][ 341 ],
   alphaCSR[ 218 ][ 342 ],
   alphaCSR[ 218 ][ 343 ],
   alphaCSR[ 218 ][ 344 ],
   alphaCSR[ 218 ][ 345 ],
   alphaCSR[ 218 ][ 346 ],
   alphaCSR[ 218 ][ 347 ],
   alphaCSR[ 218 ][ 348 ],
   alphaCSR[ 218 ][ 349 ],
   alphaCSR[ 218 ][ 350 ],
   alphaCSR[ 218 ][ 351 ],
   alphaCSR[ 218 ][ 352 ],
   alphaCSR[ 218 ][ 353 ],
   alphaCSR[ 218 ][ 354 ],
   alphaCSR[ 218 ][ 355 ],
   alphaCSR[ 218 ][ 356 ],
   alphaCSR[ 218 ][ 357 ],
   alphaCSR[ 218 ][ 358 ],
   alphaCSR[ 218 ][ 359 ],
   alphaCSR[ 218 ][ 360 ],
   alphaCSR[ 218 ][ 361 ],
   alphaCSR[ 218 ][ 362 ],
   alphaCSR[ 218 ][ 363 ],
   alphaCSR[ 218 ][ 364 ],
   alphaCSR[ 218 ][ 365 ],
   alphaCSR[ 218 ][ 366 ],
   alphaCSR[ 218 ][ 367 ],
   alphaCSR[ 218 ][ 368 ],
   alphaCSR[ 218 ][ 369 ],
   alphaCSR[ 218 ][ 370 ],
   alphaCSR[ 218 ][ 371 ],
   alphaCSR[ 218 ][ 372 ],
   alphaCSR[ 218 ][ 373 ],
   alphaCSR[ 218 ][ 374 ],
   alphaCSR[ 218 ][ 375 ],
   alphaCSR[ 218 ][ 376 ],
   alphaCSR[ 218 ][ 377 ],
   alphaCSR[ 218 ][ 378 ],
   alphaCSR[ 218 ][ 379 ],
   alphaCSR[ 218 ][ 380 ],
   alphaCSR[ 218 ][ 381 ],
   alphaCSR[ 218 ][ 382 ],
   alphaCSR[ 218 ][ 383 ],
   alphaCSR[ 219 ][ 0 ],
   alphaCSR[ 219 ][ 1 ],
   alphaCSR[ 219 ][ 2 ],
   alphaCSR[ 219 ][ 3 ],
   alphaCSR[ 219 ][ 4 ],
   alphaCSR[ 219 ][ 5 ],
   alphaCSR[ 219 ][ 6 ],
   alphaCSR[ 219 ][ 7 ],
   alphaCSR[ 219 ][ 8 ],
   alphaCSR[ 219 ][ 9 ],
   alphaCSR[ 219 ][ 10 ],
   alphaCSR[ 219 ][ 11 ],
   alphaCSR[ 219 ][ 12 ],
   alphaCSR[ 219 ][ 13 ],
   alphaCSR[ 219 ][ 14 ],
   alphaCSR[ 219 ][ 15 ],
   alphaCSR[ 219 ][ 16 ],
   alphaCSR[ 219 ][ 17 ],
   alphaCSR[ 219 ][ 18 ],
   alphaCSR[ 219 ][ 19 ],
   alphaCSR[ 219 ][ 20 ],
   alphaCSR[ 219 ][ 21 ],
   alphaCSR[ 219 ][ 22 ],
   alphaCSR[ 219 ][ 23 ],
   alphaCSR[ 219 ][ 24 ],
   alphaCSR[ 219 ][ 25 ],
   alphaCSR[ 219 ][ 26 ],
   alphaCSR[ 219 ][ 27 ],
   alphaCSR[ 219 ][ 28 ],
   alphaCSR[ 219 ][ 29 ],
   alphaCSR[ 219 ][ 30 ],
   alphaCSR[ 219 ][ 31 ],
   alphaCSR[ 219 ][ 32 ],
   alphaCSR[ 219 ][ 33 ],
   alphaCSR[ 219 ][ 34 ],
   alphaCSR[ 219 ][ 35 ],
   alphaCSR[ 219 ][ 36 ],
   alphaCSR[ 219 ][ 37 ],
   alphaCSR[ 219 ][ 38 ],
   alphaCSR[ 219 ][ 39 ],
   alphaCSR[ 219 ][ 40 ],
   alphaCSR[ 219 ][ 41 ],
   alphaCSR[ 219 ][ 42 ],
   alphaCSR[ 219 ][ 43 ],
   alphaCSR[ 219 ][ 44 ],
   alphaCSR[ 219 ][ 45 ],
   alphaCSR[ 219 ][ 46 ],
   alphaCSR[ 219 ][ 47 ],
   alphaCSR[ 219 ][ 48 ],
   alphaCSR[ 219 ][ 49 ],
   alphaCSR[ 219 ][ 50 ],
   alphaCSR[ 219 ][ 51 ],
   alphaCSR[ 219 ][ 52 ],
   alphaCSR[ 219 ][ 53 ],
   alphaCSR[ 219 ][ 54 ],
   alphaCSR[ 219 ][ 55 ],
   alphaCSR[ 219 ][ 56 ],
   alphaCSR[ 219 ][ 57 ],
   alphaCSR[ 219 ][ 58 ],
   alphaCSR[ 219 ][ 59 ],
   alphaCSR[ 219 ][ 60 ],
   alphaCSR[ 219 ][ 61 ],
   alphaCSR[ 219 ][ 62 ],
   alphaCSR[ 219 ][ 63 ],
   alphaCSR[ 219 ][ 64 ],
   alphaCSR[ 219 ][ 65 ],
   alphaCSR[ 219 ][ 66 ],
   alphaCSR[ 219 ][ 67 ],
   alphaCSR[ 219 ][ 68 ],
   alphaCSR[ 219 ][ 69 ],
   alphaCSR[ 219 ][ 70 ],
   alphaCSR[ 219 ][ 71 ],
   alphaCSR[ 219 ][ 72 ],
   alphaCSR[ 219 ][ 73 ],
   alphaCSR[ 219 ][ 74 ],
   alphaCSR[ 219 ][ 75 ],
   alphaCSR[ 219 ][ 76 ],
   alphaCSR[ 219 ][ 77 ],
   alphaCSR[ 219 ][ 78 ],
   alphaCSR[ 219 ][ 79 ],
   alphaCSR[ 219 ][ 80 ],
   alphaCSR[ 219 ][ 81 ],
   alphaCSR[ 219 ][ 82 ],
   alphaCSR[ 219 ][ 83 ],
   alphaCSR[ 219 ][ 84 ],
   alphaCSR[ 219 ][ 85 ],
   alphaCSR[ 219 ][ 86 ],
   alphaCSR[ 219 ][ 87 ],
   alphaCSR[ 219 ][ 88 ],
   alphaCSR[ 219 ][ 89 ],
   alphaCSR[ 219 ][ 90 ],
   alphaCSR[ 219 ][ 91 ],
   alphaCSR[ 219 ][ 92 ],
   alphaCSR[ 219 ][ 93 ],
   alphaCSR[ 219 ][ 94 ],
   alphaCSR[ 219 ][ 95 ],
   alphaCSR[ 219 ][ 96 ],
   alphaCSR[ 219 ][ 97 ],
   alphaCSR[ 219 ][ 98 ],
   alphaCSR[ 219 ][ 99 ],
   alphaCSR[ 219 ][ 100 ],
   alphaCSR[ 219 ][ 101 ],
   alphaCSR[ 219 ][ 102 ],
   alphaCSR[ 219 ][ 103 ],
   alphaCSR[ 219 ][ 104 ],
   alphaCSR[ 219 ][ 105 ],
   alphaCSR[ 219 ][ 106 ],
   alphaCSR[ 219 ][ 107 ],
   alphaCSR[ 219 ][ 108 ],
   alphaCSR[ 219 ][ 109 ],
   alphaCSR[ 219 ][ 110 ],
   alphaCSR[ 219 ][ 111 ],
   alphaCSR[ 219 ][ 112 ],
   alphaCSR[ 219 ][ 113 ],
   alphaCSR[ 219 ][ 114 ],
   alphaCSR[ 219 ][ 115 ],
   alphaCSR[ 219 ][ 116 ],
   alphaCSR[ 219 ][ 117 ],
   alphaCSR[ 219 ][ 118 ],
   alphaCSR[ 219 ][ 119 ],
   alphaCSR[ 219 ][ 120 ],
   alphaCSR[ 219 ][ 121 ],
   alphaCSR[ 219 ][ 122 ],
   alphaCSR[ 219 ][ 123 ],
   alphaCSR[ 219 ][ 124 ],
   alphaCSR[ 219 ][ 125 ],
   alphaCSR[ 219 ][ 126 ],
   alphaCSR[ 219 ][ 127 ],
   alphaCSR[ 219 ][ 128 ],
   alphaCSR[ 219 ][ 129 ],
   alphaCSR[ 219 ][ 130 ],
   alphaCSR[ 219 ][ 131 ],
   alphaCSR[ 219 ][ 132 ],
   alphaCSR[ 219 ][ 133 ],
   alphaCSR[ 219 ][ 134 ],
   alphaCSR[ 219 ][ 135 ],
   alphaCSR[ 219 ][ 136 ],
   alphaCSR[ 219 ][ 137 ],
   alphaCSR[ 219 ][ 138 ],
   alphaCSR[ 219 ][ 139 ],
   alphaCSR[ 219 ][ 140 ],
   alphaCSR[ 219 ][ 141 ],
   alphaCSR[ 219 ][ 142 ],
   alphaCSR[ 219 ][ 143 ],
   alphaCSR[ 219 ][ 144 ],
   alphaCSR[ 219 ][ 145 ],
   alphaCSR[ 219 ][ 146 ],
   alphaCSR[ 219 ][ 147 ],
   alphaCSR[ 219 ][ 148 ],
   alphaCSR[ 219 ][ 149 ],
   alphaCSR[ 219 ][ 150 ],
   alphaCSR[ 219 ][ 151 ],
   alphaCSR[ 219 ][ 152 ],
   alphaCSR[ 219 ][ 153 ],
   alphaCSR[ 219 ][ 154 ],
   alphaCSR[ 219 ][ 155 ],
   alphaCSR[ 219 ][ 156 ],
   alphaCSR[ 219 ][ 157 ],
   alphaCSR[ 219 ][ 158 ],
   alphaCSR[ 219 ][ 159 ],
   alphaCSR[ 219 ][ 160 ],
   alphaCSR[ 219 ][ 161 ],
   alphaCSR[ 219 ][ 162 ],
   alphaCSR[ 219 ][ 163 ],
   alphaCSR[ 219 ][ 164 ],
   alphaCSR[ 219 ][ 165 ],
   alphaCSR[ 219 ][ 166 ],
   alphaCSR[ 219 ][ 167 ],
   alphaCSR[ 219 ][ 168 ],
   alphaCSR[ 219 ][ 169 ],
   alphaCSR[ 219 ][ 170 ],
   alphaCSR[ 219 ][ 171 ],
   alphaCSR[ 219 ][ 172 ],
   alphaCSR[ 219 ][ 173 ],
   alphaCSR[ 219 ][ 174 ],
   alphaCSR[ 219 ][ 175 ],
   alphaCSR[ 219 ][ 176 ],
   alphaCSR[ 219 ][ 177 ],
   alphaCSR[ 219 ][ 178 ],
   alphaCSR[ 219 ][ 179 ],
   alphaCSR[ 219 ][ 180 ],
   alphaCSR[ 219 ][ 181 ],
   alphaCSR[ 219 ][ 182 ],
   alphaCSR[ 219 ][ 183 ],
   alphaCSR[ 219 ][ 184 ],
   alphaCSR[ 219 ][ 185 ],
   alphaCSR[ 219 ][ 186 ],
   alphaCSR[ 219 ][ 187 ],
   alphaCSR[ 219 ][ 188 ],
   alphaCSR[ 219 ][ 189 ],
   alphaCSR[ 219 ][ 190 ],
   alphaCSR[ 219 ][ 191 ],
   alphaCSR[ 219 ][ 192 ],
   alphaCSR[ 219 ][ 193 ],
   alphaCSR[ 219 ][ 194 ],
   alphaCSR[ 219 ][ 195 ],
   alphaCSR[ 219 ][ 196 ],
   alphaCSR[ 219 ][ 197 ],
   alphaCSR[ 219 ][ 198 ],
   alphaCSR[ 219 ][ 199 ],
   alphaCSR[ 219 ][ 200 ],
   alphaCSR[ 219 ][ 201 ],
   alphaCSR[ 219 ][ 202 ],
   alphaCSR[ 219 ][ 203 ],
   alphaCSR[ 219 ][ 204 ],
   alphaCSR[ 219 ][ 205 ],
   alphaCSR[ 219 ][ 206 ],
   alphaCSR[ 219 ][ 207 ],
   alphaCSR[ 219 ][ 208 ],
   alphaCSR[ 219 ][ 209 ],
   alphaCSR[ 219 ][ 210 ],
   alphaCSR[ 219 ][ 211 ],
   alphaCSR[ 219 ][ 212 ],
   alphaCSR[ 219 ][ 213 ],
   alphaCSR[ 219 ][ 214 ],
   alphaCSR[ 219 ][ 215 ],
   alphaCSR[ 219 ][ 216 ],
   alphaCSR[ 219 ][ 217 ],
   alphaCSR[ 219 ][ 218 ],
   alphaCSR[ 219 ][ 219 ],
   alphaCSR[ 219 ][ 220 ],
   alphaCSR[ 219 ][ 221 ],
   alphaCSR[ 219 ][ 222 ],
   alphaCSR[ 219 ][ 223 ],
   alphaCSR[ 219 ][ 224 ],
   alphaCSR[ 219 ][ 225 ],
   alphaCSR[ 219 ][ 226 ],
   alphaCSR[ 219 ][ 227 ],
   alphaCSR[ 219 ][ 228 ],
   alphaCSR[ 219 ][ 229 ],
   alphaCSR[ 219 ][ 230 ],
   alphaCSR[ 219 ][ 231 ],
   alphaCSR[ 219 ][ 232 ],
   alphaCSR[ 219 ][ 233 ],
   alphaCSR[ 219 ][ 234 ],
   alphaCSR[ 219 ][ 235 ],
   alphaCSR[ 219 ][ 236 ],
   alphaCSR[ 219 ][ 237 ],
   alphaCSR[ 219 ][ 238 ],
   alphaCSR[ 219 ][ 239 ],
   alphaCSR[ 219 ][ 240 ],
   alphaCSR[ 219 ][ 241 ],
   alphaCSR[ 219 ][ 242 ],
   alphaCSR[ 219 ][ 243 ],
   alphaCSR[ 219 ][ 244 ],
   alphaCSR[ 219 ][ 245 ],
   alphaCSR[ 219 ][ 246 ],
   alphaCSR[ 219 ][ 247 ],
   alphaCSR[ 219 ][ 248 ],
   alphaCSR[ 219 ][ 249 ],
   alphaCSR[ 219 ][ 250 ],
   alphaCSR[ 219 ][ 251 ],
   alphaCSR[ 219 ][ 252 ],
   alphaCSR[ 219 ][ 253 ],
   alphaCSR[ 219 ][ 254 ],
   alphaCSR[ 219 ][ 255 ],
   alphaCSR[ 219 ][ 256 ],
   alphaCSR[ 219 ][ 257 ],
   alphaCSR[ 219 ][ 258 ],
   alphaCSR[ 219 ][ 259 ],
   alphaCSR[ 219 ][ 260 ],
   alphaCSR[ 219 ][ 261 ],
   alphaCSR[ 219 ][ 262 ],
   alphaCSR[ 219 ][ 263 ],
   alphaCSR[ 219 ][ 264 ],
   alphaCSR[ 219 ][ 265 ],
   alphaCSR[ 219 ][ 266 ],
   alphaCSR[ 219 ][ 267 ],
   alphaCSR[ 219 ][ 268 ],
   alphaCSR[ 219 ][ 269 ],
   alphaCSR[ 219 ][ 270 ],
   alphaCSR[ 219 ][ 271 ],
   alphaCSR[ 219 ][ 272 ],
   alphaCSR[ 219 ][ 273 ],
   alphaCSR[ 219 ][ 274 ],
   alphaCSR[ 219 ][ 275 ],
   alphaCSR[ 219 ][ 276 ],
   alphaCSR[ 219 ][ 277 ],
   alphaCSR[ 219 ][ 278 ],
   alphaCSR[ 219 ][ 279 ],
   alphaCSR[ 219 ][ 280 ],
   alphaCSR[ 219 ][ 281 ],
   alphaCSR[ 219 ][ 282 ],
   alphaCSR[ 219 ][ 283 ],
   alphaCSR[ 219 ][ 284 ],
   alphaCSR[ 219 ][ 285 ],
   alphaCSR[ 219 ][ 286 ],
   alphaCSR[ 219 ][ 287 ],
   alphaCSR[ 219 ][ 288 ],
   alphaCSR[ 219 ][ 289 ],
   alphaCSR[ 219 ][ 290 ],
   alphaCSR[ 219 ][ 291 ],
   alphaCSR[ 219 ][ 292 ],
   alphaCSR[ 219 ][ 293 ],
   alphaCSR[ 219 ][ 294 ],
   alphaCSR[ 219 ][ 295 ],
   alphaCSR[ 219 ][ 296 ],
   alphaCSR[ 219 ][ 297 ],
   alphaCSR[ 219 ][ 298 ],
   alphaCSR[ 219 ][ 299 ],
   alphaCSR[ 219 ][ 300 ],
   alphaCSR[ 219 ][ 301 ],
   alphaCSR[ 219 ][ 302 ],
   alphaCSR[ 219 ][ 303 ],
   alphaCSR[ 219 ][ 304 ],
   alphaCSR[ 219 ][ 305 ],
   alphaCSR[ 219 ][ 306 ],
   alphaCSR[ 219 ][ 307 ],
   alphaCSR[ 219 ][ 308 ],
   alphaCSR[ 219 ][ 309 ],
   alphaCSR[ 219 ][ 310 ],
   alphaCSR[ 219 ][ 311 ],
   alphaCSR[ 219 ][ 312 ],
   alphaCSR[ 219 ][ 313 ],
   alphaCSR[ 219 ][ 314 ],
   alphaCSR[ 219 ][ 315 ],
   alphaCSR[ 219 ][ 316 ],
   alphaCSR[ 219 ][ 317 ],
   alphaCSR[ 219 ][ 318 ],
   alphaCSR[ 219 ][ 319 ],
   alphaCSR[ 219 ][ 320 ],
   alphaCSR[ 219 ][ 321 ],
   alphaCSR[ 219 ][ 322 ],
   alphaCSR[ 219 ][ 323 ],
   alphaCSR[ 219 ][ 324 ],
   alphaCSR[ 219 ][ 325 ],
   alphaCSR[ 219 ][ 326 ],
   alphaCSR[ 219 ][ 327 ],
   alphaCSR[ 219 ][ 328 ],
   alphaCSR[ 219 ][ 329 ],
   alphaCSR[ 219 ][ 330 ],
   alphaCSR[ 219 ][ 331 ],
   alphaCSR[ 219 ][ 332 ],
   alphaCSR[ 219 ][ 333 ],
   alphaCSR[ 219 ][ 334 ],
   alphaCSR[ 219 ][ 335 ],
   alphaCSR[ 219 ][ 336 ],
   alphaCSR[ 219 ][ 337 ],
   alphaCSR[ 219 ][ 338 ],
   alphaCSR[ 219 ][ 339 ],
   alphaCSR[ 219 ][ 340 ],
   alphaCSR[ 219 ][ 341 ],
   alphaCSR[ 219 ][ 342 ],
   alphaCSR[ 219 ][ 343 ],
   alphaCSR[ 219 ][ 344 ],
   alphaCSR[ 219 ][ 345 ],
   alphaCSR[ 219 ][ 346 ],
   alphaCSR[ 219 ][ 347 ],
   alphaCSR[ 219 ][ 348 ],
   alphaCSR[ 219 ][ 349 ],
   alphaCSR[ 219 ][ 350 ],
   alphaCSR[ 219 ][ 351 ],
   alphaCSR[ 219 ][ 352 ],
   alphaCSR[ 219 ][ 353 ],
   alphaCSR[ 219 ][ 354 ],
   alphaCSR[ 219 ][ 355 ],
   alphaCSR[ 219 ][ 356 ],
   alphaCSR[ 219 ][ 357 ],
   alphaCSR[ 219 ][ 358 ],
   alphaCSR[ 219 ][ 359 ],
   alphaCSR[ 219 ][ 360 ],
   alphaCSR[ 219 ][ 361 ],
   alphaCSR[ 219 ][ 362 ],
   alphaCSR[ 219 ][ 363 ],
   alphaCSR[ 219 ][ 364 ],
   alphaCSR[ 219 ][ 365 ],
   alphaCSR[ 219 ][ 366 ],
   alphaCSR[ 219 ][ 367 ],
   alphaCSR[ 219 ][ 368 ],
   alphaCSR[ 219 ][ 369 ],
   alphaCSR[ 219 ][ 370 ],
   alphaCSR[ 219 ][ 371 ],
   alphaCSR[ 219 ][ 372 ],
   alphaCSR[ 219 ][ 373 ],
   alphaCSR[ 219 ][ 374 ],
   alphaCSR[ 219 ][ 375 ],
   alphaCSR[ 219 ][ 376 ],
   alphaCSR[ 219 ][ 377 ],
   alphaCSR[ 219 ][ 378 ],
   alphaCSR[ 219 ][ 379 ],
   alphaCSR[ 219 ][ 380 ],
   alphaCSR[ 219 ][ 381 ],
   alphaCSR[ 219 ][ 382 ],
   alphaCSR[ 219 ][ 383 ],
   alphaCSR[ 220 ][ 0 ],
   alphaCSR[ 220 ][ 1 ],
   alphaCSR[ 220 ][ 2 ],
   alphaCSR[ 220 ][ 3 ],
   alphaCSR[ 220 ][ 4 ],
   alphaCSR[ 220 ][ 5 ],
   alphaCSR[ 220 ][ 6 ],
   alphaCSR[ 220 ][ 7 ],
   alphaCSR[ 220 ][ 8 ],
   alphaCSR[ 220 ][ 9 ],
   alphaCSR[ 220 ][ 10 ],
   alphaCSR[ 220 ][ 11 ],
   alphaCSR[ 220 ][ 12 ],
   alphaCSR[ 220 ][ 13 ],
   alphaCSR[ 220 ][ 14 ],
   alphaCSR[ 220 ][ 15 ],
   alphaCSR[ 220 ][ 16 ],
   alphaCSR[ 220 ][ 17 ],
   alphaCSR[ 220 ][ 18 ],
   alphaCSR[ 220 ][ 19 ],
   alphaCSR[ 220 ][ 20 ],
   alphaCSR[ 220 ][ 21 ],
   alphaCSR[ 220 ][ 22 ],
   alphaCSR[ 220 ][ 23 ],
   alphaCSR[ 220 ][ 24 ],
   alphaCSR[ 220 ][ 25 ],
   alphaCSR[ 220 ][ 26 ],
   alphaCSR[ 220 ][ 27 ],
   alphaCSR[ 220 ][ 28 ],
   alphaCSR[ 220 ][ 29 ],
   alphaCSR[ 220 ][ 30 ],
   alphaCSR[ 220 ][ 31 ],
   alphaCSR[ 220 ][ 32 ],
   alphaCSR[ 220 ][ 33 ],
   alphaCSR[ 220 ][ 34 ],
   alphaCSR[ 220 ][ 35 ],
   alphaCSR[ 220 ][ 36 ],
   alphaCSR[ 220 ][ 37 ],
   alphaCSR[ 220 ][ 38 ],
   alphaCSR[ 220 ][ 39 ],
   alphaCSR[ 220 ][ 40 ],
   alphaCSR[ 220 ][ 41 ],
   alphaCSR[ 220 ][ 42 ],
   alphaCSR[ 220 ][ 43 ],
   alphaCSR[ 220 ][ 44 ],
   alphaCSR[ 220 ][ 45 ],
   alphaCSR[ 220 ][ 46 ],
   alphaCSR[ 220 ][ 47 ],
   alphaCSR[ 220 ][ 48 ],
   alphaCSR[ 220 ][ 49 ],
   alphaCSR[ 220 ][ 50 ],
   alphaCSR[ 220 ][ 51 ],
   alphaCSR[ 220 ][ 52 ],
   alphaCSR[ 220 ][ 53 ],
   alphaCSR[ 220 ][ 54 ],
   alphaCSR[ 220 ][ 55 ],
   alphaCSR[ 220 ][ 56 ],
   alphaCSR[ 220 ][ 57 ],
   alphaCSR[ 220 ][ 58 ],
   alphaCSR[ 220 ][ 59 ],
   alphaCSR[ 220 ][ 60 ],
   alphaCSR[ 220 ][ 61 ],
   alphaCSR[ 220 ][ 62 ],
   alphaCSR[ 220 ][ 63 ],
   alphaCSR[ 220 ][ 64 ],
   alphaCSR[ 220 ][ 65 ],
   alphaCSR[ 220 ][ 66 ],
   alphaCSR[ 220 ][ 67 ],
   alphaCSR[ 220 ][ 68 ],
   alphaCSR[ 220 ][ 69 ],
   alphaCSR[ 220 ][ 70 ],
   alphaCSR[ 220 ][ 71 ],
   alphaCSR[ 220 ][ 72 ],
   alphaCSR[ 220 ][ 73 ],
   alphaCSR[ 220 ][ 74 ],
   alphaCSR[ 220 ][ 75 ],
   alphaCSR[ 220 ][ 76 ],
   alphaCSR[ 220 ][ 77 ],
   alphaCSR[ 220 ][ 78 ],
   alphaCSR[ 220 ][ 79 ],
   alphaCSR[ 220 ][ 80 ],
   alphaCSR[ 220 ][ 81 ],
   alphaCSR[ 220 ][ 82 ],
   alphaCSR[ 220 ][ 83 ],
   alphaCSR[ 220 ][ 84 ],
   alphaCSR[ 220 ][ 85 ],
   alphaCSR[ 220 ][ 86 ],
   alphaCSR[ 220 ][ 87 ],
   alphaCSR[ 220 ][ 88 ],
   alphaCSR[ 220 ][ 89 ],
   alphaCSR[ 220 ][ 90 ],
   alphaCSR[ 220 ][ 91 ],
   alphaCSR[ 220 ][ 92 ],
   alphaCSR[ 220 ][ 93 ],
   alphaCSR[ 220 ][ 94 ],
   alphaCSR[ 220 ][ 95 ],
   alphaCSR[ 220 ][ 96 ],
   alphaCSR[ 220 ][ 97 ],
   alphaCSR[ 220 ][ 98 ],
   alphaCSR[ 220 ][ 99 ],
   alphaCSR[ 220 ][ 100 ],
   alphaCSR[ 220 ][ 101 ],
   alphaCSR[ 220 ][ 102 ],
   alphaCSR[ 220 ][ 103 ],
   alphaCSR[ 220 ][ 104 ],
   alphaCSR[ 220 ][ 105 ],
   alphaCSR[ 220 ][ 106 ],
   alphaCSR[ 220 ][ 107 ],
   alphaCSR[ 220 ][ 108 ],
   alphaCSR[ 220 ][ 109 ],
   alphaCSR[ 220 ][ 110 ],
   alphaCSR[ 220 ][ 111 ],
   alphaCSR[ 220 ][ 112 ],
   alphaCSR[ 220 ][ 113 ],
   alphaCSR[ 220 ][ 114 ],
   alphaCSR[ 220 ][ 115 ],
   alphaCSR[ 220 ][ 116 ],
   alphaCSR[ 220 ][ 117 ],
   alphaCSR[ 220 ][ 118 ],
   alphaCSR[ 220 ][ 119 ],
   alphaCSR[ 220 ][ 120 ],
   alphaCSR[ 220 ][ 121 ],
   alphaCSR[ 220 ][ 122 ],
   alphaCSR[ 220 ][ 123 ],
   alphaCSR[ 220 ][ 124 ],
   alphaCSR[ 220 ][ 125 ],
   alphaCSR[ 220 ][ 126 ],
   alphaCSR[ 220 ][ 127 ],
   alphaCSR[ 220 ][ 128 ],
   alphaCSR[ 220 ][ 129 ],
   alphaCSR[ 220 ][ 130 ],
   alphaCSR[ 220 ][ 131 ],
   alphaCSR[ 220 ][ 132 ],
   alphaCSR[ 220 ][ 133 ],
   alphaCSR[ 220 ][ 134 ],
   alphaCSR[ 220 ][ 135 ],
   alphaCSR[ 220 ][ 136 ],
   alphaCSR[ 220 ][ 137 ],
   alphaCSR[ 220 ][ 138 ],
   alphaCSR[ 220 ][ 139 ],
   alphaCSR[ 220 ][ 140 ],
   alphaCSR[ 220 ][ 141 ],
   alphaCSR[ 220 ][ 142 ],
   alphaCSR[ 220 ][ 143 ],
   alphaCSR[ 220 ][ 144 ],
   alphaCSR[ 220 ][ 145 ],
   alphaCSR[ 220 ][ 146 ],
   alphaCSR[ 220 ][ 147 ],
   alphaCSR[ 220 ][ 148 ],
   alphaCSR[ 220 ][ 149 ],
   alphaCSR[ 220 ][ 150 ],
   alphaCSR[ 220 ][ 151 ],
   alphaCSR[ 220 ][ 152 ],
   alphaCSR[ 220 ][ 153 ],
   alphaCSR[ 220 ][ 154 ],
   alphaCSR[ 220 ][ 155 ],
   alphaCSR[ 220 ][ 156 ],
   alphaCSR[ 220 ][ 157 ],
   alphaCSR[ 220 ][ 158 ],
   alphaCSR[ 220 ][ 159 ],
   alphaCSR[ 220 ][ 160 ],
   alphaCSR[ 220 ][ 161 ],
   alphaCSR[ 220 ][ 162 ],
   alphaCSR[ 220 ][ 163 ],
   alphaCSR[ 220 ][ 164 ],
   alphaCSR[ 220 ][ 165 ],
   alphaCSR[ 220 ][ 166 ],
   alphaCSR[ 220 ][ 167 ],
   alphaCSR[ 220 ][ 168 ],
   alphaCSR[ 220 ][ 169 ],
   alphaCSR[ 220 ][ 170 ],
   alphaCSR[ 220 ][ 171 ],
   alphaCSR[ 220 ][ 172 ],
   alphaCSR[ 220 ][ 173 ],
   alphaCSR[ 220 ][ 174 ],
   alphaCSR[ 220 ][ 175 ],
   alphaCSR[ 220 ][ 176 ],
   alphaCSR[ 220 ][ 177 ],
   alphaCSR[ 220 ][ 178 ],
   alphaCSR[ 220 ][ 179 ],
   alphaCSR[ 220 ][ 180 ],
   alphaCSR[ 220 ][ 181 ],
   alphaCSR[ 220 ][ 182 ],
   alphaCSR[ 220 ][ 183 ],
   alphaCSR[ 220 ][ 184 ],
   alphaCSR[ 220 ][ 185 ],
   alphaCSR[ 220 ][ 186 ],
   alphaCSR[ 220 ][ 187 ],
   alphaCSR[ 220 ][ 188 ],
   alphaCSR[ 220 ][ 189 ],
   alphaCSR[ 220 ][ 190 ],
   alphaCSR[ 220 ][ 191 ],
   alphaCSR[ 220 ][ 192 ],
   alphaCSR[ 220 ][ 193 ],
   alphaCSR[ 220 ][ 194 ],
   alphaCSR[ 220 ][ 195 ],
   alphaCSR[ 220 ][ 196 ],
   alphaCSR[ 220 ][ 197 ],
   alphaCSR[ 220 ][ 198 ],
   alphaCSR[ 220 ][ 199 ],
   alphaCSR[ 220 ][ 200 ],
   alphaCSR[ 220 ][ 201 ],
   alphaCSR[ 220 ][ 202 ],
   alphaCSR[ 220 ][ 203 ],
   alphaCSR[ 220 ][ 204 ],
   alphaCSR[ 220 ][ 205 ],
   alphaCSR[ 220 ][ 206 ],
   alphaCSR[ 220 ][ 207 ],
   alphaCSR[ 220 ][ 208 ],
   alphaCSR[ 220 ][ 209 ],
   alphaCSR[ 220 ][ 210 ],
   alphaCSR[ 220 ][ 211 ],
   alphaCSR[ 220 ][ 212 ],
   alphaCSR[ 220 ][ 213 ],
   alphaCSR[ 220 ][ 214 ],
   alphaCSR[ 220 ][ 215 ],
   alphaCSR[ 220 ][ 216 ],
   alphaCSR[ 220 ][ 217 ],
   alphaCSR[ 220 ][ 218 ],
   alphaCSR[ 220 ][ 219 ],
   alphaCSR[ 220 ][ 220 ],
   alphaCSR[ 220 ][ 221 ],
   alphaCSR[ 220 ][ 222 ],
   alphaCSR[ 220 ][ 223 ],
   alphaCSR[ 220 ][ 224 ],
   alphaCSR[ 220 ][ 225 ],
   alphaCSR[ 220 ][ 226 ],
   alphaCSR[ 220 ][ 227 ],
   alphaCSR[ 220 ][ 228 ],
   alphaCSR[ 220 ][ 229 ],
   alphaCSR[ 220 ][ 230 ],
   alphaCSR[ 220 ][ 231 ],
   alphaCSR[ 220 ][ 232 ],
   alphaCSR[ 220 ][ 233 ],
   alphaCSR[ 220 ][ 234 ],
   alphaCSR[ 220 ][ 235 ],
   alphaCSR[ 220 ][ 236 ],
   alphaCSR[ 220 ][ 237 ],
   alphaCSR[ 220 ][ 238 ],
   alphaCSR[ 220 ][ 239 ],
   alphaCSR[ 220 ][ 240 ],
   alphaCSR[ 220 ][ 241 ],
   alphaCSR[ 220 ][ 242 ],
   alphaCSR[ 220 ][ 243 ],
   alphaCSR[ 220 ][ 244 ],
   alphaCSR[ 220 ][ 245 ],
   alphaCSR[ 220 ][ 246 ],
   alphaCSR[ 220 ][ 247 ],
   alphaCSR[ 220 ][ 248 ],
   alphaCSR[ 220 ][ 249 ],
   alphaCSR[ 220 ][ 250 ],
   alphaCSR[ 220 ][ 251 ],
   alphaCSR[ 220 ][ 252 ],
   alphaCSR[ 220 ][ 253 ],
   alphaCSR[ 220 ][ 254 ],
   alphaCSR[ 220 ][ 255 ],
   alphaCSR[ 220 ][ 256 ],
   alphaCSR[ 220 ][ 257 ],
   alphaCSR[ 220 ][ 258 ],
   alphaCSR[ 220 ][ 259 ],
   alphaCSR[ 220 ][ 260 ],
   alphaCSR[ 220 ][ 261 ],
   alphaCSR[ 220 ][ 262 ],
   alphaCSR[ 220 ][ 263 ],
   alphaCSR[ 220 ][ 264 ],
   alphaCSR[ 220 ][ 265 ],
   alphaCSR[ 220 ][ 266 ],
   alphaCSR[ 220 ][ 267 ],
   alphaCSR[ 220 ][ 268 ],
   alphaCSR[ 220 ][ 269 ],
   alphaCSR[ 220 ][ 270 ],
   alphaCSR[ 220 ][ 271 ],
   alphaCSR[ 220 ][ 272 ],
   alphaCSR[ 220 ][ 273 ],
   alphaCSR[ 220 ][ 274 ],
   alphaCSR[ 220 ][ 275 ],
   alphaCSR[ 220 ][ 276 ],
   alphaCSR[ 220 ][ 277 ],
   alphaCSR[ 220 ][ 278 ],
   alphaCSR[ 220 ][ 279 ],
   alphaCSR[ 220 ][ 280 ],
   alphaCSR[ 220 ][ 281 ],
   alphaCSR[ 220 ][ 282 ],
   alphaCSR[ 220 ][ 283 ],
   alphaCSR[ 220 ][ 284 ],
   alphaCSR[ 220 ][ 285 ],
   alphaCSR[ 220 ][ 286 ],
   alphaCSR[ 220 ][ 287 ],
   alphaCSR[ 220 ][ 288 ],
   alphaCSR[ 220 ][ 289 ],
   alphaCSR[ 220 ][ 290 ],
   alphaCSR[ 220 ][ 291 ],
   alphaCSR[ 220 ][ 292 ],
   alphaCSR[ 220 ][ 293 ],
   alphaCSR[ 220 ][ 294 ],
   alphaCSR[ 220 ][ 295 ],
   alphaCSR[ 220 ][ 296 ],
   alphaCSR[ 220 ][ 297 ],
   alphaCSR[ 220 ][ 298 ],
   alphaCSR[ 220 ][ 299 ],
   alphaCSR[ 220 ][ 300 ],
   alphaCSR[ 220 ][ 301 ],
   alphaCSR[ 220 ][ 302 ],
   alphaCSR[ 220 ][ 303 ],
   alphaCSR[ 220 ][ 304 ],
   alphaCSR[ 220 ][ 305 ],
   alphaCSR[ 220 ][ 306 ],
   alphaCSR[ 220 ][ 307 ],
   alphaCSR[ 220 ][ 308 ],
   alphaCSR[ 220 ][ 309 ],
   alphaCSR[ 220 ][ 310 ],
   alphaCSR[ 220 ][ 311 ],
   alphaCSR[ 220 ][ 312 ],
   alphaCSR[ 220 ][ 313 ],
   alphaCSR[ 220 ][ 314 ],
   alphaCSR[ 220 ][ 315 ],
   alphaCSR[ 220 ][ 316 ],
   alphaCSR[ 220 ][ 317 ],
   alphaCSR[ 220 ][ 318 ],
   alphaCSR[ 220 ][ 319 ],
   alphaCSR[ 220 ][ 320 ],
   alphaCSR[ 220 ][ 321 ],
   alphaCSR[ 220 ][ 322 ],
   alphaCSR[ 220 ][ 323 ],
   alphaCSR[ 220 ][ 324 ],
   alphaCSR[ 220 ][ 325 ],
   alphaCSR[ 220 ][ 326 ],
   alphaCSR[ 220 ][ 327 ],
   alphaCSR[ 220 ][ 328 ],
   alphaCSR[ 220 ][ 329 ],
   alphaCSR[ 220 ][ 330 ],
   alphaCSR[ 220 ][ 331 ],
   alphaCSR[ 220 ][ 332 ],
   alphaCSR[ 220 ][ 333 ],
   alphaCSR[ 220 ][ 334 ],
   alphaCSR[ 220 ][ 335 ],
   alphaCSR[ 220 ][ 336 ],
   alphaCSR[ 220 ][ 337 ],
   alphaCSR[ 220 ][ 338 ],
   alphaCSR[ 220 ][ 339 ],
   alphaCSR[ 220 ][ 340 ],
   alphaCSR[ 220 ][ 341 ],
   alphaCSR[ 220 ][ 342 ],
   alphaCSR[ 220 ][ 343 ],
   alphaCSR[ 220 ][ 344 ],
   alphaCSR[ 220 ][ 345 ],
   alphaCSR[ 220 ][ 346 ],
   alphaCSR[ 220 ][ 347 ],
   alphaCSR[ 220 ][ 348 ],
   alphaCSR[ 220 ][ 349 ],
   alphaCSR[ 220 ][ 350 ],
   alphaCSR[ 220 ][ 351 ],
   alphaCSR[ 220 ][ 352 ],
   alphaCSR[ 220 ][ 353 ],
   alphaCSR[ 220 ][ 354 ],
   alphaCSR[ 220 ][ 355 ],
   alphaCSR[ 220 ][ 356 ],
   alphaCSR[ 220 ][ 357 ],
   alphaCSR[ 220 ][ 358 ],
   alphaCSR[ 220 ][ 359 ],
   alphaCSR[ 220 ][ 360 ],
   alphaCSR[ 220 ][ 361 ],
   alphaCSR[ 220 ][ 362 ],
   alphaCSR[ 220 ][ 363 ],
   alphaCSR[ 220 ][ 364 ],
   alphaCSR[ 220 ][ 365 ],
   alphaCSR[ 220 ][ 366 ],
   alphaCSR[ 220 ][ 367 ],
   alphaCSR[ 220 ][ 368 ],
   alphaCSR[ 220 ][ 369 ],
   alphaCSR[ 220 ][ 370 ],
   alphaCSR[ 220 ][ 371 ],
   alphaCSR[ 220 ][ 372 ],
   alphaCSR[ 220 ][ 373 ],
   alphaCSR[ 220 ][ 374 ],
   alphaCSR[ 220 ][ 375 ],
   alphaCSR[ 220 ][ 376 ],
   alphaCSR[ 220 ][ 377 ],
   alphaCSR[ 220 ][ 378 ],
   alphaCSR[ 220 ][ 379 ],
   alphaCSR[ 220 ][ 380 ],
   alphaCSR[ 220 ][ 381 ],
   alphaCSR[ 220 ][ 382 ],
   alphaCSR[ 220 ][ 383 ],
   alphaCSR[ 221 ][ 0 ],
   alphaCSR[ 221 ][ 1 ],
   alphaCSR[ 221 ][ 2 ],
   alphaCSR[ 221 ][ 3 ],
   alphaCSR[ 221 ][ 4 ],
   alphaCSR[ 221 ][ 5 ],
   alphaCSR[ 221 ][ 6 ],
   alphaCSR[ 221 ][ 7 ],
   alphaCSR[ 221 ][ 8 ],
   alphaCSR[ 221 ][ 9 ],
   alphaCSR[ 221 ][ 10 ],
   alphaCSR[ 221 ][ 11 ],
   alphaCSR[ 221 ][ 12 ],
   alphaCSR[ 221 ][ 13 ],
   alphaCSR[ 221 ][ 14 ],
   alphaCSR[ 221 ][ 15 ],
   alphaCSR[ 221 ][ 16 ],
   alphaCSR[ 221 ][ 17 ],
   alphaCSR[ 221 ][ 18 ],
   alphaCSR[ 221 ][ 19 ],
   alphaCSR[ 221 ][ 20 ],
   alphaCSR[ 221 ][ 21 ],
   alphaCSR[ 221 ][ 22 ],
   alphaCSR[ 221 ][ 23 ],
   alphaCSR[ 221 ][ 24 ],
   alphaCSR[ 221 ][ 25 ],
   alphaCSR[ 221 ][ 26 ],
   alphaCSR[ 221 ][ 27 ],
   alphaCSR[ 221 ][ 28 ],
   alphaCSR[ 221 ][ 29 ],
   alphaCSR[ 221 ][ 30 ],
   alphaCSR[ 221 ][ 31 ],
   alphaCSR[ 221 ][ 32 ],
   alphaCSR[ 221 ][ 33 ],
   alphaCSR[ 221 ][ 34 ],
   alphaCSR[ 221 ][ 35 ],
   alphaCSR[ 221 ][ 36 ],
   alphaCSR[ 221 ][ 37 ],
   alphaCSR[ 221 ][ 38 ],
   alphaCSR[ 221 ][ 39 ],
   alphaCSR[ 221 ][ 40 ],
   alphaCSR[ 221 ][ 41 ],
   alphaCSR[ 221 ][ 42 ],
   alphaCSR[ 221 ][ 43 ],
   alphaCSR[ 221 ][ 44 ],
   alphaCSR[ 221 ][ 45 ],
   alphaCSR[ 221 ][ 46 ],
   alphaCSR[ 221 ][ 47 ],
   alphaCSR[ 221 ][ 48 ],
   alphaCSR[ 221 ][ 49 ],
   alphaCSR[ 221 ][ 50 ],
   alphaCSR[ 221 ][ 51 ],
   alphaCSR[ 221 ][ 52 ],
   alphaCSR[ 221 ][ 53 ],
   alphaCSR[ 221 ][ 54 ],
   alphaCSR[ 221 ][ 55 ],
   alphaCSR[ 221 ][ 56 ],
   alphaCSR[ 221 ][ 57 ],
   alphaCSR[ 221 ][ 58 ],
   alphaCSR[ 221 ][ 59 ],
   alphaCSR[ 221 ][ 60 ],
   alphaCSR[ 221 ][ 61 ],
   alphaCSR[ 221 ][ 62 ],
   alphaCSR[ 221 ][ 63 ],
   alphaCSR[ 221 ][ 64 ],
   alphaCSR[ 221 ][ 65 ],
   alphaCSR[ 221 ][ 66 ],
   alphaCSR[ 221 ][ 67 ],
   alphaCSR[ 221 ][ 68 ],
   alphaCSR[ 221 ][ 69 ],
   alphaCSR[ 221 ][ 70 ],
   alphaCSR[ 221 ][ 71 ],
   alphaCSR[ 221 ][ 72 ],
   alphaCSR[ 221 ][ 73 ],
   alphaCSR[ 221 ][ 74 ],
   alphaCSR[ 221 ][ 75 ],
   alphaCSR[ 221 ][ 76 ],
   alphaCSR[ 221 ][ 77 ],
   alphaCSR[ 221 ][ 78 ],
   alphaCSR[ 221 ][ 79 ],
   alphaCSR[ 221 ][ 80 ],
   alphaCSR[ 221 ][ 81 ],
   alphaCSR[ 221 ][ 82 ],
   alphaCSR[ 221 ][ 83 ],
   alphaCSR[ 221 ][ 84 ],
   alphaCSR[ 221 ][ 85 ],
   alphaCSR[ 221 ][ 86 ],
   alphaCSR[ 221 ][ 87 ],
   alphaCSR[ 221 ][ 88 ],
   alphaCSR[ 221 ][ 89 ],
   alphaCSR[ 221 ][ 90 ],
   alphaCSR[ 221 ][ 91 ],
   alphaCSR[ 221 ][ 92 ],
   alphaCSR[ 221 ][ 93 ],
   alphaCSR[ 221 ][ 94 ],
   alphaCSR[ 221 ][ 95 ],
   alphaCSR[ 221 ][ 96 ],
   alphaCSR[ 221 ][ 97 ],
   alphaCSR[ 221 ][ 98 ],
   alphaCSR[ 221 ][ 99 ],
   alphaCSR[ 221 ][ 100 ],
   alphaCSR[ 221 ][ 101 ],
   alphaCSR[ 221 ][ 102 ],
   alphaCSR[ 221 ][ 103 ],
   alphaCSR[ 221 ][ 104 ],
   alphaCSR[ 221 ][ 105 ],
   alphaCSR[ 221 ][ 106 ],
   alphaCSR[ 221 ][ 107 ],
   alphaCSR[ 221 ][ 108 ],
   alphaCSR[ 221 ][ 109 ],
   alphaCSR[ 221 ][ 110 ],
   alphaCSR[ 221 ][ 111 ],
   alphaCSR[ 221 ][ 112 ],
   alphaCSR[ 221 ][ 113 ],
   alphaCSR[ 221 ][ 114 ],
   alphaCSR[ 221 ][ 115 ],
   alphaCSR[ 221 ][ 116 ],
   alphaCSR[ 221 ][ 117 ],
   alphaCSR[ 221 ][ 118 ],
   alphaCSR[ 221 ][ 119 ],
   alphaCSR[ 221 ][ 120 ],
   alphaCSR[ 221 ][ 121 ],
   alphaCSR[ 221 ][ 122 ],
   alphaCSR[ 221 ][ 123 ],
   alphaCSR[ 221 ][ 124 ],
   alphaCSR[ 221 ][ 125 ],
   alphaCSR[ 221 ][ 126 ],
   alphaCSR[ 221 ][ 127 ],
   alphaCSR[ 221 ][ 128 ],
   alphaCSR[ 221 ][ 129 ],
   alphaCSR[ 221 ][ 130 ],
   alphaCSR[ 221 ][ 131 ],
   alphaCSR[ 221 ][ 132 ],
   alphaCSR[ 221 ][ 133 ],
   alphaCSR[ 221 ][ 134 ],
   alphaCSR[ 221 ][ 135 ],
   alphaCSR[ 221 ][ 136 ],
   alphaCSR[ 221 ][ 137 ],
   alphaCSR[ 221 ][ 138 ],
   alphaCSR[ 221 ][ 139 ],
   alphaCSR[ 221 ][ 140 ],
   alphaCSR[ 221 ][ 141 ],
   alphaCSR[ 221 ][ 142 ],
   alphaCSR[ 221 ][ 143 ],
   alphaCSR[ 221 ][ 144 ],
   alphaCSR[ 221 ][ 145 ],
   alphaCSR[ 221 ][ 146 ],
   alphaCSR[ 221 ][ 147 ],
   alphaCSR[ 221 ][ 148 ],
   alphaCSR[ 221 ][ 149 ],
   alphaCSR[ 221 ][ 150 ],
   alphaCSR[ 221 ][ 151 ],
   alphaCSR[ 221 ][ 152 ],
   alphaCSR[ 221 ][ 153 ],
   alphaCSR[ 221 ][ 154 ],
   alphaCSR[ 221 ][ 155 ],
   alphaCSR[ 221 ][ 156 ],
   alphaCSR[ 221 ][ 157 ],
   alphaCSR[ 221 ][ 158 ],
   alphaCSR[ 221 ][ 159 ],
   alphaCSR[ 221 ][ 160 ],
   alphaCSR[ 221 ][ 161 ],
   alphaCSR[ 221 ][ 162 ],
   alphaCSR[ 221 ][ 163 ],
   alphaCSR[ 221 ][ 164 ],
   alphaCSR[ 221 ][ 165 ],
   alphaCSR[ 221 ][ 166 ],
   alphaCSR[ 221 ][ 167 ],
   alphaCSR[ 221 ][ 168 ],
   alphaCSR[ 221 ][ 169 ],
   alphaCSR[ 221 ][ 170 ],
   alphaCSR[ 221 ][ 171 ],
   alphaCSR[ 221 ][ 172 ],
   alphaCSR[ 221 ][ 173 ],
   alphaCSR[ 221 ][ 174 ],
   alphaCSR[ 221 ][ 175 ],
   alphaCSR[ 221 ][ 176 ],
   alphaCSR[ 221 ][ 177 ],
   alphaCSR[ 221 ][ 178 ],
   alphaCSR[ 221 ][ 179 ],
   alphaCSR[ 221 ][ 180 ],
   alphaCSR[ 221 ][ 181 ],
   alphaCSR[ 221 ][ 182 ],
   alphaCSR[ 221 ][ 183 ],
   alphaCSR[ 221 ][ 184 ],
   alphaCSR[ 221 ][ 185 ],
   alphaCSR[ 221 ][ 186 ],
   alphaCSR[ 221 ][ 187 ],
   alphaCSR[ 221 ][ 188 ],
   alphaCSR[ 221 ][ 189 ],
   alphaCSR[ 221 ][ 190 ],
   alphaCSR[ 221 ][ 191 ],
   alphaCSR[ 221 ][ 192 ],
   alphaCSR[ 221 ][ 193 ],
   alphaCSR[ 221 ][ 194 ],
   alphaCSR[ 221 ][ 195 ],
   alphaCSR[ 221 ][ 196 ],
   alphaCSR[ 221 ][ 197 ],
   alphaCSR[ 221 ][ 198 ],
   alphaCSR[ 221 ][ 199 ],
   alphaCSR[ 221 ][ 200 ],
   alphaCSR[ 221 ][ 201 ],
   alphaCSR[ 221 ][ 202 ],
   alphaCSR[ 221 ][ 203 ],
   alphaCSR[ 221 ][ 204 ],
   alphaCSR[ 221 ][ 205 ],
   alphaCSR[ 221 ][ 206 ],
   alphaCSR[ 221 ][ 207 ],
   alphaCSR[ 221 ][ 208 ],
   alphaCSR[ 221 ][ 209 ],
   alphaCSR[ 221 ][ 210 ],
   alphaCSR[ 221 ][ 211 ],
   alphaCSR[ 221 ][ 212 ],
   alphaCSR[ 221 ][ 213 ],
   alphaCSR[ 221 ][ 214 ],
   alphaCSR[ 221 ][ 215 ],
   alphaCSR[ 221 ][ 216 ],
   alphaCSR[ 221 ][ 217 ],
   alphaCSR[ 221 ][ 218 ],
   alphaCSR[ 221 ][ 219 ],
   alphaCSR[ 221 ][ 220 ],
   alphaCSR[ 221 ][ 221 ],
   alphaCSR[ 221 ][ 222 ],
   alphaCSR[ 221 ][ 223 ],
   alphaCSR[ 221 ][ 224 ],
   alphaCSR[ 221 ][ 225 ],
   alphaCSR[ 221 ][ 226 ],
   alphaCSR[ 221 ][ 227 ],
   alphaCSR[ 221 ][ 228 ],
   alphaCSR[ 221 ][ 229 ],
   alphaCSR[ 221 ][ 230 ],
   alphaCSR[ 221 ][ 231 ],
   alphaCSR[ 221 ][ 232 ],
   alphaCSR[ 221 ][ 233 ],
   alphaCSR[ 221 ][ 234 ],
   alphaCSR[ 221 ][ 235 ],
   alphaCSR[ 221 ][ 236 ],
   alphaCSR[ 221 ][ 237 ],
   alphaCSR[ 221 ][ 238 ],
   alphaCSR[ 221 ][ 239 ],
   alphaCSR[ 221 ][ 240 ],
   alphaCSR[ 221 ][ 241 ],
   alphaCSR[ 221 ][ 242 ],
   alphaCSR[ 221 ][ 243 ],
   alphaCSR[ 221 ][ 244 ],
   alphaCSR[ 221 ][ 245 ],
   alphaCSR[ 221 ][ 246 ],
   alphaCSR[ 221 ][ 247 ],
   alphaCSR[ 221 ][ 248 ],
   alphaCSR[ 221 ][ 249 ],
   alphaCSR[ 221 ][ 250 ],
   alphaCSR[ 221 ][ 251 ],
   alphaCSR[ 221 ][ 252 ],
   alphaCSR[ 221 ][ 253 ],
   alphaCSR[ 221 ][ 254 ],
   alphaCSR[ 221 ][ 255 ],
   alphaCSR[ 221 ][ 256 ],
   alphaCSR[ 221 ][ 257 ],
   alphaCSR[ 221 ][ 258 ],
   alphaCSR[ 221 ][ 259 ],
   alphaCSR[ 221 ][ 260 ],
   alphaCSR[ 221 ][ 261 ],
   alphaCSR[ 221 ][ 262 ],
   alphaCSR[ 221 ][ 263 ],
   alphaCSR[ 221 ][ 264 ],
   alphaCSR[ 221 ][ 265 ],
   alphaCSR[ 221 ][ 266 ],
   alphaCSR[ 221 ][ 267 ],
   alphaCSR[ 221 ][ 268 ],
   alphaCSR[ 221 ][ 269 ],
   alphaCSR[ 221 ][ 270 ],
   alphaCSR[ 221 ][ 271 ],
   alphaCSR[ 221 ][ 272 ],
   alphaCSR[ 221 ][ 273 ],
   alphaCSR[ 221 ][ 274 ],
   alphaCSR[ 221 ][ 275 ],
   alphaCSR[ 221 ][ 276 ],
   alphaCSR[ 221 ][ 277 ],
   alphaCSR[ 221 ][ 278 ],
   alphaCSR[ 221 ][ 279 ],
   alphaCSR[ 221 ][ 280 ],
   alphaCSR[ 221 ][ 281 ],
   alphaCSR[ 221 ][ 282 ],
   alphaCSR[ 221 ][ 283 ],
   alphaCSR[ 221 ][ 284 ],
   alphaCSR[ 221 ][ 285 ],
   alphaCSR[ 221 ][ 286 ],
   alphaCSR[ 221 ][ 287 ],
   alphaCSR[ 221 ][ 288 ],
   alphaCSR[ 221 ][ 289 ],
   alphaCSR[ 221 ][ 290 ],
   alphaCSR[ 221 ][ 291 ],
   alphaCSR[ 221 ][ 292 ],
   alphaCSR[ 221 ][ 293 ],
   alphaCSR[ 221 ][ 294 ],
   alphaCSR[ 221 ][ 295 ],
   alphaCSR[ 221 ][ 296 ],
   alphaCSR[ 221 ][ 297 ],
   alphaCSR[ 221 ][ 298 ],
   alphaCSR[ 221 ][ 299 ],
   alphaCSR[ 221 ][ 300 ],
   alphaCSR[ 221 ][ 301 ],
   alphaCSR[ 221 ][ 302 ],
   alphaCSR[ 221 ][ 303 ],
   alphaCSR[ 221 ][ 304 ],
   alphaCSR[ 221 ][ 305 ],
   alphaCSR[ 221 ][ 306 ],
   alphaCSR[ 221 ][ 307 ],
   alphaCSR[ 221 ][ 308 ],
   alphaCSR[ 221 ][ 309 ],
   alphaCSR[ 221 ][ 310 ],
   alphaCSR[ 221 ][ 311 ],
   alphaCSR[ 221 ][ 312 ],
   alphaCSR[ 221 ][ 313 ],
   alphaCSR[ 221 ][ 314 ],
   alphaCSR[ 221 ][ 315 ],
   alphaCSR[ 221 ][ 316 ],
   alphaCSR[ 221 ][ 317 ],
   alphaCSR[ 221 ][ 318 ],
   alphaCSR[ 221 ][ 319 ],
   alphaCSR[ 221 ][ 320 ],
   alphaCSR[ 221 ][ 321 ],
   alphaCSR[ 221 ][ 322 ],
   alphaCSR[ 221 ][ 323 ],
   alphaCSR[ 221 ][ 324 ],
   alphaCSR[ 221 ][ 325 ],
   alphaCSR[ 221 ][ 326 ],
   alphaCSR[ 221 ][ 327 ],
   alphaCSR[ 221 ][ 328 ],
   alphaCSR[ 221 ][ 329 ],
   alphaCSR[ 221 ][ 330 ],
   alphaCSR[ 221 ][ 331 ],
   alphaCSR[ 221 ][ 332 ],
   alphaCSR[ 221 ][ 333 ],
   alphaCSR[ 221 ][ 334 ],
   alphaCSR[ 221 ][ 335 ],
   alphaCSR[ 221 ][ 336 ],
   alphaCSR[ 221 ][ 337 ],
   alphaCSR[ 221 ][ 338 ],
   alphaCSR[ 221 ][ 339 ],
   alphaCSR[ 221 ][ 340 ],
   alphaCSR[ 221 ][ 341 ],
   alphaCSR[ 221 ][ 342 ],
   alphaCSR[ 221 ][ 343 ],
   alphaCSR[ 221 ][ 344 ],
   alphaCSR[ 221 ][ 345 ],
   alphaCSR[ 221 ][ 346 ],
   alphaCSR[ 221 ][ 347 ],
   alphaCSR[ 221 ][ 348 ],
   alphaCSR[ 221 ][ 349 ],
   alphaCSR[ 221 ][ 350 ],
   alphaCSR[ 221 ][ 351 ],
   alphaCSR[ 221 ][ 352 ],
   alphaCSR[ 221 ][ 353 ],
   alphaCSR[ 221 ][ 354 ],
   alphaCSR[ 221 ][ 355 ],
   alphaCSR[ 221 ][ 356 ],
   alphaCSR[ 221 ][ 357 ],
   alphaCSR[ 221 ][ 358 ],
   alphaCSR[ 221 ][ 359 ],
   alphaCSR[ 221 ][ 360 ],
   alphaCSR[ 221 ][ 361 ],
   alphaCSR[ 221 ][ 362 ],
   alphaCSR[ 221 ][ 363 ],
   alphaCSR[ 221 ][ 364 ],
   alphaCSR[ 221 ][ 365 ],
   alphaCSR[ 221 ][ 366 ],
   alphaCSR[ 221 ][ 367 ],
   alphaCSR[ 221 ][ 368 ],
   alphaCSR[ 221 ][ 369 ],
   alphaCSR[ 221 ][ 370 ],
   alphaCSR[ 221 ][ 371 ],
   alphaCSR[ 221 ][ 372 ],
   alphaCSR[ 221 ][ 373 ],
   alphaCSR[ 221 ][ 374 ],
   alphaCSR[ 221 ][ 375 ],
   alphaCSR[ 221 ][ 376 ],
   alphaCSR[ 221 ][ 377 ],
   alphaCSR[ 221 ][ 378 ],
   alphaCSR[ 221 ][ 379 ],
   alphaCSR[ 221 ][ 380 ],
   alphaCSR[ 221 ][ 381 ],
   alphaCSR[ 221 ][ 382 ],
   alphaCSR[ 221 ][ 383 ],
   alphaCSR[ 222 ][ 0 ],
   alphaCSR[ 222 ][ 1 ],
   alphaCSR[ 222 ][ 2 ],
   alphaCSR[ 222 ][ 3 ],
   alphaCSR[ 222 ][ 4 ],
   alphaCSR[ 222 ][ 5 ],
   alphaCSR[ 222 ][ 6 ],
   alphaCSR[ 222 ][ 7 ],
   alphaCSR[ 222 ][ 8 ],
   alphaCSR[ 222 ][ 9 ],
   alphaCSR[ 222 ][ 10 ],
   alphaCSR[ 222 ][ 11 ],
   alphaCSR[ 222 ][ 12 ],
   alphaCSR[ 222 ][ 13 ],
   alphaCSR[ 222 ][ 14 ],
   alphaCSR[ 222 ][ 15 ],
   alphaCSR[ 222 ][ 16 ],
   alphaCSR[ 222 ][ 17 ],
   alphaCSR[ 222 ][ 18 ],
   alphaCSR[ 222 ][ 19 ],
   alphaCSR[ 222 ][ 20 ],
   alphaCSR[ 222 ][ 21 ],
   alphaCSR[ 222 ][ 22 ],
   alphaCSR[ 222 ][ 23 ],
   alphaCSR[ 222 ][ 24 ],
   alphaCSR[ 222 ][ 25 ],
   alphaCSR[ 222 ][ 26 ],
   alphaCSR[ 222 ][ 27 ],
   alphaCSR[ 222 ][ 28 ],
   alphaCSR[ 222 ][ 29 ],
   alphaCSR[ 222 ][ 30 ],
   alphaCSR[ 222 ][ 31 ],
   alphaCSR[ 222 ][ 32 ],
   alphaCSR[ 222 ][ 33 ],
   alphaCSR[ 222 ][ 34 ],
   alphaCSR[ 222 ][ 35 ],
   alphaCSR[ 222 ][ 36 ],
   alphaCSR[ 222 ][ 37 ],
   alphaCSR[ 222 ][ 38 ],
   alphaCSR[ 222 ][ 39 ],
   alphaCSR[ 222 ][ 40 ],
   alphaCSR[ 222 ][ 41 ],
   alphaCSR[ 222 ][ 42 ],
   alphaCSR[ 222 ][ 43 ],
   alphaCSR[ 222 ][ 44 ],
   alphaCSR[ 222 ][ 45 ],
   alphaCSR[ 222 ][ 46 ],
   alphaCSR[ 222 ][ 47 ],
   alphaCSR[ 222 ][ 48 ],
   alphaCSR[ 222 ][ 49 ],
   alphaCSR[ 222 ][ 50 ],
   alphaCSR[ 222 ][ 51 ],
   alphaCSR[ 222 ][ 52 ],
   alphaCSR[ 222 ][ 53 ],
   alphaCSR[ 222 ][ 54 ],
   alphaCSR[ 222 ][ 55 ],
   alphaCSR[ 222 ][ 56 ],
   alphaCSR[ 222 ][ 57 ],
   alphaCSR[ 222 ][ 58 ],
   alphaCSR[ 222 ][ 59 ],
   alphaCSR[ 222 ][ 60 ],
   alphaCSR[ 222 ][ 61 ],
   alphaCSR[ 222 ][ 62 ],
   alphaCSR[ 222 ][ 63 ],
   alphaCSR[ 222 ][ 64 ],
   alphaCSR[ 222 ][ 65 ],
   alphaCSR[ 222 ][ 66 ],
   alphaCSR[ 222 ][ 67 ],
   alphaCSR[ 222 ][ 68 ],
   alphaCSR[ 222 ][ 69 ],
   alphaCSR[ 222 ][ 70 ],
   alphaCSR[ 222 ][ 71 ],
   alphaCSR[ 222 ][ 72 ],
   alphaCSR[ 222 ][ 73 ],
   alphaCSR[ 222 ][ 74 ],
   alphaCSR[ 222 ][ 75 ],
   alphaCSR[ 222 ][ 76 ],
   alphaCSR[ 222 ][ 77 ],
   alphaCSR[ 222 ][ 78 ],
   alphaCSR[ 222 ][ 79 ],
   alphaCSR[ 222 ][ 80 ],
   alphaCSR[ 222 ][ 81 ],
   alphaCSR[ 222 ][ 82 ],
   alphaCSR[ 222 ][ 83 ],
   alphaCSR[ 222 ][ 84 ],
   alphaCSR[ 222 ][ 85 ],
   alphaCSR[ 222 ][ 86 ],
   alphaCSR[ 222 ][ 87 ],
   alphaCSR[ 222 ][ 88 ],
   alphaCSR[ 222 ][ 89 ],
   alphaCSR[ 222 ][ 90 ],
   alphaCSR[ 222 ][ 91 ],
   alphaCSR[ 222 ][ 92 ],
   alphaCSR[ 222 ][ 93 ],
   alphaCSR[ 222 ][ 94 ],
   alphaCSR[ 222 ][ 95 ],
   alphaCSR[ 222 ][ 96 ],
   alphaCSR[ 222 ][ 97 ],
   alphaCSR[ 222 ][ 98 ],
   alphaCSR[ 222 ][ 99 ],
   alphaCSR[ 222 ][ 100 ],
   alphaCSR[ 222 ][ 101 ],
   alphaCSR[ 222 ][ 102 ],
   alphaCSR[ 222 ][ 103 ],
   alphaCSR[ 222 ][ 104 ],
   alphaCSR[ 222 ][ 105 ],
   alphaCSR[ 222 ][ 106 ],
   alphaCSR[ 222 ][ 107 ],
   alphaCSR[ 222 ][ 108 ],
   alphaCSR[ 222 ][ 109 ],
   alphaCSR[ 222 ][ 110 ],
   alphaCSR[ 222 ][ 111 ],
   alphaCSR[ 222 ][ 112 ],
   alphaCSR[ 222 ][ 113 ],
   alphaCSR[ 222 ][ 114 ],
   alphaCSR[ 222 ][ 115 ],
   alphaCSR[ 222 ][ 116 ],
   alphaCSR[ 222 ][ 117 ],
   alphaCSR[ 222 ][ 118 ],
   alphaCSR[ 222 ][ 119 ],
   alphaCSR[ 222 ][ 120 ],
   alphaCSR[ 222 ][ 121 ],
   alphaCSR[ 222 ][ 122 ],
   alphaCSR[ 222 ][ 123 ],
   alphaCSR[ 222 ][ 124 ],
   alphaCSR[ 222 ][ 125 ],
   alphaCSR[ 222 ][ 126 ],
   alphaCSR[ 222 ][ 127 ],
   alphaCSR[ 222 ][ 128 ],
   alphaCSR[ 222 ][ 129 ],
   alphaCSR[ 222 ][ 130 ],
   alphaCSR[ 222 ][ 131 ],
   alphaCSR[ 222 ][ 132 ],
   alphaCSR[ 222 ][ 133 ],
   alphaCSR[ 222 ][ 134 ],
   alphaCSR[ 222 ][ 135 ],
   alphaCSR[ 222 ][ 136 ],
   alphaCSR[ 222 ][ 137 ],
   alphaCSR[ 222 ][ 138 ],
   alphaCSR[ 222 ][ 139 ],
   alphaCSR[ 222 ][ 140 ],
   alphaCSR[ 222 ][ 141 ],
   alphaCSR[ 222 ][ 142 ],
   alphaCSR[ 222 ][ 143 ],
   alphaCSR[ 222 ][ 144 ],
   alphaCSR[ 222 ][ 145 ],
   alphaCSR[ 222 ][ 146 ],
   alphaCSR[ 222 ][ 147 ],
   alphaCSR[ 222 ][ 148 ],
   alphaCSR[ 222 ][ 149 ],
   alphaCSR[ 222 ][ 150 ],
   alphaCSR[ 222 ][ 151 ],
   alphaCSR[ 222 ][ 152 ],
   alphaCSR[ 222 ][ 153 ],
   alphaCSR[ 222 ][ 154 ],
   alphaCSR[ 222 ][ 155 ],
   alphaCSR[ 222 ][ 156 ],
   alphaCSR[ 222 ][ 157 ],
   alphaCSR[ 222 ][ 158 ],
   alphaCSR[ 222 ][ 159 ],
   alphaCSR[ 222 ][ 160 ],
   alphaCSR[ 222 ][ 161 ],
   alphaCSR[ 222 ][ 162 ],
   alphaCSR[ 222 ][ 163 ],
   alphaCSR[ 222 ][ 164 ],
   alphaCSR[ 222 ][ 165 ],
   alphaCSR[ 222 ][ 166 ],
   alphaCSR[ 222 ][ 167 ],
   alphaCSR[ 222 ][ 168 ],
   alphaCSR[ 222 ][ 169 ],
   alphaCSR[ 222 ][ 170 ],
   alphaCSR[ 222 ][ 171 ],
   alphaCSR[ 222 ][ 172 ],
   alphaCSR[ 222 ][ 173 ],
   alphaCSR[ 222 ][ 174 ],
   alphaCSR[ 222 ][ 175 ],
   alphaCSR[ 222 ][ 176 ],
   alphaCSR[ 222 ][ 177 ],
   alphaCSR[ 222 ][ 178 ],
   alphaCSR[ 222 ][ 179 ],
   alphaCSR[ 222 ][ 180 ],
   alphaCSR[ 222 ][ 181 ],
   alphaCSR[ 222 ][ 182 ],
   alphaCSR[ 222 ][ 183 ],
   alphaCSR[ 222 ][ 184 ],
   alphaCSR[ 222 ][ 185 ],
   alphaCSR[ 222 ][ 186 ],
   alphaCSR[ 222 ][ 187 ],
   alphaCSR[ 222 ][ 188 ],
   alphaCSR[ 222 ][ 189 ],
   alphaCSR[ 222 ][ 190 ],
   alphaCSR[ 222 ][ 191 ],
   alphaCSR[ 222 ][ 192 ],
   alphaCSR[ 222 ][ 193 ],
   alphaCSR[ 222 ][ 194 ],
   alphaCSR[ 222 ][ 195 ],
   alphaCSR[ 222 ][ 196 ],
   alphaCSR[ 222 ][ 197 ],
   alphaCSR[ 222 ][ 198 ],
   alphaCSR[ 222 ][ 199 ],
   alphaCSR[ 222 ][ 200 ],
   alphaCSR[ 222 ][ 201 ],
   alphaCSR[ 222 ][ 202 ],
   alphaCSR[ 222 ][ 203 ],
   alphaCSR[ 222 ][ 204 ],
   alphaCSR[ 222 ][ 205 ],
   alphaCSR[ 222 ][ 206 ],
   alphaCSR[ 222 ][ 207 ],
   alphaCSR[ 222 ][ 208 ],
   alphaCSR[ 222 ][ 209 ],
   alphaCSR[ 222 ][ 210 ],
   alphaCSR[ 222 ][ 211 ],
   alphaCSR[ 222 ][ 212 ],
   alphaCSR[ 222 ][ 213 ],
   alphaCSR[ 222 ][ 214 ],
   alphaCSR[ 222 ][ 215 ],
   alphaCSR[ 222 ][ 216 ],
   alphaCSR[ 222 ][ 217 ],
   alphaCSR[ 222 ][ 218 ],
   alphaCSR[ 222 ][ 219 ],
   alphaCSR[ 222 ][ 220 ],
   alphaCSR[ 222 ][ 221 ],
   alphaCSR[ 222 ][ 222 ],
   alphaCSR[ 222 ][ 223 ],
   alphaCSR[ 222 ][ 224 ],
   alphaCSR[ 222 ][ 225 ],
   alphaCSR[ 222 ][ 226 ],
   alphaCSR[ 222 ][ 227 ],
   alphaCSR[ 222 ][ 228 ],
   alphaCSR[ 222 ][ 229 ],
   alphaCSR[ 222 ][ 230 ],
   alphaCSR[ 222 ][ 231 ],
   alphaCSR[ 222 ][ 232 ],
   alphaCSR[ 222 ][ 233 ],
   alphaCSR[ 222 ][ 234 ],
   alphaCSR[ 222 ][ 235 ],
   alphaCSR[ 222 ][ 236 ],
   alphaCSR[ 222 ][ 237 ],
   alphaCSR[ 222 ][ 238 ],
   alphaCSR[ 222 ][ 239 ],
   alphaCSR[ 222 ][ 240 ],
   alphaCSR[ 222 ][ 241 ],
   alphaCSR[ 222 ][ 242 ],
   alphaCSR[ 222 ][ 243 ],
   alphaCSR[ 222 ][ 244 ],
   alphaCSR[ 222 ][ 245 ],
   alphaCSR[ 222 ][ 246 ],
   alphaCSR[ 222 ][ 247 ],
   alphaCSR[ 222 ][ 248 ],
   alphaCSR[ 222 ][ 249 ],
   alphaCSR[ 222 ][ 250 ],
   alphaCSR[ 222 ][ 251 ],
   alphaCSR[ 222 ][ 252 ],
   alphaCSR[ 222 ][ 253 ],
   alphaCSR[ 222 ][ 254 ],
   alphaCSR[ 222 ][ 255 ],
   alphaCSR[ 222 ][ 256 ],
   alphaCSR[ 222 ][ 257 ],
   alphaCSR[ 222 ][ 258 ],
   alphaCSR[ 222 ][ 259 ],
   alphaCSR[ 222 ][ 260 ],
   alphaCSR[ 222 ][ 261 ],
   alphaCSR[ 222 ][ 262 ],
   alphaCSR[ 222 ][ 263 ],
   alphaCSR[ 222 ][ 264 ],
   alphaCSR[ 222 ][ 265 ],
   alphaCSR[ 222 ][ 266 ],
   alphaCSR[ 222 ][ 267 ],
   alphaCSR[ 222 ][ 268 ],
   alphaCSR[ 222 ][ 269 ],
   alphaCSR[ 222 ][ 270 ],
   alphaCSR[ 222 ][ 271 ],
   alphaCSR[ 222 ][ 272 ],
   alphaCSR[ 222 ][ 273 ],
   alphaCSR[ 222 ][ 274 ],
   alphaCSR[ 222 ][ 275 ],
   alphaCSR[ 222 ][ 276 ],
   alphaCSR[ 222 ][ 277 ],
   alphaCSR[ 222 ][ 278 ],
   alphaCSR[ 222 ][ 279 ],
   alphaCSR[ 222 ][ 280 ],
   alphaCSR[ 222 ][ 281 ],
   alphaCSR[ 222 ][ 282 ],
   alphaCSR[ 222 ][ 283 ],
   alphaCSR[ 222 ][ 284 ],
   alphaCSR[ 222 ][ 285 ],
   alphaCSR[ 222 ][ 286 ],
   alphaCSR[ 222 ][ 287 ],
   alphaCSR[ 222 ][ 288 ],
   alphaCSR[ 222 ][ 289 ],
   alphaCSR[ 222 ][ 290 ],
   alphaCSR[ 222 ][ 291 ],
   alphaCSR[ 222 ][ 292 ],
   alphaCSR[ 222 ][ 293 ],
   alphaCSR[ 222 ][ 294 ],
   alphaCSR[ 222 ][ 295 ],
   alphaCSR[ 222 ][ 296 ],
   alphaCSR[ 222 ][ 297 ],
   alphaCSR[ 222 ][ 298 ],
   alphaCSR[ 222 ][ 299 ],
   alphaCSR[ 222 ][ 300 ],
   alphaCSR[ 222 ][ 301 ],
   alphaCSR[ 222 ][ 302 ],
   alphaCSR[ 222 ][ 303 ],
   alphaCSR[ 222 ][ 304 ],
   alphaCSR[ 222 ][ 305 ],
   alphaCSR[ 222 ][ 306 ],
   alphaCSR[ 222 ][ 307 ],
   alphaCSR[ 222 ][ 308 ],
   alphaCSR[ 222 ][ 309 ],
   alphaCSR[ 222 ][ 310 ],
   alphaCSR[ 222 ][ 311 ],
   alphaCSR[ 222 ][ 312 ],
   alphaCSR[ 222 ][ 313 ],
   alphaCSR[ 222 ][ 314 ],
   alphaCSR[ 222 ][ 315 ],
   alphaCSR[ 222 ][ 316 ],
   alphaCSR[ 222 ][ 317 ],
   alphaCSR[ 222 ][ 318 ],
   alphaCSR[ 222 ][ 319 ],
   alphaCSR[ 222 ][ 320 ],
   alphaCSR[ 222 ][ 321 ],
   alphaCSR[ 222 ][ 322 ],
   alphaCSR[ 222 ][ 323 ],
   alphaCSR[ 222 ][ 324 ],
   alphaCSR[ 222 ][ 325 ],
   alphaCSR[ 222 ][ 326 ],
   alphaCSR[ 222 ][ 327 ],
   alphaCSR[ 222 ][ 328 ],
   alphaCSR[ 222 ][ 329 ],
   alphaCSR[ 222 ][ 330 ],
   alphaCSR[ 222 ][ 331 ],
   alphaCSR[ 222 ][ 332 ],
   alphaCSR[ 222 ][ 333 ],
   alphaCSR[ 222 ][ 334 ],
   alphaCSR[ 222 ][ 335 ],
   alphaCSR[ 222 ][ 336 ],
   alphaCSR[ 222 ][ 337 ],
   alphaCSR[ 222 ][ 338 ],
   alphaCSR[ 222 ][ 339 ],
   alphaCSR[ 222 ][ 340 ],
   alphaCSR[ 222 ][ 341 ],
   alphaCSR[ 222 ][ 342 ],
   alphaCSR[ 222 ][ 343 ],
   alphaCSR[ 222 ][ 344 ],
   alphaCSR[ 222 ][ 345 ],
   alphaCSR[ 222 ][ 346 ],
   alphaCSR[ 222 ][ 347 ],
   alphaCSR[ 222 ][ 348 ],
   alphaCSR[ 222 ][ 349 ],
   alphaCSR[ 222 ][ 350 ],
   alphaCSR[ 222 ][ 351 ],
   alphaCSR[ 222 ][ 352 ],
   alphaCSR[ 222 ][ 353 ],
   alphaCSR[ 222 ][ 354 ],
   alphaCSR[ 222 ][ 355 ],
   alphaCSR[ 222 ][ 356 ],
   alphaCSR[ 222 ][ 357 ],
   alphaCSR[ 222 ][ 358 ],
   alphaCSR[ 222 ][ 359 ],
   alphaCSR[ 222 ][ 360 ],
   alphaCSR[ 222 ][ 361 ],
   alphaCSR[ 222 ][ 362 ],
   alphaCSR[ 222 ][ 363 ],
   alphaCSR[ 222 ][ 364 ],
   alphaCSR[ 222 ][ 365 ],
   alphaCSR[ 222 ][ 366 ],
   alphaCSR[ 222 ][ 367 ],
   alphaCSR[ 222 ][ 368 ],
   alphaCSR[ 222 ][ 369 ],
   alphaCSR[ 222 ][ 370 ],
   alphaCSR[ 222 ][ 371 ],
   alphaCSR[ 222 ][ 372 ],
   alphaCSR[ 222 ][ 373 ],
   alphaCSR[ 222 ][ 374 ],
   alphaCSR[ 222 ][ 375 ],
   alphaCSR[ 222 ][ 376 ],
   alphaCSR[ 222 ][ 377 ],
   alphaCSR[ 222 ][ 378 ],
   alphaCSR[ 222 ][ 379 ],
   alphaCSR[ 222 ][ 380 ],
   alphaCSR[ 222 ][ 381 ],
   alphaCSR[ 222 ][ 382 ],
   alphaCSR[ 222 ][ 383 ],
   alphaCSR[ 223 ][ 0 ],
   alphaCSR[ 223 ][ 1 ],
   alphaCSR[ 223 ][ 2 ],
   alphaCSR[ 223 ][ 3 ],
   alphaCSR[ 223 ][ 4 ],
   alphaCSR[ 223 ][ 5 ],
   alphaCSR[ 223 ][ 6 ],
   alphaCSR[ 223 ][ 7 ],
   alphaCSR[ 223 ][ 8 ],
   alphaCSR[ 223 ][ 9 ],
   alphaCSR[ 223 ][ 10 ],
   alphaCSR[ 223 ][ 11 ],
   alphaCSR[ 223 ][ 12 ],
   alphaCSR[ 223 ][ 13 ],
   alphaCSR[ 223 ][ 14 ],
   alphaCSR[ 223 ][ 15 ],
   alphaCSR[ 223 ][ 16 ],
   alphaCSR[ 223 ][ 17 ],
   alphaCSR[ 223 ][ 18 ],
   alphaCSR[ 223 ][ 19 ],
   alphaCSR[ 223 ][ 20 ],
   alphaCSR[ 223 ][ 21 ],
   alphaCSR[ 223 ][ 22 ],
   alphaCSR[ 223 ][ 23 ],
   alphaCSR[ 223 ][ 24 ],
   alphaCSR[ 223 ][ 25 ],
   alphaCSR[ 223 ][ 26 ],
   alphaCSR[ 223 ][ 27 ],
   alphaCSR[ 223 ][ 28 ],
   alphaCSR[ 223 ][ 29 ],
   alphaCSR[ 223 ][ 30 ],
   alphaCSR[ 223 ][ 31 ],
   alphaCSR[ 223 ][ 32 ],
   alphaCSR[ 223 ][ 33 ],
   alphaCSR[ 223 ][ 34 ],
   alphaCSR[ 223 ][ 35 ],
   alphaCSR[ 223 ][ 36 ],
   alphaCSR[ 223 ][ 37 ],
   alphaCSR[ 223 ][ 38 ],
   alphaCSR[ 223 ][ 39 ],
   alphaCSR[ 223 ][ 40 ],
   alphaCSR[ 223 ][ 41 ],
   alphaCSR[ 223 ][ 42 ],
   alphaCSR[ 223 ][ 43 ],
   alphaCSR[ 223 ][ 44 ],
   alphaCSR[ 223 ][ 45 ],
   alphaCSR[ 223 ][ 46 ],
   alphaCSR[ 223 ][ 47 ],
   alphaCSR[ 223 ][ 48 ],
   alphaCSR[ 223 ][ 49 ],
   alphaCSR[ 223 ][ 50 ],
   alphaCSR[ 223 ][ 51 ],
   alphaCSR[ 223 ][ 52 ],
   alphaCSR[ 223 ][ 53 ],
   alphaCSR[ 223 ][ 54 ],
   alphaCSR[ 223 ][ 55 ],
   alphaCSR[ 223 ][ 56 ],
   alphaCSR[ 223 ][ 57 ],
   alphaCSR[ 223 ][ 58 ],
   alphaCSR[ 223 ][ 59 ],
   alphaCSR[ 223 ][ 60 ],
   alphaCSR[ 223 ][ 61 ],
   alphaCSR[ 223 ][ 62 ],
   alphaCSR[ 223 ][ 63 ],
   alphaCSR[ 223 ][ 64 ],
   alphaCSR[ 223 ][ 65 ],
   alphaCSR[ 223 ][ 66 ],
   alphaCSR[ 223 ][ 67 ],
   alphaCSR[ 223 ][ 68 ],
   alphaCSR[ 223 ][ 69 ],
   alphaCSR[ 223 ][ 70 ],
   alphaCSR[ 223 ][ 71 ],
   alphaCSR[ 223 ][ 72 ],
   alphaCSR[ 223 ][ 73 ],
   alphaCSR[ 223 ][ 74 ],
   alphaCSR[ 223 ][ 75 ],
   alphaCSR[ 223 ][ 76 ],
   alphaCSR[ 223 ][ 77 ],
   alphaCSR[ 223 ][ 78 ],
   alphaCSR[ 223 ][ 79 ],
   alphaCSR[ 223 ][ 80 ],
   alphaCSR[ 223 ][ 81 ],
   alphaCSR[ 223 ][ 82 ],
   alphaCSR[ 223 ][ 83 ],
   alphaCSR[ 223 ][ 84 ],
   alphaCSR[ 223 ][ 85 ],
   alphaCSR[ 223 ][ 86 ],
   alphaCSR[ 223 ][ 87 ],
   alphaCSR[ 223 ][ 88 ],
   alphaCSR[ 223 ][ 89 ],
   alphaCSR[ 223 ][ 90 ],
   alphaCSR[ 223 ][ 91 ],
   alphaCSR[ 223 ][ 92 ],
   alphaCSR[ 223 ][ 93 ],
   alphaCSR[ 223 ][ 94 ],
   alphaCSR[ 223 ][ 95 ],
   alphaCSR[ 223 ][ 96 ],
   alphaCSR[ 223 ][ 97 ],
   alphaCSR[ 223 ][ 98 ],
   alphaCSR[ 223 ][ 99 ],
   alphaCSR[ 223 ][ 100 ],
   alphaCSR[ 223 ][ 101 ],
   alphaCSR[ 223 ][ 102 ],
   alphaCSR[ 223 ][ 103 ],
   alphaCSR[ 223 ][ 104 ],
   alphaCSR[ 223 ][ 105 ],
   alphaCSR[ 223 ][ 106 ],
   alphaCSR[ 223 ][ 107 ],
   alphaCSR[ 223 ][ 108 ],
   alphaCSR[ 223 ][ 109 ],
   alphaCSR[ 223 ][ 110 ],
   alphaCSR[ 223 ][ 111 ],
   alphaCSR[ 223 ][ 112 ],
   alphaCSR[ 223 ][ 113 ],
   alphaCSR[ 223 ][ 114 ],
   alphaCSR[ 223 ][ 115 ],
   alphaCSR[ 223 ][ 116 ],
   alphaCSR[ 223 ][ 117 ],
   alphaCSR[ 223 ][ 118 ],
   alphaCSR[ 223 ][ 119 ],
   alphaCSR[ 223 ][ 120 ],
   alphaCSR[ 223 ][ 121 ],
   alphaCSR[ 223 ][ 122 ],
   alphaCSR[ 223 ][ 123 ],
   alphaCSR[ 223 ][ 124 ],
   alphaCSR[ 223 ][ 125 ],
   alphaCSR[ 223 ][ 126 ],
   alphaCSR[ 223 ][ 127 ],
   alphaCSR[ 223 ][ 128 ],
   alphaCSR[ 223 ][ 129 ],
   alphaCSR[ 223 ][ 130 ],
   alphaCSR[ 223 ][ 131 ],
   alphaCSR[ 223 ][ 132 ],
   alphaCSR[ 223 ][ 133 ],
   alphaCSR[ 223 ][ 134 ],
   alphaCSR[ 223 ][ 135 ],
   alphaCSR[ 223 ][ 136 ],
   alphaCSR[ 223 ][ 137 ],
   alphaCSR[ 223 ][ 138 ],
   alphaCSR[ 223 ][ 139 ],
   alphaCSR[ 223 ][ 140 ],
   alphaCSR[ 223 ][ 141 ],
   alphaCSR[ 223 ][ 142 ],
   alphaCSR[ 223 ][ 143 ],
   alphaCSR[ 223 ][ 144 ],
   alphaCSR[ 223 ][ 145 ],
   alphaCSR[ 223 ][ 146 ],
   alphaCSR[ 223 ][ 147 ],
   alphaCSR[ 223 ][ 148 ],
   alphaCSR[ 223 ][ 149 ],
   alphaCSR[ 223 ][ 150 ],
   alphaCSR[ 223 ][ 151 ],
   alphaCSR[ 223 ][ 152 ],
   alphaCSR[ 223 ][ 153 ],
   alphaCSR[ 223 ][ 154 ],
   alphaCSR[ 223 ][ 155 ],
   alphaCSR[ 223 ][ 156 ],
   alphaCSR[ 223 ][ 157 ],
   alphaCSR[ 223 ][ 158 ],
   alphaCSR[ 223 ][ 159 ],
   alphaCSR[ 223 ][ 160 ],
   alphaCSR[ 223 ][ 161 ],
   alphaCSR[ 223 ][ 162 ],
   alphaCSR[ 223 ][ 163 ],
   alphaCSR[ 223 ][ 164 ],
   alphaCSR[ 223 ][ 165 ],
   alphaCSR[ 223 ][ 166 ],
   alphaCSR[ 223 ][ 167 ],
   alphaCSR[ 223 ][ 168 ],
   alphaCSR[ 223 ][ 169 ],
   alphaCSR[ 223 ][ 170 ],
   alphaCSR[ 223 ][ 171 ],
   alphaCSR[ 223 ][ 172 ],
   alphaCSR[ 223 ][ 173 ],
   alphaCSR[ 223 ][ 174 ],
   alphaCSR[ 223 ][ 175 ],
   alphaCSR[ 223 ][ 176 ],
   alphaCSR[ 223 ][ 177 ],
   alphaCSR[ 223 ][ 178 ],
   alphaCSR[ 223 ][ 179 ],
   alphaCSR[ 223 ][ 180 ],
   alphaCSR[ 223 ][ 181 ],
   alphaCSR[ 223 ][ 182 ],
   alphaCSR[ 223 ][ 183 ],
   alphaCSR[ 223 ][ 184 ],
   alphaCSR[ 223 ][ 185 ],
   alphaCSR[ 223 ][ 186 ],
   alphaCSR[ 223 ][ 187 ],
   alphaCSR[ 223 ][ 188 ],
   alphaCSR[ 223 ][ 189 ],
   alphaCSR[ 223 ][ 190 ],
   alphaCSR[ 223 ][ 191 ],
   alphaCSR[ 223 ][ 192 ],
   alphaCSR[ 223 ][ 193 ],
   alphaCSR[ 223 ][ 194 ],
   alphaCSR[ 223 ][ 195 ],
   alphaCSR[ 223 ][ 196 ],
   alphaCSR[ 223 ][ 197 ],
   alphaCSR[ 223 ][ 198 ],
   alphaCSR[ 223 ][ 199 ],
   alphaCSR[ 223 ][ 200 ],
   alphaCSR[ 223 ][ 201 ],
   alphaCSR[ 223 ][ 202 ],
   alphaCSR[ 223 ][ 203 ],
   alphaCSR[ 223 ][ 204 ],
   alphaCSR[ 223 ][ 205 ],
   alphaCSR[ 223 ][ 206 ],
   alphaCSR[ 223 ][ 207 ],
   alphaCSR[ 223 ][ 208 ],
   alphaCSR[ 223 ][ 209 ],
   alphaCSR[ 223 ][ 210 ],
   alphaCSR[ 223 ][ 211 ],
   alphaCSR[ 223 ][ 212 ],
   alphaCSR[ 223 ][ 213 ],
   alphaCSR[ 223 ][ 214 ],
   alphaCSR[ 223 ][ 215 ],
   alphaCSR[ 223 ][ 216 ],
   alphaCSR[ 223 ][ 217 ],
   alphaCSR[ 223 ][ 218 ],
   alphaCSR[ 223 ][ 219 ],
   alphaCSR[ 223 ][ 220 ],
   alphaCSR[ 223 ][ 221 ],
   alphaCSR[ 223 ][ 222 ],
   alphaCSR[ 223 ][ 223 ],
   alphaCSR[ 223 ][ 224 ],
   alphaCSR[ 223 ][ 225 ],
   alphaCSR[ 223 ][ 226 ],
   alphaCSR[ 223 ][ 227 ],
   alphaCSR[ 223 ][ 228 ],
   alphaCSR[ 223 ][ 229 ],
   alphaCSR[ 223 ][ 230 ],
   alphaCSR[ 223 ][ 231 ],
   alphaCSR[ 223 ][ 232 ],
   alphaCSR[ 223 ][ 233 ],
   alphaCSR[ 223 ][ 234 ],
   alphaCSR[ 223 ][ 235 ],
   alphaCSR[ 223 ][ 236 ],
   alphaCSR[ 223 ][ 237 ],
   alphaCSR[ 223 ][ 238 ],
   alphaCSR[ 223 ][ 239 ],
   alphaCSR[ 223 ][ 240 ],
   alphaCSR[ 223 ][ 241 ],
   alphaCSR[ 223 ][ 242 ],
   alphaCSR[ 223 ][ 243 ],
   alphaCSR[ 223 ][ 244 ],
   alphaCSR[ 223 ][ 245 ],
   alphaCSR[ 223 ][ 246 ],
   alphaCSR[ 223 ][ 247 ],
   alphaCSR[ 223 ][ 248 ],
   alphaCSR[ 223 ][ 249 ],
   alphaCSR[ 223 ][ 250 ],
   alphaCSR[ 223 ][ 251 ],
   alphaCSR[ 223 ][ 252 ],
   alphaCSR[ 223 ][ 253 ],
   alphaCSR[ 223 ][ 254 ],
   alphaCSR[ 223 ][ 255 ],
   alphaCSR[ 223 ][ 256 ],
   alphaCSR[ 223 ][ 257 ],
   alphaCSR[ 223 ][ 258 ],
   alphaCSR[ 223 ][ 259 ],
   alphaCSR[ 223 ][ 260 ],
   alphaCSR[ 223 ][ 261 ],
   alphaCSR[ 223 ][ 262 ],
   alphaCSR[ 223 ][ 263 ],
   alphaCSR[ 223 ][ 264 ],
   alphaCSR[ 223 ][ 265 ],
   alphaCSR[ 223 ][ 266 ],
   alphaCSR[ 223 ][ 267 ],
   alphaCSR[ 223 ][ 268 ],
   alphaCSR[ 223 ][ 269 ],
   alphaCSR[ 223 ][ 270 ],
   alphaCSR[ 223 ][ 271 ],
   alphaCSR[ 223 ][ 272 ],
   alphaCSR[ 223 ][ 273 ],
   alphaCSR[ 223 ][ 274 ],
   alphaCSR[ 223 ][ 275 ],
   alphaCSR[ 223 ][ 276 ],
   alphaCSR[ 223 ][ 277 ],
   alphaCSR[ 223 ][ 278 ],
   alphaCSR[ 223 ][ 279 ],
   alphaCSR[ 223 ][ 280 ],
   alphaCSR[ 223 ][ 281 ],
   alphaCSR[ 223 ][ 282 ],
   alphaCSR[ 223 ][ 283 ],
   alphaCSR[ 223 ][ 284 ],
   alphaCSR[ 223 ][ 285 ],
   alphaCSR[ 223 ][ 286 ],
   alphaCSR[ 223 ][ 287 ],
   alphaCSR[ 223 ][ 288 ],
   alphaCSR[ 223 ][ 289 ],
   alphaCSR[ 223 ][ 290 ],
   alphaCSR[ 223 ][ 291 ],
   alphaCSR[ 223 ][ 292 ],
   alphaCSR[ 223 ][ 293 ],
   alphaCSR[ 223 ][ 294 ],
   alphaCSR[ 223 ][ 295 ],
   alphaCSR[ 223 ][ 296 ],
   alphaCSR[ 223 ][ 297 ],
   alphaCSR[ 223 ][ 298 ],
   alphaCSR[ 223 ][ 299 ],
   alphaCSR[ 223 ][ 300 ],
   alphaCSR[ 223 ][ 301 ],
   alphaCSR[ 223 ][ 302 ],
   alphaCSR[ 223 ][ 303 ],
   alphaCSR[ 223 ][ 304 ],
   alphaCSR[ 223 ][ 305 ],
   alphaCSR[ 223 ][ 306 ],
   alphaCSR[ 223 ][ 307 ],
   alphaCSR[ 223 ][ 308 ],
   alphaCSR[ 223 ][ 309 ],
   alphaCSR[ 223 ][ 310 ],
   alphaCSR[ 223 ][ 311 ],
   alphaCSR[ 223 ][ 312 ],
   alphaCSR[ 223 ][ 313 ],
   alphaCSR[ 223 ][ 314 ],
   alphaCSR[ 223 ][ 315 ],
   alphaCSR[ 223 ][ 316 ],
   alphaCSR[ 223 ][ 317 ],
   alphaCSR[ 223 ][ 318 ],
   alphaCSR[ 223 ][ 319 ],
   alphaCSR[ 223 ][ 320 ],
   alphaCSR[ 223 ][ 321 ],
   alphaCSR[ 223 ][ 322 ],
   alphaCSR[ 223 ][ 323 ],
   alphaCSR[ 223 ][ 324 ],
   alphaCSR[ 223 ][ 325 ],
   alphaCSR[ 223 ][ 326 ],
   alphaCSR[ 223 ][ 327 ],
   alphaCSR[ 223 ][ 328 ],
   alphaCSR[ 223 ][ 329 ],
   alphaCSR[ 223 ][ 330 ],
   alphaCSR[ 223 ][ 331 ],
   alphaCSR[ 223 ][ 332 ],
   alphaCSR[ 223 ][ 333 ],
   alphaCSR[ 223 ][ 334 ],
   alphaCSR[ 223 ][ 335 ],
   alphaCSR[ 223 ][ 336 ],
   alphaCSR[ 223 ][ 337 ],
   alphaCSR[ 223 ][ 338 ],
   alphaCSR[ 223 ][ 339 ],
   alphaCSR[ 223 ][ 340 ],
   alphaCSR[ 223 ][ 341 ],
   alphaCSR[ 223 ][ 342 ],
   alphaCSR[ 223 ][ 343 ],
   alphaCSR[ 223 ][ 344 ],
   alphaCSR[ 223 ][ 345 ],
   alphaCSR[ 223 ][ 346 ],
   alphaCSR[ 223 ][ 347 ],
   alphaCSR[ 223 ][ 348 ],
   alphaCSR[ 223 ][ 349 ],
   alphaCSR[ 223 ][ 350 ],
   alphaCSR[ 223 ][ 351 ],
   alphaCSR[ 223 ][ 352 ],
   alphaCSR[ 223 ][ 353 ],
   alphaCSR[ 223 ][ 354 ],
   alphaCSR[ 223 ][ 355 ],
   alphaCSR[ 223 ][ 356 ],
   alphaCSR[ 223 ][ 357 ],
   alphaCSR[ 223 ][ 358 ],
   alphaCSR[ 223 ][ 359 ],
   alphaCSR[ 223 ][ 360 ],
   alphaCSR[ 223 ][ 361 ],
   alphaCSR[ 223 ][ 362 ],
   alphaCSR[ 223 ][ 363 ],
   alphaCSR[ 223 ][ 364 ],
   alphaCSR[ 223 ][ 365 ],
   alphaCSR[ 223 ][ 366 ],
   alphaCSR[ 223 ][ 367 ],
   alphaCSR[ 223 ][ 368 ],
   alphaCSR[ 223 ][ 369 ],
   alphaCSR[ 223 ][ 370 ],
   alphaCSR[ 223 ][ 371 ],
   alphaCSR[ 223 ][ 372 ],
   alphaCSR[ 223 ][ 373 ],
   alphaCSR[ 223 ][ 374 ],
   alphaCSR[ 223 ][ 375 ],
   alphaCSR[ 223 ][ 376 ],
   alphaCSR[ 223 ][ 377 ],
   alphaCSR[ 223 ][ 378 ],
   alphaCSR[ 223 ][ 379 ],
   alphaCSR[ 223 ][ 380 ],
   alphaCSR[ 223 ][ 381 ],
   alphaCSR[ 223 ][ 382 ],
   alphaCSR[ 223 ][ 383 ],
   alphaCSR[ 224 ][ 0 ],
   alphaCSR[ 224 ][ 1 ],
   alphaCSR[ 224 ][ 2 ],
   alphaCSR[ 224 ][ 3 ],
   alphaCSR[ 224 ][ 4 ],
   alphaCSR[ 224 ][ 5 ],
   alphaCSR[ 224 ][ 6 ],
   alphaCSR[ 224 ][ 7 ],
   alphaCSR[ 224 ][ 8 ],
   alphaCSR[ 224 ][ 9 ],
   alphaCSR[ 224 ][ 10 ],
   alphaCSR[ 224 ][ 11 ],
   alphaCSR[ 224 ][ 12 ],
   alphaCSR[ 224 ][ 13 ],
   alphaCSR[ 224 ][ 14 ],
   alphaCSR[ 224 ][ 15 ],
   alphaCSR[ 224 ][ 16 ],
   alphaCSR[ 224 ][ 17 ],
   alphaCSR[ 224 ][ 18 ],
   alphaCSR[ 224 ][ 19 ],
   alphaCSR[ 224 ][ 20 ],
   alphaCSR[ 224 ][ 21 ],
   alphaCSR[ 224 ][ 22 ],
   alphaCSR[ 224 ][ 23 ],
   alphaCSR[ 224 ][ 24 ],
   alphaCSR[ 224 ][ 25 ],
   alphaCSR[ 224 ][ 26 ],
   alphaCSR[ 224 ][ 27 ],
   alphaCSR[ 224 ][ 28 ],
   alphaCSR[ 224 ][ 29 ],
   alphaCSR[ 224 ][ 30 ],
   alphaCSR[ 224 ][ 31 ],
   alphaCSR[ 224 ][ 32 ],
   alphaCSR[ 224 ][ 33 ],
   alphaCSR[ 224 ][ 34 ],
   alphaCSR[ 224 ][ 35 ],
   alphaCSR[ 224 ][ 36 ],
   alphaCSR[ 224 ][ 37 ],
   alphaCSR[ 224 ][ 38 ],
   alphaCSR[ 224 ][ 39 ],
   alphaCSR[ 224 ][ 40 ],
   alphaCSR[ 224 ][ 41 ],
   alphaCSR[ 224 ][ 42 ],
   alphaCSR[ 224 ][ 43 ],
   alphaCSR[ 224 ][ 44 ],
   alphaCSR[ 224 ][ 45 ],
   alphaCSR[ 224 ][ 46 ],
   alphaCSR[ 224 ][ 47 ],
   alphaCSR[ 224 ][ 48 ],
   alphaCSR[ 224 ][ 49 ],
   alphaCSR[ 224 ][ 50 ],
   alphaCSR[ 224 ][ 51 ],
   alphaCSR[ 224 ][ 52 ],
   alphaCSR[ 224 ][ 53 ],
   alphaCSR[ 224 ][ 54 ],
   alphaCSR[ 224 ][ 55 ],
   alphaCSR[ 224 ][ 56 ],
   alphaCSR[ 224 ][ 57 ],
   alphaCSR[ 224 ][ 58 ],
   alphaCSR[ 224 ][ 59 ],
   alphaCSR[ 224 ][ 60 ],
   alphaCSR[ 224 ][ 61 ],
   alphaCSR[ 224 ][ 62 ],
   alphaCSR[ 224 ][ 63 ],
   alphaCSR[ 224 ][ 64 ],
   alphaCSR[ 224 ][ 65 ],
   alphaCSR[ 224 ][ 66 ],
   alphaCSR[ 224 ][ 67 ],
   alphaCSR[ 224 ][ 68 ],
   alphaCSR[ 224 ][ 69 ],
   alphaCSR[ 224 ][ 70 ],
   alphaCSR[ 224 ][ 71 ],
   alphaCSR[ 224 ][ 72 ],
   alphaCSR[ 224 ][ 73 ],
   alphaCSR[ 224 ][ 74 ],
   alphaCSR[ 224 ][ 75 ],
   alphaCSR[ 224 ][ 76 ],
   alphaCSR[ 224 ][ 77 ],
   alphaCSR[ 224 ][ 78 ],
   alphaCSR[ 224 ][ 79 ],
   alphaCSR[ 224 ][ 80 ],
   alphaCSR[ 224 ][ 81 ],
   alphaCSR[ 224 ][ 82 ],
   alphaCSR[ 224 ][ 83 ],
   alphaCSR[ 224 ][ 84 ],
   alphaCSR[ 224 ][ 85 ],
   alphaCSR[ 224 ][ 86 ],
   alphaCSR[ 224 ][ 87 ],
   alphaCSR[ 224 ][ 88 ],
   alphaCSR[ 224 ][ 89 ],
   alphaCSR[ 224 ][ 90 ],
   alphaCSR[ 224 ][ 91 ],
   alphaCSR[ 224 ][ 92 ],
   alphaCSR[ 224 ][ 93 ],
   alphaCSR[ 224 ][ 94 ],
   alphaCSR[ 224 ][ 95 ],
   alphaCSR[ 224 ][ 96 ],
   alphaCSR[ 224 ][ 97 ],
   alphaCSR[ 224 ][ 98 ],
   alphaCSR[ 224 ][ 99 ],
   alphaCSR[ 224 ][ 100 ],
   alphaCSR[ 224 ][ 101 ],
   alphaCSR[ 224 ][ 102 ],
   alphaCSR[ 224 ][ 103 ],
   alphaCSR[ 224 ][ 104 ],
   alphaCSR[ 224 ][ 105 ],
   alphaCSR[ 224 ][ 106 ],
   alphaCSR[ 224 ][ 107 ],
   alphaCSR[ 224 ][ 108 ],
   alphaCSR[ 224 ][ 109 ],
   alphaCSR[ 224 ][ 110 ],
   alphaCSR[ 224 ][ 111 ],
   alphaCSR[ 224 ][ 112 ],
   alphaCSR[ 224 ][ 113 ],
   alphaCSR[ 224 ][ 114 ],
   alphaCSR[ 224 ][ 115 ],
   alphaCSR[ 224 ][ 116 ],
   alphaCSR[ 224 ][ 117 ],
   alphaCSR[ 224 ][ 118 ],
   alphaCSR[ 224 ][ 119 ],
   alphaCSR[ 224 ][ 120 ],
   alphaCSR[ 224 ][ 121 ],
   alphaCSR[ 224 ][ 122 ],
   alphaCSR[ 224 ][ 123 ],
   alphaCSR[ 224 ][ 124 ],
   alphaCSR[ 224 ][ 125 ],
   alphaCSR[ 224 ][ 126 ],
   alphaCSR[ 224 ][ 127 ],
   alphaCSR[ 224 ][ 128 ],
   alphaCSR[ 224 ][ 129 ],
   alphaCSR[ 224 ][ 130 ],
   alphaCSR[ 224 ][ 131 ],
   alphaCSR[ 224 ][ 132 ],
   alphaCSR[ 224 ][ 133 ],
   alphaCSR[ 224 ][ 134 ],
   alphaCSR[ 224 ][ 135 ],
   alphaCSR[ 224 ][ 136 ],
   alphaCSR[ 224 ][ 137 ],
   alphaCSR[ 224 ][ 138 ],
   alphaCSR[ 224 ][ 139 ],
   alphaCSR[ 224 ][ 140 ],
   alphaCSR[ 224 ][ 141 ],
   alphaCSR[ 224 ][ 142 ],
   alphaCSR[ 224 ][ 143 ],
   alphaCSR[ 224 ][ 144 ],
   alphaCSR[ 224 ][ 145 ],
   alphaCSR[ 224 ][ 146 ],
   alphaCSR[ 224 ][ 147 ],
   alphaCSR[ 224 ][ 148 ],
   alphaCSR[ 224 ][ 149 ],
   alphaCSR[ 224 ][ 150 ],
   alphaCSR[ 224 ][ 151 ],
   alphaCSR[ 224 ][ 152 ],
   alphaCSR[ 224 ][ 153 ],
   alphaCSR[ 224 ][ 154 ],
   alphaCSR[ 224 ][ 155 ],
   alphaCSR[ 224 ][ 156 ],
   alphaCSR[ 224 ][ 157 ],
   alphaCSR[ 224 ][ 158 ],
   alphaCSR[ 224 ][ 159 ],
   alphaCSR[ 224 ][ 160 ],
   alphaCSR[ 224 ][ 161 ],
   alphaCSR[ 224 ][ 162 ],
   alphaCSR[ 224 ][ 163 ],
   alphaCSR[ 224 ][ 164 ],
   alphaCSR[ 224 ][ 165 ],
   alphaCSR[ 224 ][ 166 ],
   alphaCSR[ 224 ][ 167 ],
   alphaCSR[ 224 ][ 168 ],
   alphaCSR[ 224 ][ 169 ],
   alphaCSR[ 224 ][ 170 ],
   alphaCSR[ 224 ][ 171 ],
   alphaCSR[ 224 ][ 172 ],
   alphaCSR[ 224 ][ 173 ],
   alphaCSR[ 224 ][ 174 ],
   alphaCSR[ 224 ][ 175 ],
   alphaCSR[ 224 ][ 176 ],
   alphaCSR[ 224 ][ 177 ],
   alphaCSR[ 224 ][ 178 ],
   alphaCSR[ 224 ][ 179 ],
   alphaCSR[ 224 ][ 180 ],
   alphaCSR[ 224 ][ 181 ],
   alphaCSR[ 224 ][ 182 ],
   alphaCSR[ 224 ][ 183 ],
   alphaCSR[ 224 ][ 184 ],
   alphaCSR[ 224 ][ 185 ],
   alphaCSR[ 224 ][ 186 ],
   alphaCSR[ 224 ][ 187 ],
   alphaCSR[ 224 ][ 188 ],
   alphaCSR[ 224 ][ 189 ],
   alphaCSR[ 224 ][ 190 ],
   alphaCSR[ 224 ][ 191 ],
   alphaCSR[ 224 ][ 192 ],
   alphaCSR[ 224 ][ 193 ],
   alphaCSR[ 224 ][ 194 ],
   alphaCSR[ 224 ][ 195 ],
   alphaCSR[ 224 ][ 196 ],
   alphaCSR[ 224 ][ 197 ],
   alphaCSR[ 224 ][ 198 ],
   alphaCSR[ 224 ][ 199 ],
   alphaCSR[ 224 ][ 200 ],
   alphaCSR[ 224 ][ 201 ],
   alphaCSR[ 224 ][ 202 ],
   alphaCSR[ 224 ][ 203 ],
   alphaCSR[ 224 ][ 204 ],
   alphaCSR[ 224 ][ 205 ],
   alphaCSR[ 224 ][ 206 ],
   alphaCSR[ 224 ][ 207 ],
   alphaCSR[ 224 ][ 208 ],
   alphaCSR[ 224 ][ 209 ],
   alphaCSR[ 224 ][ 210 ],
   alphaCSR[ 224 ][ 211 ],
   alphaCSR[ 224 ][ 212 ],
   alphaCSR[ 224 ][ 213 ],
   alphaCSR[ 224 ][ 214 ],
   alphaCSR[ 224 ][ 215 ],
   alphaCSR[ 224 ][ 216 ],
   alphaCSR[ 224 ][ 217 ],
   alphaCSR[ 224 ][ 218 ],
   alphaCSR[ 224 ][ 219 ],
   alphaCSR[ 224 ][ 220 ],
   alphaCSR[ 224 ][ 221 ],
   alphaCSR[ 224 ][ 222 ],
   alphaCSR[ 224 ][ 223 ],
   alphaCSR[ 224 ][ 224 ],
   alphaCSR[ 224 ][ 225 ],
   alphaCSR[ 224 ][ 226 ],
   alphaCSR[ 224 ][ 227 ],
   alphaCSR[ 224 ][ 228 ],
   alphaCSR[ 224 ][ 229 ],
   alphaCSR[ 224 ][ 230 ],
   alphaCSR[ 224 ][ 231 ],
   alphaCSR[ 224 ][ 232 ],
   alphaCSR[ 224 ][ 233 ],
   alphaCSR[ 224 ][ 234 ],
   alphaCSR[ 224 ][ 235 ],
   alphaCSR[ 224 ][ 236 ],
   alphaCSR[ 224 ][ 237 ],
   alphaCSR[ 224 ][ 238 ],
   alphaCSR[ 224 ][ 239 ],
   alphaCSR[ 224 ][ 240 ],
   alphaCSR[ 224 ][ 241 ],
   alphaCSR[ 224 ][ 242 ],
   alphaCSR[ 224 ][ 243 ],
   alphaCSR[ 224 ][ 244 ],
   alphaCSR[ 224 ][ 245 ],
   alphaCSR[ 224 ][ 246 ],
   alphaCSR[ 224 ][ 247 ],
   alphaCSR[ 224 ][ 248 ],
   alphaCSR[ 224 ][ 249 ],
   alphaCSR[ 224 ][ 250 ],
   alphaCSR[ 224 ][ 251 ],
   alphaCSR[ 224 ][ 252 ],
   alphaCSR[ 224 ][ 253 ],
   alphaCSR[ 224 ][ 254 ],
   alphaCSR[ 224 ][ 255 ],
   alphaCSR[ 224 ][ 256 ],
   alphaCSR[ 224 ][ 257 ],
   alphaCSR[ 224 ][ 258 ],
   alphaCSR[ 224 ][ 259 ],
   alphaCSR[ 224 ][ 260 ],
   alphaCSR[ 224 ][ 261 ],
   alphaCSR[ 224 ][ 262 ],
   alphaCSR[ 224 ][ 263 ],
   alphaCSR[ 224 ][ 264 ],
   alphaCSR[ 224 ][ 265 ],
   alphaCSR[ 224 ][ 266 ],
   alphaCSR[ 224 ][ 267 ],
   alphaCSR[ 224 ][ 268 ],
   alphaCSR[ 224 ][ 269 ],
   alphaCSR[ 224 ][ 270 ],
   alphaCSR[ 224 ][ 271 ],
   alphaCSR[ 224 ][ 272 ],
   alphaCSR[ 224 ][ 273 ],
   alphaCSR[ 224 ][ 274 ],
   alphaCSR[ 224 ][ 275 ],
   alphaCSR[ 224 ][ 276 ],
   alphaCSR[ 224 ][ 277 ],
   alphaCSR[ 224 ][ 278 ],
   alphaCSR[ 224 ][ 279 ],
   alphaCSR[ 224 ][ 280 ],
   alphaCSR[ 224 ][ 281 ],
   alphaCSR[ 224 ][ 282 ],
   alphaCSR[ 224 ][ 283 ],
   alphaCSR[ 224 ][ 284 ],
   alphaCSR[ 224 ][ 285 ],
   alphaCSR[ 224 ][ 286 ],
   alphaCSR[ 224 ][ 287 ],
   alphaCSR[ 224 ][ 288 ],
   alphaCSR[ 224 ][ 289 ],
   alphaCSR[ 224 ][ 290 ],
   alphaCSR[ 224 ][ 291 ],
   alphaCSR[ 224 ][ 292 ],
   alphaCSR[ 224 ][ 293 ],
   alphaCSR[ 224 ][ 294 ],
   alphaCSR[ 224 ][ 295 ],
   alphaCSR[ 224 ][ 296 ],
   alphaCSR[ 224 ][ 297 ],
   alphaCSR[ 224 ][ 298 ],
   alphaCSR[ 224 ][ 299 ],
   alphaCSR[ 224 ][ 300 ],
   alphaCSR[ 224 ][ 301 ],
   alphaCSR[ 224 ][ 302 ],
   alphaCSR[ 224 ][ 303 ],
   alphaCSR[ 224 ][ 304 ],
   alphaCSR[ 224 ][ 305 ],
   alphaCSR[ 224 ][ 306 ],
   alphaCSR[ 224 ][ 307 ],
   alphaCSR[ 224 ][ 308 ],
   alphaCSR[ 224 ][ 309 ],
   alphaCSR[ 224 ][ 310 ],
   alphaCSR[ 224 ][ 311 ],
   alphaCSR[ 224 ][ 312 ],
   alphaCSR[ 224 ][ 313 ],
   alphaCSR[ 224 ][ 314 ],
   alphaCSR[ 224 ][ 315 ],
   alphaCSR[ 224 ][ 316 ],
   alphaCSR[ 224 ][ 317 ],
   alphaCSR[ 224 ][ 318 ],
   alphaCSR[ 224 ][ 319 ],
   alphaCSR[ 224 ][ 320 ],
   alphaCSR[ 224 ][ 321 ],
   alphaCSR[ 224 ][ 322 ],
   alphaCSR[ 224 ][ 323 ],
   alphaCSR[ 224 ][ 324 ],
   alphaCSR[ 224 ][ 325 ],
   alphaCSR[ 224 ][ 326 ],
   alphaCSR[ 224 ][ 327 ],
   alphaCSR[ 224 ][ 328 ],
   alphaCSR[ 224 ][ 329 ],
   alphaCSR[ 224 ][ 330 ],
   alphaCSR[ 224 ][ 331 ],
   alphaCSR[ 224 ][ 332 ],
   alphaCSR[ 224 ][ 333 ],
   alphaCSR[ 224 ][ 334 ],
   alphaCSR[ 224 ][ 335 ],
   alphaCSR[ 224 ][ 336 ],
   alphaCSR[ 224 ][ 337 ],
   alphaCSR[ 224 ][ 338 ],
   alphaCSR[ 224 ][ 339 ],
   alphaCSR[ 224 ][ 340 ],
   alphaCSR[ 224 ][ 341 ],
   alphaCSR[ 224 ][ 342 ],
   alphaCSR[ 224 ][ 343 ],
   alphaCSR[ 224 ][ 344 ],
   alphaCSR[ 224 ][ 345 ],
   alphaCSR[ 224 ][ 346 ],
   alphaCSR[ 224 ][ 347 ],
   alphaCSR[ 224 ][ 348 ],
   alphaCSR[ 224 ][ 349 ],
   alphaCSR[ 224 ][ 350 ],
   alphaCSR[ 224 ][ 351 ],
   alphaCSR[ 224 ][ 352 ],
   alphaCSR[ 224 ][ 353 ],
   alphaCSR[ 224 ][ 354 ],
   alphaCSR[ 224 ][ 355 ],
   alphaCSR[ 224 ][ 356 ],
   alphaCSR[ 224 ][ 357 ],
   alphaCSR[ 224 ][ 358 ],
   alphaCSR[ 224 ][ 359 ],
   alphaCSR[ 224 ][ 360 ],
   alphaCSR[ 224 ][ 361 ],
   alphaCSR[ 224 ][ 362 ],
   alphaCSR[ 224 ][ 363 ],
   alphaCSR[ 224 ][ 364 ],
   alphaCSR[ 224 ][ 365 ],
   alphaCSR[ 224 ][ 366 ],
   alphaCSR[ 224 ][ 367 ],
   alphaCSR[ 224 ][ 368 ],
   alphaCSR[ 224 ][ 369 ],
   alphaCSR[ 224 ][ 370 ],
   alphaCSR[ 224 ][ 371 ],
   alphaCSR[ 224 ][ 372 ],
   alphaCSR[ 224 ][ 373 ],
   alphaCSR[ 224 ][ 374 ],
   alphaCSR[ 224 ][ 375 ],
   alphaCSR[ 224 ][ 376 ],
   alphaCSR[ 224 ][ 377 ],
   alphaCSR[ 224 ][ 378 ],
   alphaCSR[ 224 ][ 379 ],
   alphaCSR[ 224 ][ 380 ],
   alphaCSR[ 224 ][ 381 ],
   alphaCSR[ 224 ][ 382 ],
   alphaCSR[ 224 ][ 383 ],
   alphaCSR[ 225 ][ 0 ],
   alphaCSR[ 225 ][ 1 ],
   alphaCSR[ 225 ][ 2 ],
   alphaCSR[ 225 ][ 3 ],
   alphaCSR[ 225 ][ 4 ],
   alphaCSR[ 225 ][ 5 ],
   alphaCSR[ 225 ][ 6 ],
   alphaCSR[ 225 ][ 7 ],
   alphaCSR[ 225 ][ 8 ],
   alphaCSR[ 225 ][ 9 ],
   alphaCSR[ 225 ][ 10 ],
   alphaCSR[ 225 ][ 11 ],
   alphaCSR[ 225 ][ 12 ],
   alphaCSR[ 225 ][ 13 ],
   alphaCSR[ 225 ][ 14 ],
   alphaCSR[ 225 ][ 15 ],
   alphaCSR[ 225 ][ 16 ],
   alphaCSR[ 225 ][ 17 ],
   alphaCSR[ 225 ][ 18 ],
   alphaCSR[ 225 ][ 19 ],
   alphaCSR[ 225 ][ 20 ],
   alphaCSR[ 225 ][ 21 ],
   alphaCSR[ 225 ][ 22 ],
   alphaCSR[ 225 ][ 23 ],
   alphaCSR[ 225 ][ 24 ],
   alphaCSR[ 225 ][ 25 ],
   alphaCSR[ 225 ][ 26 ],
   alphaCSR[ 225 ][ 27 ],
   alphaCSR[ 225 ][ 28 ],
   alphaCSR[ 225 ][ 29 ],
   alphaCSR[ 225 ][ 30 ],
   alphaCSR[ 225 ][ 31 ],
   alphaCSR[ 225 ][ 32 ],
   alphaCSR[ 225 ][ 33 ],
   alphaCSR[ 225 ][ 34 ],
   alphaCSR[ 225 ][ 35 ],
   alphaCSR[ 225 ][ 36 ],
   alphaCSR[ 225 ][ 37 ],
   alphaCSR[ 225 ][ 38 ],
   alphaCSR[ 225 ][ 39 ],
   alphaCSR[ 225 ][ 40 ],
   alphaCSR[ 225 ][ 41 ],
   alphaCSR[ 225 ][ 42 ],
   alphaCSR[ 225 ][ 43 ],
   alphaCSR[ 225 ][ 44 ],
   alphaCSR[ 225 ][ 45 ],
   alphaCSR[ 225 ][ 46 ],
   alphaCSR[ 225 ][ 47 ],
   alphaCSR[ 225 ][ 48 ],
   alphaCSR[ 225 ][ 49 ],
   alphaCSR[ 225 ][ 50 ],
   alphaCSR[ 225 ][ 51 ],
   alphaCSR[ 225 ][ 52 ],
   alphaCSR[ 225 ][ 53 ],
   alphaCSR[ 225 ][ 54 ],
   alphaCSR[ 225 ][ 55 ],
   alphaCSR[ 225 ][ 56 ],
   alphaCSR[ 225 ][ 57 ],
   alphaCSR[ 225 ][ 58 ],
   alphaCSR[ 225 ][ 59 ],
   alphaCSR[ 225 ][ 60 ],
   alphaCSR[ 225 ][ 61 ],
   alphaCSR[ 225 ][ 62 ],
   alphaCSR[ 225 ][ 63 ],
   alphaCSR[ 225 ][ 64 ],
   alphaCSR[ 225 ][ 65 ],
   alphaCSR[ 225 ][ 66 ],
   alphaCSR[ 225 ][ 67 ],
   alphaCSR[ 225 ][ 68 ],
   alphaCSR[ 225 ][ 69 ],
   alphaCSR[ 225 ][ 70 ],
   alphaCSR[ 225 ][ 71 ],
   alphaCSR[ 225 ][ 72 ],
   alphaCSR[ 225 ][ 73 ],
   alphaCSR[ 225 ][ 74 ],
   alphaCSR[ 225 ][ 75 ],
   alphaCSR[ 225 ][ 76 ],
   alphaCSR[ 225 ][ 77 ],
   alphaCSR[ 225 ][ 78 ],
   alphaCSR[ 225 ][ 79 ],
   alphaCSR[ 225 ][ 80 ],
   alphaCSR[ 225 ][ 81 ],
   alphaCSR[ 225 ][ 82 ],
   alphaCSR[ 225 ][ 83 ],
   alphaCSR[ 225 ][ 84 ],
   alphaCSR[ 225 ][ 85 ],
   alphaCSR[ 225 ][ 86 ],
   alphaCSR[ 225 ][ 87 ],
   alphaCSR[ 225 ][ 88 ],
   alphaCSR[ 225 ][ 89 ],
   alphaCSR[ 225 ][ 90 ],
   alphaCSR[ 225 ][ 91 ],
   alphaCSR[ 225 ][ 92 ],
   alphaCSR[ 225 ][ 93 ],
   alphaCSR[ 225 ][ 94 ],
   alphaCSR[ 225 ][ 95 ],
   alphaCSR[ 225 ][ 96 ],
   alphaCSR[ 225 ][ 97 ],
   alphaCSR[ 225 ][ 98 ],
   alphaCSR[ 225 ][ 99 ],
   alphaCSR[ 225 ][ 100 ],
   alphaCSR[ 225 ][ 101 ],
   alphaCSR[ 225 ][ 102 ],
   alphaCSR[ 225 ][ 103 ],
   alphaCSR[ 225 ][ 104 ],
   alphaCSR[ 225 ][ 105 ],
   alphaCSR[ 225 ][ 106 ],
   alphaCSR[ 225 ][ 107 ],
   alphaCSR[ 225 ][ 108 ],
   alphaCSR[ 225 ][ 109 ],
   alphaCSR[ 225 ][ 110 ],
   alphaCSR[ 225 ][ 111 ],
   alphaCSR[ 225 ][ 112 ],
   alphaCSR[ 225 ][ 113 ],
   alphaCSR[ 225 ][ 114 ],
   alphaCSR[ 225 ][ 115 ],
   alphaCSR[ 225 ][ 116 ],
   alphaCSR[ 225 ][ 117 ],
   alphaCSR[ 225 ][ 118 ],
   alphaCSR[ 225 ][ 119 ],
   alphaCSR[ 225 ][ 120 ],
   alphaCSR[ 225 ][ 121 ],
   alphaCSR[ 225 ][ 122 ],
   alphaCSR[ 225 ][ 123 ],
   alphaCSR[ 225 ][ 124 ],
   alphaCSR[ 225 ][ 125 ],
   alphaCSR[ 225 ][ 126 ],
   alphaCSR[ 225 ][ 127 ],
   alphaCSR[ 225 ][ 128 ],
   alphaCSR[ 225 ][ 129 ],
   alphaCSR[ 225 ][ 130 ],
   alphaCSR[ 225 ][ 131 ],
   alphaCSR[ 225 ][ 132 ],
   alphaCSR[ 225 ][ 133 ],
   alphaCSR[ 225 ][ 134 ],
   alphaCSR[ 225 ][ 135 ],
   alphaCSR[ 225 ][ 136 ],
   alphaCSR[ 225 ][ 137 ],
   alphaCSR[ 225 ][ 138 ],
   alphaCSR[ 225 ][ 139 ],
   alphaCSR[ 225 ][ 140 ],
   alphaCSR[ 225 ][ 141 ],
   alphaCSR[ 225 ][ 142 ],
   alphaCSR[ 225 ][ 143 ],
   alphaCSR[ 225 ][ 144 ],
   alphaCSR[ 225 ][ 145 ],
   alphaCSR[ 225 ][ 146 ],
   alphaCSR[ 225 ][ 147 ],
   alphaCSR[ 225 ][ 148 ],
   alphaCSR[ 225 ][ 149 ],
   alphaCSR[ 225 ][ 150 ],
   alphaCSR[ 225 ][ 151 ],
   alphaCSR[ 225 ][ 152 ],
   alphaCSR[ 225 ][ 153 ],
   alphaCSR[ 225 ][ 154 ],
   alphaCSR[ 225 ][ 155 ],
   alphaCSR[ 225 ][ 156 ],
   alphaCSR[ 225 ][ 157 ],
   alphaCSR[ 225 ][ 158 ],
   alphaCSR[ 225 ][ 159 ],
   alphaCSR[ 225 ][ 160 ],
   alphaCSR[ 225 ][ 161 ],
   alphaCSR[ 225 ][ 162 ],
   alphaCSR[ 225 ][ 163 ],
   alphaCSR[ 225 ][ 164 ],
   alphaCSR[ 225 ][ 165 ],
   alphaCSR[ 225 ][ 166 ],
   alphaCSR[ 225 ][ 167 ],
   alphaCSR[ 225 ][ 168 ],
   alphaCSR[ 225 ][ 169 ],
   alphaCSR[ 225 ][ 170 ],
   alphaCSR[ 225 ][ 171 ],
   alphaCSR[ 225 ][ 172 ],
   alphaCSR[ 225 ][ 173 ],
   alphaCSR[ 225 ][ 174 ],
   alphaCSR[ 225 ][ 175 ],
   alphaCSR[ 225 ][ 176 ],
   alphaCSR[ 225 ][ 177 ],
   alphaCSR[ 225 ][ 178 ],
   alphaCSR[ 225 ][ 179 ],
   alphaCSR[ 225 ][ 180 ],
   alphaCSR[ 225 ][ 181 ],
   alphaCSR[ 225 ][ 182 ],
   alphaCSR[ 225 ][ 183 ],
   alphaCSR[ 225 ][ 184 ],
   alphaCSR[ 225 ][ 185 ],
   alphaCSR[ 225 ][ 186 ],
   alphaCSR[ 225 ][ 187 ],
   alphaCSR[ 225 ][ 188 ],
   alphaCSR[ 225 ][ 189 ],
   alphaCSR[ 225 ][ 190 ],
   alphaCSR[ 225 ][ 191 ],
   alphaCSR[ 225 ][ 192 ],
   alphaCSR[ 225 ][ 193 ],
   alphaCSR[ 225 ][ 194 ],
   alphaCSR[ 225 ][ 195 ],
   alphaCSR[ 225 ][ 196 ],
   alphaCSR[ 225 ][ 197 ],
   alphaCSR[ 225 ][ 198 ],
   alphaCSR[ 225 ][ 199 ],
   alphaCSR[ 225 ][ 200 ],
   alphaCSR[ 225 ][ 201 ],
   alphaCSR[ 225 ][ 202 ],
   alphaCSR[ 225 ][ 203 ],
   alphaCSR[ 225 ][ 204 ],
   alphaCSR[ 225 ][ 205 ],
   alphaCSR[ 225 ][ 206 ],
   alphaCSR[ 225 ][ 207 ],
   alphaCSR[ 225 ][ 208 ],
   alphaCSR[ 225 ][ 209 ],
   alphaCSR[ 225 ][ 210 ],
   alphaCSR[ 225 ][ 211 ],
   alphaCSR[ 225 ][ 212 ],
   alphaCSR[ 225 ][ 213 ],
   alphaCSR[ 225 ][ 214 ],
   alphaCSR[ 225 ][ 215 ],
   alphaCSR[ 225 ][ 216 ],
   alphaCSR[ 225 ][ 217 ],
   alphaCSR[ 225 ][ 218 ],
   alphaCSR[ 225 ][ 219 ],
   alphaCSR[ 225 ][ 220 ],
   alphaCSR[ 225 ][ 221 ],
   alphaCSR[ 225 ][ 222 ],
   alphaCSR[ 225 ][ 223 ],
   alphaCSR[ 225 ][ 224 ],
   alphaCSR[ 225 ][ 225 ],
   alphaCSR[ 225 ][ 226 ],
   alphaCSR[ 225 ][ 227 ],
   alphaCSR[ 225 ][ 228 ],
   alphaCSR[ 225 ][ 229 ],
   alphaCSR[ 225 ][ 230 ],
   alphaCSR[ 225 ][ 231 ],
   alphaCSR[ 225 ][ 232 ],
   alphaCSR[ 225 ][ 233 ],
   alphaCSR[ 225 ][ 234 ],
   alphaCSR[ 225 ][ 235 ],
   alphaCSR[ 225 ][ 236 ],
   alphaCSR[ 225 ][ 237 ],
   alphaCSR[ 225 ][ 238 ],
   alphaCSR[ 225 ][ 239 ],
   alphaCSR[ 225 ][ 240 ],
   alphaCSR[ 225 ][ 241 ],
   alphaCSR[ 225 ][ 242 ],
   alphaCSR[ 225 ][ 243 ],
   alphaCSR[ 225 ][ 244 ],
   alphaCSR[ 225 ][ 245 ],
   alphaCSR[ 225 ][ 246 ],
   alphaCSR[ 225 ][ 247 ],
   alphaCSR[ 225 ][ 248 ],
   alphaCSR[ 225 ][ 249 ],
   alphaCSR[ 225 ][ 250 ],
   alphaCSR[ 225 ][ 251 ],
   alphaCSR[ 225 ][ 252 ],
   alphaCSR[ 225 ][ 253 ],
   alphaCSR[ 225 ][ 254 ],
   alphaCSR[ 225 ][ 255 ],
   alphaCSR[ 225 ][ 256 ],
   alphaCSR[ 225 ][ 257 ],
   alphaCSR[ 225 ][ 258 ],
   alphaCSR[ 225 ][ 259 ],
   alphaCSR[ 225 ][ 260 ],
   alphaCSR[ 225 ][ 261 ],
   alphaCSR[ 225 ][ 262 ],
   alphaCSR[ 225 ][ 263 ],
   alphaCSR[ 225 ][ 264 ],
   alphaCSR[ 225 ][ 265 ],
   alphaCSR[ 225 ][ 266 ],
   alphaCSR[ 225 ][ 267 ],
   alphaCSR[ 225 ][ 268 ],
   alphaCSR[ 225 ][ 269 ],
   alphaCSR[ 225 ][ 270 ],
   alphaCSR[ 225 ][ 271 ],
   alphaCSR[ 225 ][ 272 ],
   alphaCSR[ 225 ][ 273 ],
   alphaCSR[ 225 ][ 274 ],
   alphaCSR[ 225 ][ 275 ],
   alphaCSR[ 225 ][ 276 ],
   alphaCSR[ 225 ][ 277 ],
   alphaCSR[ 225 ][ 278 ],
   alphaCSR[ 225 ][ 279 ],
   alphaCSR[ 225 ][ 280 ],
   alphaCSR[ 225 ][ 281 ],
   alphaCSR[ 225 ][ 282 ],
   alphaCSR[ 225 ][ 283 ],
   alphaCSR[ 225 ][ 284 ],
   alphaCSR[ 225 ][ 285 ],
   alphaCSR[ 225 ][ 286 ],
   alphaCSR[ 225 ][ 287 ],
   alphaCSR[ 225 ][ 288 ],
   alphaCSR[ 225 ][ 289 ],
   alphaCSR[ 225 ][ 290 ],
   alphaCSR[ 225 ][ 291 ],
   alphaCSR[ 225 ][ 292 ],
   alphaCSR[ 225 ][ 293 ],
   alphaCSR[ 225 ][ 294 ],
   alphaCSR[ 225 ][ 295 ],
   alphaCSR[ 225 ][ 296 ],
   alphaCSR[ 225 ][ 297 ],
   alphaCSR[ 225 ][ 298 ],
   alphaCSR[ 225 ][ 299 ],
   alphaCSR[ 225 ][ 300 ],
   alphaCSR[ 225 ][ 301 ],
   alphaCSR[ 225 ][ 302 ],
   alphaCSR[ 225 ][ 303 ],
   alphaCSR[ 225 ][ 304 ],
   alphaCSR[ 225 ][ 305 ],
   alphaCSR[ 225 ][ 306 ],
   alphaCSR[ 225 ][ 307 ],
   alphaCSR[ 225 ][ 308 ],
   alphaCSR[ 225 ][ 309 ],
   alphaCSR[ 225 ][ 310 ],
   alphaCSR[ 225 ][ 311 ],
   alphaCSR[ 225 ][ 312 ],
   alphaCSR[ 225 ][ 313 ],
   alphaCSR[ 225 ][ 314 ],
   alphaCSR[ 225 ][ 315 ],
   alphaCSR[ 225 ][ 316 ],
   alphaCSR[ 225 ][ 317 ],
   alphaCSR[ 225 ][ 318 ],
   alphaCSR[ 225 ][ 319 ],
   alphaCSR[ 225 ][ 320 ],
   alphaCSR[ 225 ][ 321 ],
   alphaCSR[ 225 ][ 322 ],
   alphaCSR[ 225 ][ 323 ],
   alphaCSR[ 225 ][ 324 ],
   alphaCSR[ 225 ][ 325 ],
   alphaCSR[ 225 ][ 326 ],
   alphaCSR[ 225 ][ 327 ],
   alphaCSR[ 225 ][ 328 ],
   alphaCSR[ 225 ][ 329 ],
   alphaCSR[ 225 ][ 330 ],
   alphaCSR[ 225 ][ 331 ],
   alphaCSR[ 225 ][ 332 ],
   alphaCSR[ 225 ][ 333 ],
   alphaCSR[ 225 ][ 334 ],
   alphaCSR[ 225 ][ 335 ],
   alphaCSR[ 225 ][ 336 ],
   alphaCSR[ 225 ][ 337 ],
   alphaCSR[ 225 ][ 338 ],
   alphaCSR[ 225 ][ 339 ],
   alphaCSR[ 225 ][ 340 ],
   alphaCSR[ 225 ][ 341 ],
   alphaCSR[ 225 ][ 342 ],
   alphaCSR[ 225 ][ 343 ],
   alphaCSR[ 225 ][ 344 ],
   alphaCSR[ 225 ][ 345 ],
   alphaCSR[ 225 ][ 346 ],
   alphaCSR[ 225 ][ 347 ],
   alphaCSR[ 225 ][ 348 ],
   alphaCSR[ 225 ][ 349 ],
   alphaCSR[ 225 ][ 350 ],
   alphaCSR[ 225 ][ 351 ],
   alphaCSR[ 225 ][ 352 ],
   alphaCSR[ 225 ][ 353 ],
   alphaCSR[ 225 ][ 354 ],
   alphaCSR[ 225 ][ 355 ],
   alphaCSR[ 225 ][ 356 ],
   alphaCSR[ 225 ][ 357 ],
   alphaCSR[ 225 ][ 358 ],
   alphaCSR[ 225 ][ 359 ],
   alphaCSR[ 225 ][ 360 ],
   alphaCSR[ 225 ][ 361 ],
   alphaCSR[ 225 ][ 362 ],
   alphaCSR[ 225 ][ 363 ],
   alphaCSR[ 225 ][ 364 ],
   alphaCSR[ 225 ][ 365 ],
   alphaCSR[ 225 ][ 366 ],
   alphaCSR[ 225 ][ 367 ],
   alphaCSR[ 225 ][ 368 ],
   alphaCSR[ 225 ][ 369 ],
   alphaCSR[ 225 ][ 370 ],
   alphaCSR[ 225 ][ 371 ],
   alphaCSR[ 225 ][ 372 ],
   alphaCSR[ 225 ][ 373 ],
   alphaCSR[ 225 ][ 374 ],
   alphaCSR[ 225 ][ 375 ],
   alphaCSR[ 225 ][ 376 ],
   alphaCSR[ 225 ][ 377 ],
   alphaCSR[ 225 ][ 378 ],
   alphaCSR[ 225 ][ 379 ],
   alphaCSR[ 225 ][ 380 ],
   alphaCSR[ 225 ][ 381 ],
   alphaCSR[ 225 ][ 382 ],
   alphaCSR[ 225 ][ 383 ],
   alphaCSR[ 226 ][ 0 ],
   alphaCSR[ 226 ][ 1 ],
   alphaCSR[ 226 ][ 2 ],
   alphaCSR[ 226 ][ 3 ],
   alphaCSR[ 226 ][ 4 ],
   alphaCSR[ 226 ][ 5 ],
   alphaCSR[ 226 ][ 6 ],
   alphaCSR[ 226 ][ 7 ],
   alphaCSR[ 226 ][ 8 ],
   alphaCSR[ 226 ][ 9 ],
   alphaCSR[ 226 ][ 10 ],
   alphaCSR[ 226 ][ 11 ],
   alphaCSR[ 226 ][ 12 ],
   alphaCSR[ 226 ][ 13 ],
   alphaCSR[ 226 ][ 14 ],
   alphaCSR[ 226 ][ 15 ],
   alphaCSR[ 226 ][ 16 ],
   alphaCSR[ 226 ][ 17 ],
   alphaCSR[ 226 ][ 18 ],
   alphaCSR[ 226 ][ 19 ],
   alphaCSR[ 226 ][ 20 ],
   alphaCSR[ 226 ][ 21 ],
   alphaCSR[ 226 ][ 22 ],
   alphaCSR[ 226 ][ 23 ],
   alphaCSR[ 226 ][ 24 ],
   alphaCSR[ 226 ][ 25 ],
   alphaCSR[ 226 ][ 26 ],
   alphaCSR[ 226 ][ 27 ],
   alphaCSR[ 226 ][ 28 ],
   alphaCSR[ 226 ][ 29 ],
   alphaCSR[ 226 ][ 30 ],
   alphaCSR[ 226 ][ 31 ],
   alphaCSR[ 226 ][ 32 ],
   alphaCSR[ 226 ][ 33 ],
   alphaCSR[ 226 ][ 34 ],
   alphaCSR[ 226 ][ 35 ],
   alphaCSR[ 226 ][ 36 ],
   alphaCSR[ 226 ][ 37 ],
   alphaCSR[ 226 ][ 38 ],
   alphaCSR[ 226 ][ 39 ],
   alphaCSR[ 226 ][ 40 ],
   alphaCSR[ 226 ][ 41 ],
   alphaCSR[ 226 ][ 42 ],
   alphaCSR[ 226 ][ 43 ],
   alphaCSR[ 226 ][ 44 ],
   alphaCSR[ 226 ][ 45 ],
   alphaCSR[ 226 ][ 46 ],
   alphaCSR[ 226 ][ 47 ],
   alphaCSR[ 226 ][ 48 ],
   alphaCSR[ 226 ][ 49 ],
   alphaCSR[ 226 ][ 50 ],
   alphaCSR[ 226 ][ 51 ],
   alphaCSR[ 226 ][ 52 ],
   alphaCSR[ 226 ][ 53 ],
   alphaCSR[ 226 ][ 54 ],
   alphaCSR[ 226 ][ 55 ],
   alphaCSR[ 226 ][ 56 ],
   alphaCSR[ 226 ][ 57 ],
   alphaCSR[ 226 ][ 58 ],
   alphaCSR[ 226 ][ 59 ],
   alphaCSR[ 226 ][ 60 ],
   alphaCSR[ 226 ][ 61 ],
   alphaCSR[ 226 ][ 62 ],
   alphaCSR[ 226 ][ 63 ],
   alphaCSR[ 226 ][ 64 ],
   alphaCSR[ 226 ][ 65 ],
   alphaCSR[ 226 ][ 66 ],
   alphaCSR[ 226 ][ 67 ],
   alphaCSR[ 226 ][ 68 ],
   alphaCSR[ 226 ][ 69 ],
   alphaCSR[ 226 ][ 70 ],
   alphaCSR[ 226 ][ 71 ],
   alphaCSR[ 226 ][ 72 ],
   alphaCSR[ 226 ][ 73 ],
   alphaCSR[ 226 ][ 74 ],
   alphaCSR[ 226 ][ 75 ],
   alphaCSR[ 226 ][ 76 ],
   alphaCSR[ 226 ][ 77 ],
   alphaCSR[ 226 ][ 78 ],
   alphaCSR[ 226 ][ 79 ],
   alphaCSR[ 226 ][ 80 ],
   alphaCSR[ 226 ][ 81 ],
   alphaCSR[ 226 ][ 82 ],
   alphaCSR[ 226 ][ 83 ],
   alphaCSR[ 226 ][ 84 ],
   alphaCSR[ 226 ][ 85 ],
   alphaCSR[ 226 ][ 86 ],
   alphaCSR[ 226 ][ 87 ],
   alphaCSR[ 226 ][ 88 ],
   alphaCSR[ 226 ][ 89 ],
   alphaCSR[ 226 ][ 90 ],
   alphaCSR[ 226 ][ 91 ],
   alphaCSR[ 226 ][ 92 ],
   alphaCSR[ 226 ][ 93 ],
   alphaCSR[ 226 ][ 94 ],
   alphaCSR[ 226 ][ 95 ],
   alphaCSR[ 226 ][ 96 ],
   alphaCSR[ 226 ][ 97 ],
   alphaCSR[ 226 ][ 98 ],
   alphaCSR[ 226 ][ 99 ],
   alphaCSR[ 226 ][ 100 ],
   alphaCSR[ 226 ][ 101 ],
   alphaCSR[ 226 ][ 102 ],
   alphaCSR[ 226 ][ 103 ],
   alphaCSR[ 226 ][ 104 ],
   alphaCSR[ 226 ][ 105 ],
   alphaCSR[ 226 ][ 106 ],
   alphaCSR[ 226 ][ 107 ],
   alphaCSR[ 226 ][ 108 ],
   alphaCSR[ 226 ][ 109 ],
   alphaCSR[ 226 ][ 110 ],
   alphaCSR[ 226 ][ 111 ],
   alphaCSR[ 226 ][ 112 ],
   alphaCSR[ 226 ][ 113 ],
   alphaCSR[ 226 ][ 114 ],
   alphaCSR[ 226 ][ 115 ],
   alphaCSR[ 226 ][ 116 ],
   alphaCSR[ 226 ][ 117 ],
   alphaCSR[ 226 ][ 118 ],
   alphaCSR[ 226 ][ 119 ],
   alphaCSR[ 226 ][ 120 ],
   alphaCSR[ 226 ][ 121 ],
   alphaCSR[ 226 ][ 122 ],
   alphaCSR[ 226 ][ 123 ],
   alphaCSR[ 226 ][ 124 ],
   alphaCSR[ 226 ][ 125 ],
   alphaCSR[ 226 ][ 126 ],
   alphaCSR[ 226 ][ 127 ],
   alphaCSR[ 226 ][ 128 ],
   alphaCSR[ 226 ][ 129 ],
   alphaCSR[ 226 ][ 130 ],
   alphaCSR[ 226 ][ 131 ],
   alphaCSR[ 226 ][ 132 ],
   alphaCSR[ 226 ][ 133 ],
   alphaCSR[ 226 ][ 134 ],
   alphaCSR[ 226 ][ 135 ],
   alphaCSR[ 226 ][ 136 ],
   alphaCSR[ 226 ][ 137 ],
   alphaCSR[ 226 ][ 138 ],
   alphaCSR[ 226 ][ 139 ],
   alphaCSR[ 226 ][ 140 ],
   alphaCSR[ 226 ][ 141 ],
   alphaCSR[ 226 ][ 142 ],
   alphaCSR[ 226 ][ 143 ],
   alphaCSR[ 226 ][ 144 ],
   alphaCSR[ 226 ][ 145 ],
   alphaCSR[ 226 ][ 146 ],
   alphaCSR[ 226 ][ 147 ],
   alphaCSR[ 226 ][ 148 ],
   alphaCSR[ 226 ][ 149 ],
   alphaCSR[ 226 ][ 150 ],
   alphaCSR[ 226 ][ 151 ],
   alphaCSR[ 226 ][ 152 ],
   alphaCSR[ 226 ][ 153 ],
   alphaCSR[ 226 ][ 154 ],
   alphaCSR[ 226 ][ 155 ],
   alphaCSR[ 226 ][ 156 ],
   alphaCSR[ 226 ][ 157 ],
   alphaCSR[ 226 ][ 158 ],
   alphaCSR[ 226 ][ 159 ],
   alphaCSR[ 226 ][ 160 ],
   alphaCSR[ 226 ][ 161 ],
   alphaCSR[ 226 ][ 162 ],
   alphaCSR[ 226 ][ 163 ],
   alphaCSR[ 226 ][ 164 ],
   alphaCSR[ 226 ][ 165 ],
   alphaCSR[ 226 ][ 166 ],
   alphaCSR[ 226 ][ 167 ],
   alphaCSR[ 226 ][ 168 ],
   alphaCSR[ 226 ][ 169 ],
   alphaCSR[ 226 ][ 170 ],
   alphaCSR[ 226 ][ 171 ],
   alphaCSR[ 226 ][ 172 ],
   alphaCSR[ 226 ][ 173 ],
   alphaCSR[ 226 ][ 174 ],
   alphaCSR[ 226 ][ 175 ],
   alphaCSR[ 226 ][ 176 ],
   alphaCSR[ 226 ][ 177 ],
   alphaCSR[ 226 ][ 178 ],
   alphaCSR[ 226 ][ 179 ],
   alphaCSR[ 226 ][ 180 ],
   alphaCSR[ 226 ][ 181 ],
   alphaCSR[ 226 ][ 182 ],
   alphaCSR[ 226 ][ 183 ],
   alphaCSR[ 226 ][ 184 ],
   alphaCSR[ 226 ][ 185 ],
   alphaCSR[ 226 ][ 186 ],
   alphaCSR[ 226 ][ 187 ],
   alphaCSR[ 226 ][ 188 ],
   alphaCSR[ 226 ][ 189 ],
   alphaCSR[ 226 ][ 190 ],
   alphaCSR[ 226 ][ 191 ],
   alphaCSR[ 226 ][ 192 ],
   alphaCSR[ 226 ][ 193 ],
   alphaCSR[ 226 ][ 194 ],
   alphaCSR[ 226 ][ 195 ],
   alphaCSR[ 226 ][ 196 ],
   alphaCSR[ 226 ][ 197 ],
   alphaCSR[ 226 ][ 198 ],
   alphaCSR[ 226 ][ 199 ],
   alphaCSR[ 226 ][ 200 ],
   alphaCSR[ 226 ][ 201 ],
   alphaCSR[ 226 ][ 202 ],
   alphaCSR[ 226 ][ 203 ],
   alphaCSR[ 226 ][ 204 ],
   alphaCSR[ 226 ][ 205 ],
   alphaCSR[ 226 ][ 206 ],
   alphaCSR[ 226 ][ 207 ],
   alphaCSR[ 226 ][ 208 ],
   alphaCSR[ 226 ][ 209 ],
   alphaCSR[ 226 ][ 210 ],
   alphaCSR[ 226 ][ 211 ],
   alphaCSR[ 226 ][ 212 ],
   alphaCSR[ 226 ][ 213 ],
   alphaCSR[ 226 ][ 214 ],
   alphaCSR[ 226 ][ 215 ],
   alphaCSR[ 226 ][ 216 ],
   alphaCSR[ 226 ][ 217 ],
   alphaCSR[ 226 ][ 218 ],
   alphaCSR[ 226 ][ 219 ],
   alphaCSR[ 226 ][ 220 ],
   alphaCSR[ 226 ][ 221 ],
   alphaCSR[ 226 ][ 222 ],
   alphaCSR[ 226 ][ 223 ],
   alphaCSR[ 226 ][ 224 ],
   alphaCSR[ 226 ][ 225 ],
   alphaCSR[ 226 ][ 226 ],
   alphaCSR[ 226 ][ 227 ],
   alphaCSR[ 226 ][ 228 ],
   alphaCSR[ 226 ][ 229 ],
   alphaCSR[ 226 ][ 230 ],
   alphaCSR[ 226 ][ 231 ],
   alphaCSR[ 226 ][ 232 ],
   alphaCSR[ 226 ][ 233 ],
   alphaCSR[ 226 ][ 234 ],
   alphaCSR[ 226 ][ 235 ],
   alphaCSR[ 226 ][ 236 ],
   alphaCSR[ 226 ][ 237 ],
   alphaCSR[ 226 ][ 238 ],
   alphaCSR[ 226 ][ 239 ],
   alphaCSR[ 226 ][ 240 ],
   alphaCSR[ 226 ][ 241 ],
   alphaCSR[ 226 ][ 242 ],
   alphaCSR[ 226 ][ 243 ],
   alphaCSR[ 226 ][ 244 ],
   alphaCSR[ 226 ][ 245 ],
   alphaCSR[ 226 ][ 246 ],
   alphaCSR[ 226 ][ 247 ],
   alphaCSR[ 226 ][ 248 ],
   alphaCSR[ 226 ][ 249 ],
   alphaCSR[ 226 ][ 250 ],
   alphaCSR[ 226 ][ 251 ],
   alphaCSR[ 226 ][ 252 ],
   alphaCSR[ 226 ][ 253 ],
   alphaCSR[ 226 ][ 254 ],
   alphaCSR[ 226 ][ 255 ],
   alphaCSR[ 226 ][ 256 ],
   alphaCSR[ 226 ][ 257 ],
   alphaCSR[ 226 ][ 258 ],
   alphaCSR[ 226 ][ 259 ],
   alphaCSR[ 226 ][ 260 ],
   alphaCSR[ 226 ][ 261 ],
   alphaCSR[ 226 ][ 262 ],
   alphaCSR[ 226 ][ 263 ],
   alphaCSR[ 226 ][ 264 ],
   alphaCSR[ 226 ][ 265 ],
   alphaCSR[ 226 ][ 266 ],
   alphaCSR[ 226 ][ 267 ],
   alphaCSR[ 226 ][ 268 ],
   alphaCSR[ 226 ][ 269 ],
   alphaCSR[ 226 ][ 270 ],
   alphaCSR[ 226 ][ 271 ],
   alphaCSR[ 226 ][ 272 ],
   alphaCSR[ 226 ][ 273 ],
   alphaCSR[ 226 ][ 274 ],
   alphaCSR[ 226 ][ 275 ],
   alphaCSR[ 226 ][ 276 ],
   alphaCSR[ 226 ][ 277 ],
   alphaCSR[ 226 ][ 278 ],
   alphaCSR[ 226 ][ 279 ],
   alphaCSR[ 226 ][ 280 ],
   alphaCSR[ 226 ][ 281 ],
   alphaCSR[ 226 ][ 282 ],
   alphaCSR[ 226 ][ 283 ],
   alphaCSR[ 226 ][ 284 ],
   alphaCSR[ 226 ][ 285 ],
   alphaCSR[ 226 ][ 286 ],
   alphaCSR[ 226 ][ 287 ],
   alphaCSR[ 226 ][ 288 ],
   alphaCSR[ 226 ][ 289 ],
   alphaCSR[ 226 ][ 290 ],
   alphaCSR[ 226 ][ 291 ],
   alphaCSR[ 226 ][ 292 ],
   alphaCSR[ 226 ][ 293 ],
   alphaCSR[ 226 ][ 294 ],
   alphaCSR[ 226 ][ 295 ],
   alphaCSR[ 226 ][ 296 ],
   alphaCSR[ 226 ][ 297 ],
   alphaCSR[ 226 ][ 298 ],
   alphaCSR[ 226 ][ 299 ],
   alphaCSR[ 226 ][ 300 ],
   alphaCSR[ 226 ][ 301 ],
   alphaCSR[ 226 ][ 302 ],
   alphaCSR[ 226 ][ 303 ],
   alphaCSR[ 226 ][ 304 ],
   alphaCSR[ 226 ][ 305 ],
   alphaCSR[ 226 ][ 306 ],
   alphaCSR[ 226 ][ 307 ],
   alphaCSR[ 226 ][ 308 ],
   alphaCSR[ 226 ][ 309 ],
   alphaCSR[ 226 ][ 310 ],
   alphaCSR[ 226 ][ 311 ],
   alphaCSR[ 226 ][ 312 ],
   alphaCSR[ 226 ][ 313 ],
   alphaCSR[ 226 ][ 314 ],
   alphaCSR[ 226 ][ 315 ],
   alphaCSR[ 226 ][ 316 ],
   alphaCSR[ 226 ][ 317 ],
   alphaCSR[ 226 ][ 318 ],
   alphaCSR[ 226 ][ 319 ],
   alphaCSR[ 226 ][ 320 ],
   alphaCSR[ 226 ][ 321 ],
   alphaCSR[ 226 ][ 322 ],
   alphaCSR[ 226 ][ 323 ],
   alphaCSR[ 226 ][ 324 ],
   alphaCSR[ 226 ][ 325 ],
   alphaCSR[ 226 ][ 326 ],
   alphaCSR[ 226 ][ 327 ],
   alphaCSR[ 226 ][ 328 ],
   alphaCSR[ 226 ][ 329 ],
   alphaCSR[ 226 ][ 330 ],
   alphaCSR[ 226 ][ 331 ],
   alphaCSR[ 226 ][ 332 ],
   alphaCSR[ 226 ][ 333 ],
   alphaCSR[ 226 ][ 334 ],
   alphaCSR[ 226 ][ 335 ],
   alphaCSR[ 226 ][ 336 ],
   alphaCSR[ 226 ][ 337 ],
   alphaCSR[ 226 ][ 338 ],
   alphaCSR[ 226 ][ 339 ],
   alphaCSR[ 226 ][ 340 ],
   alphaCSR[ 226 ][ 341 ],
   alphaCSR[ 226 ][ 342 ],
   alphaCSR[ 226 ][ 343 ],
   alphaCSR[ 226 ][ 344 ],
   alphaCSR[ 226 ][ 345 ],
   alphaCSR[ 226 ][ 346 ],
   alphaCSR[ 226 ][ 347 ],
   alphaCSR[ 226 ][ 348 ],
   alphaCSR[ 226 ][ 349 ],
   alphaCSR[ 226 ][ 350 ],
   alphaCSR[ 226 ][ 351 ],
   alphaCSR[ 226 ][ 352 ],
   alphaCSR[ 226 ][ 353 ],
   alphaCSR[ 226 ][ 354 ],
   alphaCSR[ 226 ][ 355 ],
   alphaCSR[ 226 ][ 356 ],
   alphaCSR[ 226 ][ 357 ],
   alphaCSR[ 226 ][ 358 ],
   alphaCSR[ 226 ][ 359 ],
   alphaCSR[ 226 ][ 360 ],
   alphaCSR[ 226 ][ 361 ],
   alphaCSR[ 226 ][ 362 ],
   alphaCSR[ 226 ][ 363 ],
   alphaCSR[ 226 ][ 364 ],
   alphaCSR[ 226 ][ 365 ],
   alphaCSR[ 226 ][ 366 ],
   alphaCSR[ 226 ][ 367 ],
   alphaCSR[ 226 ][ 368 ],
   alphaCSR[ 226 ][ 369 ],
   alphaCSR[ 226 ][ 370 ],
   alphaCSR[ 226 ][ 371 ],
   alphaCSR[ 226 ][ 372 ],
   alphaCSR[ 226 ][ 373 ],
   alphaCSR[ 226 ][ 374 ],
   alphaCSR[ 226 ][ 375 ],
   alphaCSR[ 226 ][ 376 ],
   alphaCSR[ 226 ][ 377 ],
   alphaCSR[ 226 ][ 378 ],
   alphaCSR[ 226 ][ 379 ],
   alphaCSR[ 226 ][ 380 ],
   alphaCSR[ 226 ][ 381 ],
   alphaCSR[ 226 ][ 382 ],
   alphaCSR[ 226 ][ 383 ],
   alphaCSR[ 227 ][ 0 ],
   alphaCSR[ 227 ][ 1 ],
   alphaCSR[ 227 ][ 2 ],
   alphaCSR[ 227 ][ 3 ],
   alphaCSR[ 227 ][ 4 ],
   alphaCSR[ 227 ][ 5 ],
   alphaCSR[ 227 ][ 6 ],
   alphaCSR[ 227 ][ 7 ],
   alphaCSR[ 227 ][ 8 ],
   alphaCSR[ 227 ][ 9 ],
   alphaCSR[ 227 ][ 10 ],
   alphaCSR[ 227 ][ 11 ],
   alphaCSR[ 227 ][ 12 ],
   alphaCSR[ 227 ][ 13 ],
   alphaCSR[ 227 ][ 14 ],
   alphaCSR[ 227 ][ 15 ],
   alphaCSR[ 227 ][ 16 ],
   alphaCSR[ 227 ][ 17 ],
   alphaCSR[ 227 ][ 18 ],
   alphaCSR[ 227 ][ 19 ],
   alphaCSR[ 227 ][ 20 ],
   alphaCSR[ 227 ][ 21 ],
   alphaCSR[ 227 ][ 22 ],
   alphaCSR[ 227 ][ 23 ],
   alphaCSR[ 227 ][ 24 ],
   alphaCSR[ 227 ][ 25 ],
   alphaCSR[ 227 ][ 26 ],
   alphaCSR[ 227 ][ 27 ],
   alphaCSR[ 227 ][ 28 ],
   alphaCSR[ 227 ][ 29 ],
   alphaCSR[ 227 ][ 30 ],
   alphaCSR[ 227 ][ 31 ],
   alphaCSR[ 227 ][ 32 ],
   alphaCSR[ 227 ][ 33 ],
   alphaCSR[ 227 ][ 34 ],
   alphaCSR[ 227 ][ 35 ],
   alphaCSR[ 227 ][ 36 ],
   alphaCSR[ 227 ][ 37 ],
   alphaCSR[ 227 ][ 38 ],
   alphaCSR[ 227 ][ 39 ],
   alphaCSR[ 227 ][ 40 ],
   alphaCSR[ 227 ][ 41 ],
   alphaCSR[ 227 ][ 42 ],
   alphaCSR[ 227 ][ 43 ],
   alphaCSR[ 227 ][ 44 ],
   alphaCSR[ 227 ][ 45 ],
   alphaCSR[ 227 ][ 46 ],
   alphaCSR[ 227 ][ 47 ],
   alphaCSR[ 227 ][ 48 ],
   alphaCSR[ 227 ][ 49 ],
   alphaCSR[ 227 ][ 50 ],
   alphaCSR[ 227 ][ 51 ],
   alphaCSR[ 227 ][ 52 ],
   alphaCSR[ 227 ][ 53 ],
   alphaCSR[ 227 ][ 54 ],
   alphaCSR[ 227 ][ 55 ],
   alphaCSR[ 227 ][ 56 ],
   alphaCSR[ 227 ][ 57 ],
   alphaCSR[ 227 ][ 58 ],
   alphaCSR[ 227 ][ 59 ],
   alphaCSR[ 227 ][ 60 ],
   alphaCSR[ 227 ][ 61 ],
   alphaCSR[ 227 ][ 62 ],
   alphaCSR[ 227 ][ 63 ],
   alphaCSR[ 227 ][ 64 ],
   alphaCSR[ 227 ][ 65 ],
   alphaCSR[ 227 ][ 66 ],
   alphaCSR[ 227 ][ 67 ],
   alphaCSR[ 227 ][ 68 ],
   alphaCSR[ 227 ][ 69 ],
   alphaCSR[ 227 ][ 70 ],
   alphaCSR[ 227 ][ 71 ],
   alphaCSR[ 227 ][ 72 ],
   alphaCSR[ 227 ][ 73 ],
   alphaCSR[ 227 ][ 74 ],
   alphaCSR[ 227 ][ 75 ],
   alphaCSR[ 227 ][ 76 ],
   alphaCSR[ 227 ][ 77 ],
   alphaCSR[ 227 ][ 78 ],
   alphaCSR[ 227 ][ 79 ],
   alphaCSR[ 227 ][ 80 ],
   alphaCSR[ 227 ][ 81 ],
   alphaCSR[ 227 ][ 82 ],
   alphaCSR[ 227 ][ 83 ],
   alphaCSR[ 227 ][ 84 ],
   alphaCSR[ 227 ][ 85 ],
   alphaCSR[ 227 ][ 86 ],
   alphaCSR[ 227 ][ 87 ],
   alphaCSR[ 227 ][ 88 ],
   alphaCSR[ 227 ][ 89 ],
   alphaCSR[ 227 ][ 90 ],
   alphaCSR[ 227 ][ 91 ],
   alphaCSR[ 227 ][ 92 ],
   alphaCSR[ 227 ][ 93 ],
   alphaCSR[ 227 ][ 94 ],
   alphaCSR[ 227 ][ 95 ],
   alphaCSR[ 227 ][ 96 ],
   alphaCSR[ 227 ][ 97 ],
   alphaCSR[ 227 ][ 98 ],
   alphaCSR[ 227 ][ 99 ],
   alphaCSR[ 227 ][ 100 ],
   alphaCSR[ 227 ][ 101 ],
   alphaCSR[ 227 ][ 102 ],
   alphaCSR[ 227 ][ 103 ],
   alphaCSR[ 227 ][ 104 ],
   alphaCSR[ 227 ][ 105 ],
   alphaCSR[ 227 ][ 106 ],
   alphaCSR[ 227 ][ 107 ],
   alphaCSR[ 227 ][ 108 ],
   alphaCSR[ 227 ][ 109 ],
   alphaCSR[ 227 ][ 110 ],
   alphaCSR[ 227 ][ 111 ],
   alphaCSR[ 227 ][ 112 ],
   alphaCSR[ 227 ][ 113 ],
   alphaCSR[ 227 ][ 114 ],
   alphaCSR[ 227 ][ 115 ],
   alphaCSR[ 227 ][ 116 ],
   alphaCSR[ 227 ][ 117 ],
   alphaCSR[ 227 ][ 118 ],
   alphaCSR[ 227 ][ 119 ],
   alphaCSR[ 227 ][ 120 ],
   alphaCSR[ 227 ][ 121 ],
   alphaCSR[ 227 ][ 122 ],
   alphaCSR[ 227 ][ 123 ],
   alphaCSR[ 227 ][ 124 ],
   alphaCSR[ 227 ][ 125 ],
   alphaCSR[ 227 ][ 126 ],
   alphaCSR[ 227 ][ 127 ],
   alphaCSR[ 227 ][ 128 ],
   alphaCSR[ 227 ][ 129 ],
   alphaCSR[ 227 ][ 130 ],
   alphaCSR[ 227 ][ 131 ],
   alphaCSR[ 227 ][ 132 ],
   alphaCSR[ 227 ][ 133 ],
   alphaCSR[ 227 ][ 134 ],
   alphaCSR[ 227 ][ 135 ],
   alphaCSR[ 227 ][ 136 ],
   alphaCSR[ 227 ][ 137 ],
   alphaCSR[ 227 ][ 138 ],
   alphaCSR[ 227 ][ 139 ],
   alphaCSR[ 227 ][ 140 ],
   alphaCSR[ 227 ][ 141 ],
   alphaCSR[ 227 ][ 142 ],
   alphaCSR[ 227 ][ 143 ],
   alphaCSR[ 227 ][ 144 ],
   alphaCSR[ 227 ][ 145 ],
   alphaCSR[ 227 ][ 146 ],
   alphaCSR[ 227 ][ 147 ],
   alphaCSR[ 227 ][ 148 ],
   alphaCSR[ 227 ][ 149 ],
   alphaCSR[ 227 ][ 150 ],
   alphaCSR[ 227 ][ 151 ],
   alphaCSR[ 227 ][ 152 ],
   alphaCSR[ 227 ][ 153 ],
   alphaCSR[ 227 ][ 154 ],
   alphaCSR[ 227 ][ 155 ],
   alphaCSR[ 227 ][ 156 ],
   alphaCSR[ 227 ][ 157 ],
   alphaCSR[ 227 ][ 158 ],
   alphaCSR[ 227 ][ 159 ],
   alphaCSR[ 227 ][ 160 ],
   alphaCSR[ 227 ][ 161 ],
   alphaCSR[ 227 ][ 162 ],
   alphaCSR[ 227 ][ 163 ],
   alphaCSR[ 227 ][ 164 ],
   alphaCSR[ 227 ][ 165 ],
   alphaCSR[ 227 ][ 166 ],
   alphaCSR[ 227 ][ 167 ],
   alphaCSR[ 227 ][ 168 ],
   alphaCSR[ 227 ][ 169 ],
   alphaCSR[ 227 ][ 170 ],
   alphaCSR[ 227 ][ 171 ],
   alphaCSR[ 227 ][ 172 ],
   alphaCSR[ 227 ][ 173 ],
   alphaCSR[ 227 ][ 174 ],
   alphaCSR[ 227 ][ 175 ],
   alphaCSR[ 227 ][ 176 ],
   alphaCSR[ 227 ][ 177 ],
   alphaCSR[ 227 ][ 178 ],
   alphaCSR[ 227 ][ 179 ],
   alphaCSR[ 227 ][ 180 ],
   alphaCSR[ 227 ][ 181 ],
   alphaCSR[ 227 ][ 182 ],
   alphaCSR[ 227 ][ 183 ],
   alphaCSR[ 227 ][ 184 ],
   alphaCSR[ 227 ][ 185 ],
   alphaCSR[ 227 ][ 186 ],
   alphaCSR[ 227 ][ 187 ],
   alphaCSR[ 227 ][ 188 ],
   alphaCSR[ 227 ][ 189 ],
   alphaCSR[ 227 ][ 190 ],
   alphaCSR[ 227 ][ 191 ],
   alphaCSR[ 227 ][ 192 ],
   alphaCSR[ 227 ][ 193 ],
   alphaCSR[ 227 ][ 194 ],
   alphaCSR[ 227 ][ 195 ],
   alphaCSR[ 227 ][ 196 ],
   alphaCSR[ 227 ][ 197 ],
   alphaCSR[ 227 ][ 198 ],
   alphaCSR[ 227 ][ 199 ],
   alphaCSR[ 227 ][ 200 ],
   alphaCSR[ 227 ][ 201 ],
   alphaCSR[ 227 ][ 202 ],
   alphaCSR[ 227 ][ 203 ],
   alphaCSR[ 227 ][ 204 ],
   alphaCSR[ 227 ][ 205 ],
   alphaCSR[ 227 ][ 206 ],
   alphaCSR[ 227 ][ 207 ],
   alphaCSR[ 227 ][ 208 ],
   alphaCSR[ 227 ][ 209 ],
   alphaCSR[ 227 ][ 210 ],
   alphaCSR[ 227 ][ 211 ],
   alphaCSR[ 227 ][ 212 ],
   alphaCSR[ 227 ][ 213 ],
   alphaCSR[ 227 ][ 214 ],
   alphaCSR[ 227 ][ 215 ],
   alphaCSR[ 227 ][ 216 ],
   alphaCSR[ 227 ][ 217 ],
   alphaCSR[ 227 ][ 218 ],
   alphaCSR[ 227 ][ 219 ],
   alphaCSR[ 227 ][ 220 ],
   alphaCSR[ 227 ][ 221 ],
   alphaCSR[ 227 ][ 222 ],
   alphaCSR[ 227 ][ 223 ],
   alphaCSR[ 227 ][ 224 ],
   alphaCSR[ 227 ][ 225 ],
   alphaCSR[ 227 ][ 226 ],
   alphaCSR[ 227 ][ 227 ],
   alphaCSR[ 227 ][ 228 ],
   alphaCSR[ 227 ][ 229 ],
   alphaCSR[ 227 ][ 230 ],
   alphaCSR[ 227 ][ 231 ],
   alphaCSR[ 227 ][ 232 ],
   alphaCSR[ 227 ][ 233 ],
   alphaCSR[ 227 ][ 234 ],
   alphaCSR[ 227 ][ 235 ],
   alphaCSR[ 227 ][ 236 ],
   alphaCSR[ 227 ][ 237 ],
   alphaCSR[ 227 ][ 238 ],
   alphaCSR[ 227 ][ 239 ],
   alphaCSR[ 227 ][ 240 ],
   alphaCSR[ 227 ][ 241 ],
   alphaCSR[ 227 ][ 242 ],
   alphaCSR[ 227 ][ 243 ],
   alphaCSR[ 227 ][ 244 ],
   alphaCSR[ 227 ][ 245 ],
   alphaCSR[ 227 ][ 246 ],
   alphaCSR[ 227 ][ 247 ],
   alphaCSR[ 227 ][ 248 ],
   alphaCSR[ 227 ][ 249 ],
   alphaCSR[ 227 ][ 250 ],
   alphaCSR[ 227 ][ 251 ],
   alphaCSR[ 227 ][ 252 ],
   alphaCSR[ 227 ][ 253 ],
   alphaCSR[ 227 ][ 254 ],
   alphaCSR[ 227 ][ 255 ],
   alphaCSR[ 227 ][ 256 ],
   alphaCSR[ 227 ][ 257 ],
   alphaCSR[ 227 ][ 258 ],
   alphaCSR[ 227 ][ 259 ],
   alphaCSR[ 227 ][ 260 ],
   alphaCSR[ 227 ][ 261 ],
   alphaCSR[ 227 ][ 262 ],
   alphaCSR[ 227 ][ 263 ],
   alphaCSR[ 227 ][ 264 ],
   alphaCSR[ 227 ][ 265 ],
   alphaCSR[ 227 ][ 266 ],
   alphaCSR[ 227 ][ 267 ],
   alphaCSR[ 227 ][ 268 ],
   alphaCSR[ 227 ][ 269 ],
   alphaCSR[ 227 ][ 270 ],
   alphaCSR[ 227 ][ 271 ],
   alphaCSR[ 227 ][ 272 ],
   alphaCSR[ 227 ][ 273 ],
   alphaCSR[ 227 ][ 274 ],
   alphaCSR[ 227 ][ 275 ],
   alphaCSR[ 227 ][ 276 ],
   alphaCSR[ 227 ][ 277 ],
   alphaCSR[ 227 ][ 278 ],
   alphaCSR[ 227 ][ 279 ],
   alphaCSR[ 227 ][ 280 ],
   alphaCSR[ 227 ][ 281 ],
   alphaCSR[ 227 ][ 282 ],
   alphaCSR[ 227 ][ 283 ],
   alphaCSR[ 227 ][ 284 ],
   alphaCSR[ 227 ][ 285 ],
   alphaCSR[ 227 ][ 286 ],
   alphaCSR[ 227 ][ 287 ],
   alphaCSR[ 227 ][ 288 ],
   alphaCSR[ 227 ][ 289 ],
   alphaCSR[ 227 ][ 290 ],
   alphaCSR[ 227 ][ 291 ],
   alphaCSR[ 227 ][ 292 ],
   alphaCSR[ 227 ][ 293 ],
   alphaCSR[ 227 ][ 294 ],
   alphaCSR[ 227 ][ 295 ],
   alphaCSR[ 227 ][ 296 ],
   alphaCSR[ 227 ][ 297 ],
   alphaCSR[ 227 ][ 298 ],
   alphaCSR[ 227 ][ 299 ],
   alphaCSR[ 227 ][ 300 ],
   alphaCSR[ 227 ][ 301 ],
   alphaCSR[ 227 ][ 302 ],
   alphaCSR[ 227 ][ 303 ],
   alphaCSR[ 227 ][ 304 ],
   alphaCSR[ 227 ][ 305 ],
   alphaCSR[ 227 ][ 306 ],
   alphaCSR[ 227 ][ 307 ],
   alphaCSR[ 227 ][ 308 ],
   alphaCSR[ 227 ][ 309 ],
   alphaCSR[ 227 ][ 310 ],
   alphaCSR[ 227 ][ 311 ],
   alphaCSR[ 227 ][ 312 ],
   alphaCSR[ 227 ][ 313 ],
   alphaCSR[ 227 ][ 314 ],
   alphaCSR[ 227 ][ 315 ],
   alphaCSR[ 227 ][ 316 ],
   alphaCSR[ 227 ][ 317 ],
   alphaCSR[ 227 ][ 318 ],
   alphaCSR[ 227 ][ 319 ],
   alphaCSR[ 227 ][ 320 ],
   alphaCSR[ 227 ][ 321 ],
   alphaCSR[ 227 ][ 322 ],
   alphaCSR[ 227 ][ 323 ],
   alphaCSR[ 227 ][ 324 ],
   alphaCSR[ 227 ][ 325 ],
   alphaCSR[ 227 ][ 326 ],
   alphaCSR[ 227 ][ 327 ],
   alphaCSR[ 227 ][ 328 ],
   alphaCSR[ 227 ][ 329 ],
   alphaCSR[ 227 ][ 330 ],
   alphaCSR[ 227 ][ 331 ],
   alphaCSR[ 227 ][ 332 ],
   alphaCSR[ 227 ][ 333 ],
   alphaCSR[ 227 ][ 334 ],
   alphaCSR[ 227 ][ 335 ],
   alphaCSR[ 227 ][ 336 ],
   alphaCSR[ 227 ][ 337 ],
   alphaCSR[ 227 ][ 338 ],
   alphaCSR[ 227 ][ 339 ],
   alphaCSR[ 227 ][ 340 ],
   alphaCSR[ 227 ][ 341 ],
   alphaCSR[ 227 ][ 342 ],
   alphaCSR[ 227 ][ 343 ],
   alphaCSR[ 227 ][ 344 ],
   alphaCSR[ 227 ][ 345 ],
   alphaCSR[ 227 ][ 346 ],
   alphaCSR[ 227 ][ 347 ],
   alphaCSR[ 227 ][ 348 ],
   alphaCSR[ 227 ][ 349 ],
   alphaCSR[ 227 ][ 350 ],
   alphaCSR[ 227 ][ 351 ],
   alphaCSR[ 227 ][ 352 ],
   alphaCSR[ 227 ][ 353 ],
   alphaCSR[ 227 ][ 354 ],
   alphaCSR[ 227 ][ 355 ],
   alphaCSR[ 227 ][ 356 ],
   alphaCSR[ 227 ][ 357 ],
   alphaCSR[ 227 ][ 358 ],
   alphaCSR[ 227 ][ 359 ],
   alphaCSR[ 227 ][ 360 ],
   alphaCSR[ 227 ][ 361 ],
   alphaCSR[ 227 ][ 362 ],
   alphaCSR[ 227 ][ 363 ],
   alphaCSR[ 227 ][ 364 ],
   alphaCSR[ 227 ][ 365 ],
   alphaCSR[ 227 ][ 366 ],
   alphaCSR[ 227 ][ 367 ],
   alphaCSR[ 227 ][ 368 ],
   alphaCSR[ 227 ][ 369 ],
   alphaCSR[ 227 ][ 370 ],
   alphaCSR[ 227 ][ 371 ],
   alphaCSR[ 227 ][ 372 ],
   alphaCSR[ 227 ][ 373 ],
   alphaCSR[ 227 ][ 374 ],
   alphaCSR[ 227 ][ 375 ],
   alphaCSR[ 227 ][ 376 ],
   alphaCSR[ 227 ][ 377 ],
   alphaCSR[ 227 ][ 378 ],
   alphaCSR[ 227 ][ 379 ],
   alphaCSR[ 227 ][ 380 ],
   alphaCSR[ 227 ][ 381 ],
   alphaCSR[ 227 ][ 382 ],
   alphaCSR[ 227 ][ 383 ],
   alphaCSR[ 228 ][ 0 ],
   alphaCSR[ 228 ][ 1 ],
   alphaCSR[ 228 ][ 2 ],
   alphaCSR[ 228 ][ 3 ],
   alphaCSR[ 228 ][ 4 ],
   alphaCSR[ 228 ][ 5 ],
   alphaCSR[ 228 ][ 6 ],
   alphaCSR[ 228 ][ 7 ],
   alphaCSR[ 228 ][ 8 ],
   alphaCSR[ 228 ][ 9 ],
   alphaCSR[ 228 ][ 10 ],
   alphaCSR[ 228 ][ 11 ],
   alphaCSR[ 228 ][ 12 ],
   alphaCSR[ 228 ][ 13 ],
   alphaCSR[ 228 ][ 14 ],
   alphaCSR[ 228 ][ 15 ],
   alphaCSR[ 228 ][ 16 ],
   alphaCSR[ 228 ][ 17 ],
   alphaCSR[ 228 ][ 18 ],
   alphaCSR[ 228 ][ 19 ],
   alphaCSR[ 228 ][ 20 ],
   alphaCSR[ 228 ][ 21 ],
   alphaCSR[ 228 ][ 22 ],
   alphaCSR[ 228 ][ 23 ],
   alphaCSR[ 228 ][ 24 ],
   alphaCSR[ 228 ][ 25 ],
   alphaCSR[ 228 ][ 26 ],
   alphaCSR[ 228 ][ 27 ],
   alphaCSR[ 228 ][ 28 ],
   alphaCSR[ 228 ][ 29 ],
   alphaCSR[ 228 ][ 30 ],
   alphaCSR[ 228 ][ 31 ],
   alphaCSR[ 228 ][ 32 ],
   alphaCSR[ 228 ][ 33 ],
   alphaCSR[ 228 ][ 34 ],
   alphaCSR[ 228 ][ 35 ],
   alphaCSR[ 228 ][ 36 ],
   alphaCSR[ 228 ][ 37 ],
   alphaCSR[ 228 ][ 38 ],
   alphaCSR[ 228 ][ 39 ],
   alphaCSR[ 228 ][ 40 ],
   alphaCSR[ 228 ][ 41 ],
   alphaCSR[ 228 ][ 42 ],
   alphaCSR[ 228 ][ 43 ],
   alphaCSR[ 228 ][ 44 ],
   alphaCSR[ 228 ][ 45 ],
   alphaCSR[ 228 ][ 46 ],
   alphaCSR[ 228 ][ 47 ],
   alphaCSR[ 228 ][ 48 ],
   alphaCSR[ 228 ][ 49 ],
   alphaCSR[ 228 ][ 50 ],
   alphaCSR[ 228 ][ 51 ],
   alphaCSR[ 228 ][ 52 ],
   alphaCSR[ 228 ][ 53 ],
   alphaCSR[ 228 ][ 54 ],
   alphaCSR[ 228 ][ 55 ],
   alphaCSR[ 228 ][ 56 ],
   alphaCSR[ 228 ][ 57 ],
   alphaCSR[ 228 ][ 58 ],
   alphaCSR[ 228 ][ 59 ],
   alphaCSR[ 228 ][ 60 ],
   alphaCSR[ 228 ][ 61 ],
   alphaCSR[ 228 ][ 62 ],
   alphaCSR[ 228 ][ 63 ],
   alphaCSR[ 228 ][ 64 ],
   alphaCSR[ 228 ][ 65 ],
   alphaCSR[ 228 ][ 66 ],
   alphaCSR[ 228 ][ 67 ],
   alphaCSR[ 228 ][ 68 ],
   alphaCSR[ 228 ][ 69 ],
   alphaCSR[ 228 ][ 70 ],
   alphaCSR[ 228 ][ 71 ],
   alphaCSR[ 228 ][ 72 ],
   alphaCSR[ 228 ][ 73 ],
   alphaCSR[ 228 ][ 74 ],
   alphaCSR[ 228 ][ 75 ],
   alphaCSR[ 228 ][ 76 ],
   alphaCSR[ 228 ][ 77 ],
   alphaCSR[ 228 ][ 78 ],
   alphaCSR[ 228 ][ 79 ],
   alphaCSR[ 228 ][ 80 ],
   alphaCSR[ 228 ][ 81 ],
   alphaCSR[ 228 ][ 82 ],
   alphaCSR[ 228 ][ 83 ],
   alphaCSR[ 228 ][ 84 ],
   alphaCSR[ 228 ][ 85 ],
   alphaCSR[ 228 ][ 86 ],
   alphaCSR[ 228 ][ 87 ],
   alphaCSR[ 228 ][ 88 ],
   alphaCSR[ 228 ][ 89 ],
   alphaCSR[ 228 ][ 90 ],
   alphaCSR[ 228 ][ 91 ],
   alphaCSR[ 228 ][ 92 ],
   alphaCSR[ 228 ][ 93 ],
   alphaCSR[ 228 ][ 94 ],
   alphaCSR[ 228 ][ 95 ],
   alphaCSR[ 228 ][ 96 ],
   alphaCSR[ 228 ][ 97 ],
   alphaCSR[ 228 ][ 98 ],
   alphaCSR[ 228 ][ 99 ],
   alphaCSR[ 228 ][ 100 ],
   alphaCSR[ 228 ][ 101 ],
   alphaCSR[ 228 ][ 102 ],
   alphaCSR[ 228 ][ 103 ],
   alphaCSR[ 228 ][ 104 ],
   alphaCSR[ 228 ][ 105 ],
   alphaCSR[ 228 ][ 106 ],
   alphaCSR[ 228 ][ 107 ],
   alphaCSR[ 228 ][ 108 ],
   alphaCSR[ 228 ][ 109 ],
   alphaCSR[ 228 ][ 110 ],
   alphaCSR[ 228 ][ 111 ],
   alphaCSR[ 228 ][ 112 ],
   alphaCSR[ 228 ][ 113 ],
   alphaCSR[ 228 ][ 114 ],
   alphaCSR[ 228 ][ 115 ],
   alphaCSR[ 228 ][ 116 ],
   alphaCSR[ 228 ][ 117 ],
   alphaCSR[ 228 ][ 118 ],
   alphaCSR[ 228 ][ 119 ],
   alphaCSR[ 228 ][ 120 ],
   alphaCSR[ 228 ][ 121 ],
   alphaCSR[ 228 ][ 122 ],
   alphaCSR[ 228 ][ 123 ],
   alphaCSR[ 228 ][ 124 ],
   alphaCSR[ 228 ][ 125 ],
   alphaCSR[ 228 ][ 126 ],
   alphaCSR[ 228 ][ 127 ],
   alphaCSR[ 228 ][ 128 ],
   alphaCSR[ 228 ][ 129 ],
   alphaCSR[ 228 ][ 130 ],
   alphaCSR[ 228 ][ 131 ],
   alphaCSR[ 228 ][ 132 ],
   alphaCSR[ 228 ][ 133 ],
   alphaCSR[ 228 ][ 134 ],
   alphaCSR[ 228 ][ 135 ],
   alphaCSR[ 228 ][ 136 ],
   alphaCSR[ 228 ][ 137 ],
   alphaCSR[ 228 ][ 138 ],
   alphaCSR[ 228 ][ 139 ],
   alphaCSR[ 228 ][ 140 ],
   alphaCSR[ 228 ][ 141 ],
   alphaCSR[ 228 ][ 142 ],
   alphaCSR[ 228 ][ 143 ],
   alphaCSR[ 228 ][ 144 ],
   alphaCSR[ 228 ][ 145 ],
   alphaCSR[ 228 ][ 146 ],
   alphaCSR[ 228 ][ 147 ],
   alphaCSR[ 228 ][ 148 ],
   alphaCSR[ 228 ][ 149 ],
   alphaCSR[ 228 ][ 150 ],
   alphaCSR[ 228 ][ 151 ],
   alphaCSR[ 228 ][ 152 ],
   alphaCSR[ 228 ][ 153 ],
   alphaCSR[ 228 ][ 154 ],
   alphaCSR[ 228 ][ 155 ],
   alphaCSR[ 228 ][ 156 ],
   alphaCSR[ 228 ][ 157 ],
   alphaCSR[ 228 ][ 158 ],
   alphaCSR[ 228 ][ 159 ],
   alphaCSR[ 228 ][ 160 ],
   alphaCSR[ 228 ][ 161 ],
   alphaCSR[ 228 ][ 162 ],
   alphaCSR[ 228 ][ 163 ],
   alphaCSR[ 228 ][ 164 ],
   alphaCSR[ 228 ][ 165 ],
   alphaCSR[ 228 ][ 166 ],
   alphaCSR[ 228 ][ 167 ],
   alphaCSR[ 228 ][ 168 ],
   alphaCSR[ 228 ][ 169 ],
   alphaCSR[ 228 ][ 170 ],
   alphaCSR[ 228 ][ 171 ],
   alphaCSR[ 228 ][ 172 ],
   alphaCSR[ 228 ][ 173 ],
   alphaCSR[ 228 ][ 174 ],
   alphaCSR[ 228 ][ 175 ],
   alphaCSR[ 228 ][ 176 ],
   alphaCSR[ 228 ][ 177 ],
   alphaCSR[ 228 ][ 178 ],
   alphaCSR[ 228 ][ 179 ],
   alphaCSR[ 228 ][ 180 ],
   alphaCSR[ 228 ][ 181 ],
   alphaCSR[ 228 ][ 182 ],
   alphaCSR[ 228 ][ 183 ],
   alphaCSR[ 228 ][ 184 ],
   alphaCSR[ 228 ][ 185 ],
   alphaCSR[ 228 ][ 186 ],
   alphaCSR[ 228 ][ 187 ],
   alphaCSR[ 228 ][ 188 ],
   alphaCSR[ 228 ][ 189 ],
   alphaCSR[ 228 ][ 190 ],
   alphaCSR[ 228 ][ 191 ],
   alphaCSR[ 228 ][ 192 ],
   alphaCSR[ 228 ][ 193 ],
   alphaCSR[ 228 ][ 194 ],
   alphaCSR[ 228 ][ 195 ],
   alphaCSR[ 228 ][ 196 ],
   alphaCSR[ 228 ][ 197 ],
   alphaCSR[ 228 ][ 198 ],
   alphaCSR[ 228 ][ 199 ],
   alphaCSR[ 228 ][ 200 ],
   alphaCSR[ 228 ][ 201 ],
   alphaCSR[ 228 ][ 202 ],
   alphaCSR[ 228 ][ 203 ],
   alphaCSR[ 228 ][ 204 ],
   alphaCSR[ 228 ][ 205 ],
   alphaCSR[ 228 ][ 206 ],
   alphaCSR[ 228 ][ 207 ],
   alphaCSR[ 228 ][ 208 ],
   alphaCSR[ 228 ][ 209 ],
   alphaCSR[ 228 ][ 210 ],
   alphaCSR[ 228 ][ 211 ],
   alphaCSR[ 228 ][ 212 ],
   alphaCSR[ 228 ][ 213 ],
   alphaCSR[ 228 ][ 214 ],
   alphaCSR[ 228 ][ 215 ],
   alphaCSR[ 228 ][ 216 ],
   alphaCSR[ 228 ][ 217 ],
   alphaCSR[ 228 ][ 218 ],
   alphaCSR[ 228 ][ 219 ],
   alphaCSR[ 228 ][ 220 ],
   alphaCSR[ 228 ][ 221 ],
   alphaCSR[ 228 ][ 222 ],
   alphaCSR[ 228 ][ 223 ],
   alphaCSR[ 228 ][ 224 ],
   alphaCSR[ 228 ][ 225 ],
   alphaCSR[ 228 ][ 226 ],
   alphaCSR[ 228 ][ 227 ],
   alphaCSR[ 228 ][ 228 ],
   alphaCSR[ 228 ][ 229 ],
   alphaCSR[ 228 ][ 230 ],
   alphaCSR[ 228 ][ 231 ],
   alphaCSR[ 228 ][ 232 ],
   alphaCSR[ 228 ][ 233 ],
   alphaCSR[ 228 ][ 234 ],
   alphaCSR[ 228 ][ 235 ],
   alphaCSR[ 228 ][ 236 ],
   alphaCSR[ 228 ][ 237 ],
   alphaCSR[ 228 ][ 238 ],
   alphaCSR[ 228 ][ 239 ],
   alphaCSR[ 228 ][ 240 ],
   alphaCSR[ 228 ][ 241 ],
   alphaCSR[ 228 ][ 242 ],
   alphaCSR[ 228 ][ 243 ],
   alphaCSR[ 228 ][ 244 ],
   alphaCSR[ 228 ][ 245 ],
   alphaCSR[ 228 ][ 246 ],
   alphaCSR[ 228 ][ 247 ],
   alphaCSR[ 228 ][ 248 ],
   alphaCSR[ 228 ][ 249 ],
   alphaCSR[ 228 ][ 250 ],
   alphaCSR[ 228 ][ 251 ],
   alphaCSR[ 228 ][ 252 ],
   alphaCSR[ 228 ][ 253 ],
   alphaCSR[ 228 ][ 254 ],
   alphaCSR[ 228 ][ 255 ],
   alphaCSR[ 228 ][ 256 ],
   alphaCSR[ 228 ][ 257 ],
   alphaCSR[ 228 ][ 258 ],
   alphaCSR[ 228 ][ 259 ],
   alphaCSR[ 228 ][ 260 ],
   alphaCSR[ 228 ][ 261 ],
   alphaCSR[ 228 ][ 262 ],
   alphaCSR[ 228 ][ 263 ],
   alphaCSR[ 228 ][ 264 ],
   alphaCSR[ 228 ][ 265 ],
   alphaCSR[ 228 ][ 266 ],
   alphaCSR[ 228 ][ 267 ],
   alphaCSR[ 228 ][ 268 ],
   alphaCSR[ 228 ][ 269 ],
   alphaCSR[ 228 ][ 270 ],
   alphaCSR[ 228 ][ 271 ],
   alphaCSR[ 228 ][ 272 ],
   alphaCSR[ 228 ][ 273 ],
   alphaCSR[ 228 ][ 274 ],
   alphaCSR[ 228 ][ 275 ],
   alphaCSR[ 228 ][ 276 ],
   alphaCSR[ 228 ][ 277 ],
   alphaCSR[ 228 ][ 278 ],
   alphaCSR[ 228 ][ 279 ],
   alphaCSR[ 228 ][ 280 ],
   alphaCSR[ 228 ][ 281 ],
   alphaCSR[ 228 ][ 282 ],
   alphaCSR[ 228 ][ 283 ],
   alphaCSR[ 228 ][ 284 ],
   alphaCSR[ 228 ][ 285 ],
   alphaCSR[ 228 ][ 286 ],
   alphaCSR[ 228 ][ 287 ],
   alphaCSR[ 228 ][ 288 ],
   alphaCSR[ 228 ][ 289 ],
   alphaCSR[ 228 ][ 290 ],
   alphaCSR[ 228 ][ 291 ],
   alphaCSR[ 228 ][ 292 ],
   alphaCSR[ 228 ][ 293 ],
   alphaCSR[ 228 ][ 294 ],
   alphaCSR[ 228 ][ 295 ],
   alphaCSR[ 228 ][ 296 ],
   alphaCSR[ 228 ][ 297 ],
   alphaCSR[ 228 ][ 298 ],
   alphaCSR[ 228 ][ 299 ],
   alphaCSR[ 228 ][ 300 ],
   alphaCSR[ 228 ][ 301 ],
   alphaCSR[ 228 ][ 302 ],
   alphaCSR[ 228 ][ 303 ],
   alphaCSR[ 228 ][ 304 ],
   alphaCSR[ 228 ][ 305 ],
   alphaCSR[ 228 ][ 306 ],
   alphaCSR[ 228 ][ 307 ],
   alphaCSR[ 228 ][ 308 ],
   alphaCSR[ 228 ][ 309 ],
   alphaCSR[ 228 ][ 310 ],
   alphaCSR[ 228 ][ 311 ],
   alphaCSR[ 228 ][ 312 ],
   alphaCSR[ 228 ][ 313 ],
   alphaCSR[ 228 ][ 314 ],
   alphaCSR[ 228 ][ 315 ],
   alphaCSR[ 228 ][ 316 ],
   alphaCSR[ 228 ][ 317 ],
   alphaCSR[ 228 ][ 318 ],
   alphaCSR[ 228 ][ 319 ],
   alphaCSR[ 228 ][ 320 ],
   alphaCSR[ 228 ][ 321 ],
   alphaCSR[ 228 ][ 322 ],
   alphaCSR[ 228 ][ 323 ],
   alphaCSR[ 228 ][ 324 ],
   alphaCSR[ 228 ][ 325 ],
   alphaCSR[ 228 ][ 326 ],
   alphaCSR[ 228 ][ 327 ],
   alphaCSR[ 228 ][ 328 ],
   alphaCSR[ 228 ][ 329 ],
   alphaCSR[ 228 ][ 330 ],
   alphaCSR[ 228 ][ 331 ],
   alphaCSR[ 228 ][ 332 ],
   alphaCSR[ 228 ][ 333 ],
   alphaCSR[ 228 ][ 334 ],
   alphaCSR[ 228 ][ 335 ],
   alphaCSR[ 228 ][ 336 ],
   alphaCSR[ 228 ][ 337 ],
   alphaCSR[ 228 ][ 338 ],
   alphaCSR[ 228 ][ 339 ],
   alphaCSR[ 228 ][ 340 ],
   alphaCSR[ 228 ][ 341 ],
   alphaCSR[ 228 ][ 342 ],
   alphaCSR[ 228 ][ 343 ],
   alphaCSR[ 228 ][ 344 ],
   alphaCSR[ 228 ][ 345 ],
   alphaCSR[ 228 ][ 346 ],
   alphaCSR[ 228 ][ 347 ],
   alphaCSR[ 228 ][ 348 ],
   alphaCSR[ 228 ][ 349 ],
   alphaCSR[ 228 ][ 350 ],
   alphaCSR[ 228 ][ 351 ],
   alphaCSR[ 228 ][ 352 ],
   alphaCSR[ 228 ][ 353 ],
   alphaCSR[ 228 ][ 354 ],
   alphaCSR[ 228 ][ 355 ],
   alphaCSR[ 228 ][ 356 ],
   alphaCSR[ 228 ][ 357 ],
   alphaCSR[ 228 ][ 358 ],
   alphaCSR[ 228 ][ 359 ],
   alphaCSR[ 228 ][ 360 ],
   alphaCSR[ 228 ][ 361 ],
   alphaCSR[ 228 ][ 362 ],
   alphaCSR[ 228 ][ 363 ],
   alphaCSR[ 228 ][ 364 ],
   alphaCSR[ 228 ][ 365 ],
   alphaCSR[ 228 ][ 366 ],
   alphaCSR[ 228 ][ 367 ],
   alphaCSR[ 228 ][ 368 ],
   alphaCSR[ 228 ][ 369 ],
   alphaCSR[ 228 ][ 370 ],
   alphaCSR[ 228 ][ 371 ],
   alphaCSR[ 228 ][ 372 ],
   alphaCSR[ 228 ][ 373 ],
   alphaCSR[ 228 ][ 374 ],
   alphaCSR[ 228 ][ 375 ],
   alphaCSR[ 228 ][ 376 ],
   alphaCSR[ 228 ][ 377 ],
   alphaCSR[ 228 ][ 378 ],
   alphaCSR[ 228 ][ 379 ],
   alphaCSR[ 228 ][ 380 ],
   alphaCSR[ 228 ][ 381 ],
   alphaCSR[ 228 ][ 382 ],
   alphaCSR[ 228 ][ 383 ],
   alphaCSR[ 229 ][ 0 ],
   alphaCSR[ 229 ][ 1 ],
   alphaCSR[ 229 ][ 2 ],
   alphaCSR[ 229 ][ 3 ],
   alphaCSR[ 229 ][ 4 ],
   alphaCSR[ 229 ][ 5 ],
   alphaCSR[ 229 ][ 6 ],
   alphaCSR[ 229 ][ 7 ],
   alphaCSR[ 229 ][ 8 ],
   alphaCSR[ 229 ][ 9 ],
   alphaCSR[ 229 ][ 10 ],
   alphaCSR[ 229 ][ 11 ],
   alphaCSR[ 229 ][ 12 ],
   alphaCSR[ 229 ][ 13 ],
   alphaCSR[ 229 ][ 14 ],
   alphaCSR[ 229 ][ 15 ],
   alphaCSR[ 229 ][ 16 ],
   alphaCSR[ 229 ][ 17 ],
   alphaCSR[ 229 ][ 18 ],
   alphaCSR[ 229 ][ 19 ],
   alphaCSR[ 229 ][ 20 ],
   alphaCSR[ 229 ][ 21 ],
   alphaCSR[ 229 ][ 22 ],
   alphaCSR[ 229 ][ 23 ],
   alphaCSR[ 229 ][ 24 ],
   alphaCSR[ 229 ][ 25 ],
   alphaCSR[ 229 ][ 26 ],
   alphaCSR[ 229 ][ 27 ],
   alphaCSR[ 229 ][ 28 ],
   alphaCSR[ 229 ][ 29 ],
   alphaCSR[ 229 ][ 30 ],
   alphaCSR[ 229 ][ 31 ],
   alphaCSR[ 229 ][ 32 ],
   alphaCSR[ 229 ][ 33 ],
   alphaCSR[ 229 ][ 34 ],
   alphaCSR[ 229 ][ 35 ],
   alphaCSR[ 229 ][ 36 ],
   alphaCSR[ 229 ][ 37 ],
   alphaCSR[ 229 ][ 38 ],
   alphaCSR[ 229 ][ 39 ],
   alphaCSR[ 229 ][ 40 ],
   alphaCSR[ 229 ][ 41 ],
   alphaCSR[ 229 ][ 42 ],
   alphaCSR[ 229 ][ 43 ],
   alphaCSR[ 229 ][ 44 ],
   alphaCSR[ 229 ][ 45 ],
   alphaCSR[ 229 ][ 46 ],
   alphaCSR[ 229 ][ 47 ],
   alphaCSR[ 229 ][ 48 ],
   alphaCSR[ 229 ][ 49 ],
   alphaCSR[ 229 ][ 50 ],
   alphaCSR[ 229 ][ 51 ],
   alphaCSR[ 229 ][ 52 ],
   alphaCSR[ 229 ][ 53 ],
   alphaCSR[ 229 ][ 54 ],
   alphaCSR[ 229 ][ 55 ],
   alphaCSR[ 229 ][ 56 ],
   alphaCSR[ 229 ][ 57 ],
   alphaCSR[ 229 ][ 58 ],
   alphaCSR[ 229 ][ 59 ],
   alphaCSR[ 229 ][ 60 ],
   alphaCSR[ 229 ][ 61 ],
   alphaCSR[ 229 ][ 62 ],
   alphaCSR[ 229 ][ 63 ],
   alphaCSR[ 229 ][ 64 ],
   alphaCSR[ 229 ][ 65 ],
   alphaCSR[ 229 ][ 66 ],
   alphaCSR[ 229 ][ 67 ],
   alphaCSR[ 229 ][ 68 ],
   alphaCSR[ 229 ][ 69 ],
   alphaCSR[ 229 ][ 70 ],
   alphaCSR[ 229 ][ 71 ],
   alphaCSR[ 229 ][ 72 ],
   alphaCSR[ 229 ][ 73 ],
   alphaCSR[ 229 ][ 74 ],
   alphaCSR[ 229 ][ 75 ],
   alphaCSR[ 229 ][ 76 ],
   alphaCSR[ 229 ][ 77 ],
   alphaCSR[ 229 ][ 78 ],
   alphaCSR[ 229 ][ 79 ],
   alphaCSR[ 229 ][ 80 ],
   alphaCSR[ 229 ][ 81 ],
   alphaCSR[ 229 ][ 82 ],
   alphaCSR[ 229 ][ 83 ],
   alphaCSR[ 229 ][ 84 ],
   alphaCSR[ 229 ][ 85 ],
   alphaCSR[ 229 ][ 86 ],
   alphaCSR[ 229 ][ 87 ],
   alphaCSR[ 229 ][ 88 ],
   alphaCSR[ 229 ][ 89 ],
   alphaCSR[ 229 ][ 90 ],
   alphaCSR[ 229 ][ 91 ],
   alphaCSR[ 229 ][ 92 ],
   alphaCSR[ 229 ][ 93 ],
   alphaCSR[ 229 ][ 94 ],
   alphaCSR[ 229 ][ 95 ],
   alphaCSR[ 229 ][ 96 ],
   alphaCSR[ 229 ][ 97 ],
   alphaCSR[ 229 ][ 98 ],
   alphaCSR[ 229 ][ 99 ],
   alphaCSR[ 229 ][ 100 ],
   alphaCSR[ 229 ][ 101 ],
   alphaCSR[ 229 ][ 102 ],
   alphaCSR[ 229 ][ 103 ],
   alphaCSR[ 229 ][ 104 ],
   alphaCSR[ 229 ][ 105 ],
   alphaCSR[ 229 ][ 106 ],
   alphaCSR[ 229 ][ 107 ],
   alphaCSR[ 229 ][ 108 ],
   alphaCSR[ 229 ][ 109 ],
   alphaCSR[ 229 ][ 110 ],
   alphaCSR[ 229 ][ 111 ],
   alphaCSR[ 229 ][ 112 ],
   alphaCSR[ 229 ][ 113 ],
   alphaCSR[ 229 ][ 114 ],
   alphaCSR[ 229 ][ 115 ],
   alphaCSR[ 229 ][ 116 ],
   alphaCSR[ 229 ][ 117 ],
   alphaCSR[ 229 ][ 118 ],
   alphaCSR[ 229 ][ 119 ],
   alphaCSR[ 229 ][ 120 ],
   alphaCSR[ 229 ][ 121 ],
   alphaCSR[ 229 ][ 122 ],
   alphaCSR[ 229 ][ 123 ],
   alphaCSR[ 229 ][ 124 ],
   alphaCSR[ 229 ][ 125 ],
   alphaCSR[ 229 ][ 126 ],
   alphaCSR[ 229 ][ 127 ],
   alphaCSR[ 229 ][ 128 ],
   alphaCSR[ 229 ][ 129 ],
   alphaCSR[ 229 ][ 130 ],
   alphaCSR[ 229 ][ 131 ],
   alphaCSR[ 229 ][ 132 ],
   alphaCSR[ 229 ][ 133 ],
   alphaCSR[ 229 ][ 134 ],
   alphaCSR[ 229 ][ 135 ],
   alphaCSR[ 229 ][ 136 ],
   alphaCSR[ 229 ][ 137 ],
   alphaCSR[ 229 ][ 138 ],
   alphaCSR[ 229 ][ 139 ],
   alphaCSR[ 229 ][ 140 ],
   alphaCSR[ 229 ][ 141 ],
   alphaCSR[ 229 ][ 142 ],
   alphaCSR[ 229 ][ 143 ],
   alphaCSR[ 229 ][ 144 ],
   alphaCSR[ 229 ][ 145 ],
   alphaCSR[ 229 ][ 146 ],
   alphaCSR[ 229 ][ 147 ],
   alphaCSR[ 229 ][ 148 ],
   alphaCSR[ 229 ][ 149 ],
   alphaCSR[ 229 ][ 150 ],
   alphaCSR[ 229 ][ 151 ],
   alphaCSR[ 229 ][ 152 ],
   alphaCSR[ 229 ][ 153 ],
   alphaCSR[ 229 ][ 154 ],
   alphaCSR[ 229 ][ 155 ],
   alphaCSR[ 229 ][ 156 ],
   alphaCSR[ 229 ][ 157 ],
   alphaCSR[ 229 ][ 158 ],
   alphaCSR[ 229 ][ 159 ],
   alphaCSR[ 229 ][ 160 ],
   alphaCSR[ 229 ][ 161 ],
   alphaCSR[ 229 ][ 162 ],
   alphaCSR[ 229 ][ 163 ],
   alphaCSR[ 229 ][ 164 ],
   alphaCSR[ 229 ][ 165 ],
   alphaCSR[ 229 ][ 166 ],
   alphaCSR[ 229 ][ 167 ],
   alphaCSR[ 229 ][ 168 ],
   alphaCSR[ 229 ][ 169 ],
   alphaCSR[ 229 ][ 170 ],
   alphaCSR[ 229 ][ 171 ],
   alphaCSR[ 229 ][ 172 ],
   alphaCSR[ 229 ][ 173 ],
   alphaCSR[ 229 ][ 174 ],
   alphaCSR[ 229 ][ 175 ],
   alphaCSR[ 229 ][ 176 ],
   alphaCSR[ 229 ][ 177 ],
   alphaCSR[ 229 ][ 178 ],
   alphaCSR[ 229 ][ 179 ],
   alphaCSR[ 229 ][ 180 ],
   alphaCSR[ 229 ][ 181 ],
   alphaCSR[ 229 ][ 182 ],
   alphaCSR[ 229 ][ 183 ],
   alphaCSR[ 229 ][ 184 ],
   alphaCSR[ 229 ][ 185 ],
   alphaCSR[ 229 ][ 186 ],
   alphaCSR[ 229 ][ 187 ],
   alphaCSR[ 229 ][ 188 ],
   alphaCSR[ 229 ][ 189 ],
   alphaCSR[ 229 ][ 190 ],
   alphaCSR[ 229 ][ 191 ],
   alphaCSR[ 229 ][ 192 ],
   alphaCSR[ 229 ][ 193 ],
   alphaCSR[ 229 ][ 194 ],
   alphaCSR[ 229 ][ 195 ],
   alphaCSR[ 229 ][ 196 ],
   alphaCSR[ 229 ][ 197 ],
   alphaCSR[ 229 ][ 198 ],
   alphaCSR[ 229 ][ 199 ],
   alphaCSR[ 229 ][ 200 ],
   alphaCSR[ 229 ][ 201 ],
   alphaCSR[ 229 ][ 202 ],
   alphaCSR[ 229 ][ 203 ],
   alphaCSR[ 229 ][ 204 ],
   alphaCSR[ 229 ][ 205 ],
   alphaCSR[ 229 ][ 206 ],
   alphaCSR[ 229 ][ 207 ],
   alphaCSR[ 229 ][ 208 ],
   alphaCSR[ 229 ][ 209 ],
   alphaCSR[ 229 ][ 210 ],
   alphaCSR[ 229 ][ 211 ],
   alphaCSR[ 229 ][ 212 ],
   alphaCSR[ 229 ][ 213 ],
   alphaCSR[ 229 ][ 214 ],
   alphaCSR[ 229 ][ 215 ],
   alphaCSR[ 229 ][ 216 ],
   alphaCSR[ 229 ][ 217 ],
   alphaCSR[ 229 ][ 218 ],
   alphaCSR[ 229 ][ 219 ],
   alphaCSR[ 229 ][ 220 ],
   alphaCSR[ 229 ][ 221 ],
   alphaCSR[ 229 ][ 222 ],
   alphaCSR[ 229 ][ 223 ],
   alphaCSR[ 229 ][ 224 ],
   alphaCSR[ 229 ][ 225 ],
   alphaCSR[ 229 ][ 226 ],
   alphaCSR[ 229 ][ 227 ],
   alphaCSR[ 229 ][ 228 ],
   alphaCSR[ 229 ][ 229 ],
   alphaCSR[ 229 ][ 230 ],
   alphaCSR[ 229 ][ 231 ],
   alphaCSR[ 229 ][ 232 ],
   alphaCSR[ 229 ][ 233 ],
   alphaCSR[ 229 ][ 234 ],
   alphaCSR[ 229 ][ 235 ],
   alphaCSR[ 229 ][ 236 ],
   alphaCSR[ 229 ][ 237 ],
   alphaCSR[ 229 ][ 238 ],
   alphaCSR[ 229 ][ 239 ],
   alphaCSR[ 229 ][ 240 ],
   alphaCSR[ 229 ][ 241 ],
   alphaCSR[ 229 ][ 242 ],
   alphaCSR[ 229 ][ 243 ],
   alphaCSR[ 229 ][ 244 ],
   alphaCSR[ 229 ][ 245 ],
   alphaCSR[ 229 ][ 246 ],
   alphaCSR[ 229 ][ 247 ],
   alphaCSR[ 229 ][ 248 ],
   alphaCSR[ 229 ][ 249 ],
   alphaCSR[ 229 ][ 250 ],
   alphaCSR[ 229 ][ 251 ],
   alphaCSR[ 229 ][ 252 ],
   alphaCSR[ 229 ][ 253 ],
   alphaCSR[ 229 ][ 254 ],
   alphaCSR[ 229 ][ 255 ],
   alphaCSR[ 229 ][ 256 ],
   alphaCSR[ 229 ][ 257 ],
   alphaCSR[ 229 ][ 258 ],
   alphaCSR[ 229 ][ 259 ],
   alphaCSR[ 229 ][ 260 ],
   alphaCSR[ 229 ][ 261 ],
   alphaCSR[ 229 ][ 262 ],
   alphaCSR[ 229 ][ 263 ],
   alphaCSR[ 229 ][ 264 ],
   alphaCSR[ 229 ][ 265 ],
   alphaCSR[ 229 ][ 266 ],
   alphaCSR[ 229 ][ 267 ],
   alphaCSR[ 229 ][ 268 ],
   alphaCSR[ 229 ][ 269 ],
   alphaCSR[ 229 ][ 270 ],
   alphaCSR[ 229 ][ 271 ],
   alphaCSR[ 229 ][ 272 ],
   alphaCSR[ 229 ][ 273 ],
   alphaCSR[ 229 ][ 274 ],
   alphaCSR[ 229 ][ 275 ],
   alphaCSR[ 229 ][ 276 ],
   alphaCSR[ 229 ][ 277 ],
   alphaCSR[ 229 ][ 278 ],
   alphaCSR[ 229 ][ 279 ],
   alphaCSR[ 229 ][ 280 ],
   alphaCSR[ 229 ][ 281 ],
   alphaCSR[ 229 ][ 282 ],
   alphaCSR[ 229 ][ 283 ],
   alphaCSR[ 229 ][ 284 ],
   alphaCSR[ 229 ][ 285 ],
   alphaCSR[ 229 ][ 286 ],
   alphaCSR[ 229 ][ 287 ],
   alphaCSR[ 229 ][ 288 ],
   alphaCSR[ 229 ][ 289 ],
   alphaCSR[ 229 ][ 290 ],
   alphaCSR[ 229 ][ 291 ],
   alphaCSR[ 229 ][ 292 ],
   alphaCSR[ 229 ][ 293 ],
   alphaCSR[ 229 ][ 294 ],
   alphaCSR[ 229 ][ 295 ],
   alphaCSR[ 229 ][ 296 ],
   alphaCSR[ 229 ][ 297 ],
   alphaCSR[ 229 ][ 298 ],
   alphaCSR[ 229 ][ 299 ],
   alphaCSR[ 229 ][ 300 ],
   alphaCSR[ 229 ][ 301 ],
   alphaCSR[ 229 ][ 302 ],
   alphaCSR[ 229 ][ 303 ],
   alphaCSR[ 229 ][ 304 ],
   alphaCSR[ 229 ][ 305 ],
   alphaCSR[ 229 ][ 306 ],
   alphaCSR[ 229 ][ 307 ],
   alphaCSR[ 229 ][ 308 ],
   alphaCSR[ 229 ][ 309 ],
   alphaCSR[ 229 ][ 310 ],
   alphaCSR[ 229 ][ 311 ],
   alphaCSR[ 229 ][ 312 ],
   alphaCSR[ 229 ][ 313 ],
   alphaCSR[ 229 ][ 314 ],
   alphaCSR[ 229 ][ 315 ],
   alphaCSR[ 229 ][ 316 ],
   alphaCSR[ 229 ][ 317 ],
   alphaCSR[ 229 ][ 318 ],
   alphaCSR[ 229 ][ 319 ],
   alphaCSR[ 229 ][ 320 ],
   alphaCSR[ 229 ][ 321 ],
   alphaCSR[ 229 ][ 322 ],
   alphaCSR[ 229 ][ 323 ],
   alphaCSR[ 229 ][ 324 ],
   alphaCSR[ 229 ][ 325 ],
   alphaCSR[ 229 ][ 326 ],
   alphaCSR[ 229 ][ 327 ],
   alphaCSR[ 229 ][ 328 ],
   alphaCSR[ 229 ][ 329 ],
   alphaCSR[ 229 ][ 330 ],
   alphaCSR[ 229 ][ 331 ],
   alphaCSR[ 229 ][ 332 ],
   alphaCSR[ 229 ][ 333 ],
   alphaCSR[ 229 ][ 334 ],
   alphaCSR[ 229 ][ 335 ],
   alphaCSR[ 229 ][ 336 ],
   alphaCSR[ 229 ][ 337 ],
   alphaCSR[ 229 ][ 338 ],
   alphaCSR[ 229 ][ 339 ],
   alphaCSR[ 229 ][ 340 ],
   alphaCSR[ 229 ][ 341 ],
   alphaCSR[ 229 ][ 342 ],
   alphaCSR[ 229 ][ 343 ],
   alphaCSR[ 229 ][ 344 ],
   alphaCSR[ 229 ][ 345 ],
   alphaCSR[ 229 ][ 346 ],
   alphaCSR[ 229 ][ 347 ],
   alphaCSR[ 229 ][ 348 ],
   alphaCSR[ 229 ][ 349 ],
   alphaCSR[ 229 ][ 350 ],
   alphaCSR[ 229 ][ 351 ],
   alphaCSR[ 229 ][ 352 ],
   alphaCSR[ 229 ][ 353 ],
   alphaCSR[ 229 ][ 354 ],
   alphaCSR[ 229 ][ 355 ],
   alphaCSR[ 229 ][ 356 ],
   alphaCSR[ 229 ][ 357 ],
   alphaCSR[ 229 ][ 358 ],
   alphaCSR[ 229 ][ 359 ],
   alphaCSR[ 229 ][ 360 ],
   alphaCSR[ 229 ][ 361 ],
   alphaCSR[ 229 ][ 362 ],
   alphaCSR[ 229 ][ 363 ],
   alphaCSR[ 229 ][ 364 ],
   alphaCSR[ 229 ][ 365 ],
   alphaCSR[ 229 ][ 366 ],
   alphaCSR[ 229 ][ 367 ],
   alphaCSR[ 229 ][ 368 ],
   alphaCSR[ 229 ][ 369 ],
   alphaCSR[ 229 ][ 370 ],
   alphaCSR[ 229 ][ 371 ],
   alphaCSR[ 229 ][ 372 ],
   alphaCSR[ 229 ][ 373 ],
   alphaCSR[ 229 ][ 374 ],
   alphaCSR[ 229 ][ 375 ],
   alphaCSR[ 229 ][ 376 ],
   alphaCSR[ 229 ][ 377 ],
   alphaCSR[ 229 ][ 378 ],
   alphaCSR[ 229 ][ 379 ],
   alphaCSR[ 229 ][ 380 ],
   alphaCSR[ 229 ][ 381 ],
   alphaCSR[ 229 ][ 382 ],
   alphaCSR[ 229 ][ 383 ],
   alphaCSR[ 230 ][ 0 ],
   alphaCSR[ 230 ][ 1 ],
   alphaCSR[ 230 ][ 2 ],
   alphaCSR[ 230 ][ 3 ],
   alphaCSR[ 230 ][ 4 ],
   alphaCSR[ 230 ][ 5 ],
   alphaCSR[ 230 ][ 6 ],
   alphaCSR[ 230 ][ 7 ],
   alphaCSR[ 230 ][ 8 ],
   alphaCSR[ 230 ][ 9 ],
   alphaCSR[ 230 ][ 10 ],
   alphaCSR[ 230 ][ 11 ],
   alphaCSR[ 230 ][ 12 ],
   alphaCSR[ 230 ][ 13 ],
   alphaCSR[ 230 ][ 14 ],
   alphaCSR[ 230 ][ 15 ],
   alphaCSR[ 230 ][ 16 ],
   alphaCSR[ 230 ][ 17 ],
   alphaCSR[ 230 ][ 18 ],
   alphaCSR[ 230 ][ 19 ],
   alphaCSR[ 230 ][ 20 ],
   alphaCSR[ 230 ][ 21 ],
   alphaCSR[ 230 ][ 22 ],
   alphaCSR[ 230 ][ 23 ],
   alphaCSR[ 230 ][ 24 ],
   alphaCSR[ 230 ][ 25 ],
   alphaCSR[ 230 ][ 26 ],
   alphaCSR[ 230 ][ 27 ],
   alphaCSR[ 230 ][ 28 ],
   alphaCSR[ 230 ][ 29 ],
   alphaCSR[ 230 ][ 30 ],
   alphaCSR[ 230 ][ 31 ],
   alphaCSR[ 230 ][ 32 ],
   alphaCSR[ 230 ][ 33 ],
   alphaCSR[ 230 ][ 34 ],
   alphaCSR[ 230 ][ 35 ],
   alphaCSR[ 230 ][ 36 ],
   alphaCSR[ 230 ][ 37 ],
   alphaCSR[ 230 ][ 38 ],
   alphaCSR[ 230 ][ 39 ],
   alphaCSR[ 230 ][ 40 ],
   alphaCSR[ 230 ][ 41 ],
   alphaCSR[ 230 ][ 42 ],
   alphaCSR[ 230 ][ 43 ],
   alphaCSR[ 230 ][ 44 ],
   alphaCSR[ 230 ][ 45 ],
   alphaCSR[ 230 ][ 46 ],
   alphaCSR[ 230 ][ 47 ],
   alphaCSR[ 230 ][ 48 ],
   alphaCSR[ 230 ][ 49 ],
   alphaCSR[ 230 ][ 50 ],
   alphaCSR[ 230 ][ 51 ],
   alphaCSR[ 230 ][ 52 ],
   alphaCSR[ 230 ][ 53 ],
   alphaCSR[ 230 ][ 54 ],
   alphaCSR[ 230 ][ 55 ],
   alphaCSR[ 230 ][ 56 ],
   alphaCSR[ 230 ][ 57 ],
   alphaCSR[ 230 ][ 58 ],
   alphaCSR[ 230 ][ 59 ],
   alphaCSR[ 230 ][ 60 ],
   alphaCSR[ 230 ][ 61 ],
   alphaCSR[ 230 ][ 62 ],
   alphaCSR[ 230 ][ 63 ],
   alphaCSR[ 230 ][ 64 ],
   alphaCSR[ 230 ][ 65 ],
   alphaCSR[ 230 ][ 66 ],
   alphaCSR[ 230 ][ 67 ],
   alphaCSR[ 230 ][ 68 ],
   alphaCSR[ 230 ][ 69 ],
   alphaCSR[ 230 ][ 70 ],
   alphaCSR[ 230 ][ 71 ],
   alphaCSR[ 230 ][ 72 ],
   alphaCSR[ 230 ][ 73 ],
   alphaCSR[ 230 ][ 74 ],
   alphaCSR[ 230 ][ 75 ],
   alphaCSR[ 230 ][ 76 ],
   alphaCSR[ 230 ][ 77 ],
   alphaCSR[ 230 ][ 78 ],
   alphaCSR[ 230 ][ 79 ],
   alphaCSR[ 230 ][ 80 ],
   alphaCSR[ 230 ][ 81 ],
   alphaCSR[ 230 ][ 82 ],
   alphaCSR[ 230 ][ 83 ],
   alphaCSR[ 230 ][ 84 ],
   alphaCSR[ 230 ][ 85 ],
   alphaCSR[ 230 ][ 86 ],
   alphaCSR[ 230 ][ 87 ],
   alphaCSR[ 230 ][ 88 ],
   alphaCSR[ 230 ][ 89 ],
   alphaCSR[ 230 ][ 90 ],
   alphaCSR[ 230 ][ 91 ],
   alphaCSR[ 230 ][ 92 ],
   alphaCSR[ 230 ][ 93 ],
   alphaCSR[ 230 ][ 94 ],
   alphaCSR[ 230 ][ 95 ],
   alphaCSR[ 230 ][ 96 ],
   alphaCSR[ 230 ][ 97 ],
   alphaCSR[ 230 ][ 98 ],
   alphaCSR[ 230 ][ 99 ],
   alphaCSR[ 230 ][ 100 ],
   alphaCSR[ 230 ][ 101 ],
   alphaCSR[ 230 ][ 102 ],
   alphaCSR[ 230 ][ 103 ],
   alphaCSR[ 230 ][ 104 ],
   alphaCSR[ 230 ][ 105 ],
   alphaCSR[ 230 ][ 106 ],
   alphaCSR[ 230 ][ 107 ],
   alphaCSR[ 230 ][ 108 ],
   alphaCSR[ 230 ][ 109 ],
   alphaCSR[ 230 ][ 110 ],
   alphaCSR[ 230 ][ 111 ],
   alphaCSR[ 230 ][ 112 ],
   alphaCSR[ 230 ][ 113 ],
   alphaCSR[ 230 ][ 114 ],
   alphaCSR[ 230 ][ 115 ],
   alphaCSR[ 230 ][ 116 ],
   alphaCSR[ 230 ][ 117 ],
   alphaCSR[ 230 ][ 118 ],
   alphaCSR[ 230 ][ 119 ],
   alphaCSR[ 230 ][ 120 ],
   alphaCSR[ 230 ][ 121 ],
   alphaCSR[ 230 ][ 122 ],
   alphaCSR[ 230 ][ 123 ],
   alphaCSR[ 230 ][ 124 ],
   alphaCSR[ 230 ][ 125 ],
   alphaCSR[ 230 ][ 126 ],
   alphaCSR[ 230 ][ 127 ],
   alphaCSR[ 230 ][ 128 ],
   alphaCSR[ 230 ][ 129 ],
   alphaCSR[ 230 ][ 130 ],
   alphaCSR[ 230 ][ 131 ],
   alphaCSR[ 230 ][ 132 ],
   alphaCSR[ 230 ][ 133 ],
   alphaCSR[ 230 ][ 134 ],
   alphaCSR[ 230 ][ 135 ],
   alphaCSR[ 230 ][ 136 ],
   alphaCSR[ 230 ][ 137 ],
   alphaCSR[ 230 ][ 138 ],
   alphaCSR[ 230 ][ 139 ],
   alphaCSR[ 230 ][ 140 ],
   alphaCSR[ 230 ][ 141 ],
   alphaCSR[ 230 ][ 142 ],
   alphaCSR[ 230 ][ 143 ],
   alphaCSR[ 230 ][ 144 ],
   alphaCSR[ 230 ][ 145 ],
   alphaCSR[ 230 ][ 146 ],
   alphaCSR[ 230 ][ 147 ],
   alphaCSR[ 230 ][ 148 ],
   alphaCSR[ 230 ][ 149 ],
   alphaCSR[ 230 ][ 150 ],
   alphaCSR[ 230 ][ 151 ],
   alphaCSR[ 230 ][ 152 ],
   alphaCSR[ 230 ][ 153 ],
   alphaCSR[ 230 ][ 154 ],
   alphaCSR[ 230 ][ 155 ],
   alphaCSR[ 230 ][ 156 ],
   alphaCSR[ 230 ][ 157 ],
   alphaCSR[ 230 ][ 158 ],
   alphaCSR[ 230 ][ 159 ],
   alphaCSR[ 230 ][ 160 ],
   alphaCSR[ 230 ][ 161 ],
   alphaCSR[ 230 ][ 162 ],
   alphaCSR[ 230 ][ 163 ],
   alphaCSR[ 230 ][ 164 ],
   alphaCSR[ 230 ][ 165 ],
   alphaCSR[ 230 ][ 166 ],
   alphaCSR[ 230 ][ 167 ],
   alphaCSR[ 230 ][ 168 ],
   alphaCSR[ 230 ][ 169 ],
   alphaCSR[ 230 ][ 170 ],
   alphaCSR[ 230 ][ 171 ],
   alphaCSR[ 230 ][ 172 ],
   alphaCSR[ 230 ][ 173 ],
   alphaCSR[ 230 ][ 174 ],
   alphaCSR[ 230 ][ 175 ],
   alphaCSR[ 230 ][ 176 ],
   alphaCSR[ 230 ][ 177 ],
   alphaCSR[ 230 ][ 178 ],
   alphaCSR[ 230 ][ 179 ],
   alphaCSR[ 230 ][ 180 ],
   alphaCSR[ 230 ][ 181 ],
   alphaCSR[ 230 ][ 182 ],
   alphaCSR[ 230 ][ 183 ],
   alphaCSR[ 230 ][ 184 ],
   alphaCSR[ 230 ][ 185 ],
   alphaCSR[ 230 ][ 186 ],
   alphaCSR[ 230 ][ 187 ],
   alphaCSR[ 230 ][ 188 ],
   alphaCSR[ 230 ][ 189 ],
   alphaCSR[ 230 ][ 190 ],
   alphaCSR[ 230 ][ 191 ],
   alphaCSR[ 230 ][ 192 ],
   alphaCSR[ 230 ][ 193 ],
   alphaCSR[ 230 ][ 194 ],
   alphaCSR[ 230 ][ 195 ],
   alphaCSR[ 230 ][ 196 ],
   alphaCSR[ 230 ][ 197 ],
   alphaCSR[ 230 ][ 198 ],
   alphaCSR[ 230 ][ 199 ],
   alphaCSR[ 230 ][ 200 ],
   alphaCSR[ 230 ][ 201 ],
   alphaCSR[ 230 ][ 202 ],
   alphaCSR[ 230 ][ 203 ],
   alphaCSR[ 230 ][ 204 ],
   alphaCSR[ 230 ][ 205 ],
   alphaCSR[ 230 ][ 206 ],
   alphaCSR[ 230 ][ 207 ],
   alphaCSR[ 230 ][ 208 ],
   alphaCSR[ 230 ][ 209 ],
   alphaCSR[ 230 ][ 210 ],
   alphaCSR[ 230 ][ 211 ],
   alphaCSR[ 230 ][ 212 ],
   alphaCSR[ 230 ][ 213 ],
   alphaCSR[ 230 ][ 214 ],
   alphaCSR[ 230 ][ 215 ],
   alphaCSR[ 230 ][ 216 ],
   alphaCSR[ 230 ][ 217 ],
   alphaCSR[ 230 ][ 218 ],
   alphaCSR[ 230 ][ 219 ],
   alphaCSR[ 230 ][ 220 ],
   alphaCSR[ 230 ][ 221 ],
   alphaCSR[ 230 ][ 222 ],
   alphaCSR[ 230 ][ 223 ],
   alphaCSR[ 230 ][ 224 ],
   alphaCSR[ 230 ][ 225 ],
   alphaCSR[ 230 ][ 226 ],
   alphaCSR[ 230 ][ 227 ],
   alphaCSR[ 230 ][ 228 ],
   alphaCSR[ 230 ][ 229 ],
   alphaCSR[ 230 ][ 230 ],
   alphaCSR[ 230 ][ 231 ],
   alphaCSR[ 230 ][ 232 ],
   alphaCSR[ 230 ][ 233 ],
   alphaCSR[ 230 ][ 234 ],
   alphaCSR[ 230 ][ 235 ],
   alphaCSR[ 230 ][ 236 ],
   alphaCSR[ 230 ][ 237 ],
   alphaCSR[ 230 ][ 238 ],
   alphaCSR[ 230 ][ 239 ],
   alphaCSR[ 230 ][ 240 ],
   alphaCSR[ 230 ][ 241 ],
   alphaCSR[ 230 ][ 242 ],
   alphaCSR[ 230 ][ 243 ],
   alphaCSR[ 230 ][ 244 ],
   alphaCSR[ 230 ][ 245 ],
   alphaCSR[ 230 ][ 246 ],
   alphaCSR[ 230 ][ 247 ],
   alphaCSR[ 230 ][ 248 ],
   alphaCSR[ 230 ][ 249 ],
   alphaCSR[ 230 ][ 250 ],
   alphaCSR[ 230 ][ 251 ],
   alphaCSR[ 230 ][ 252 ],
   alphaCSR[ 230 ][ 253 ],
   alphaCSR[ 230 ][ 254 ],
   alphaCSR[ 230 ][ 255 ],
   alphaCSR[ 230 ][ 256 ],
   alphaCSR[ 230 ][ 257 ],
   alphaCSR[ 230 ][ 258 ],
   alphaCSR[ 230 ][ 259 ],
   alphaCSR[ 230 ][ 260 ],
   alphaCSR[ 230 ][ 261 ],
   alphaCSR[ 230 ][ 262 ],
   alphaCSR[ 230 ][ 263 ],
   alphaCSR[ 230 ][ 264 ],
   alphaCSR[ 230 ][ 265 ],
   alphaCSR[ 230 ][ 266 ],
   alphaCSR[ 230 ][ 267 ],
   alphaCSR[ 230 ][ 268 ],
   alphaCSR[ 230 ][ 269 ],
   alphaCSR[ 230 ][ 270 ],
   alphaCSR[ 230 ][ 271 ],
   alphaCSR[ 230 ][ 272 ],
   alphaCSR[ 230 ][ 273 ],
   alphaCSR[ 230 ][ 274 ],
   alphaCSR[ 230 ][ 275 ],
   alphaCSR[ 230 ][ 276 ],
   alphaCSR[ 230 ][ 277 ],
   alphaCSR[ 230 ][ 278 ],
   alphaCSR[ 230 ][ 279 ],
   alphaCSR[ 230 ][ 280 ],
   alphaCSR[ 230 ][ 281 ],
   alphaCSR[ 230 ][ 282 ],
   alphaCSR[ 230 ][ 283 ],
   alphaCSR[ 230 ][ 284 ],
   alphaCSR[ 230 ][ 285 ],
   alphaCSR[ 230 ][ 286 ],
   alphaCSR[ 230 ][ 287 ],
   alphaCSR[ 230 ][ 288 ],
   alphaCSR[ 230 ][ 289 ],
   alphaCSR[ 230 ][ 290 ],
   alphaCSR[ 230 ][ 291 ],
   alphaCSR[ 230 ][ 292 ],
   alphaCSR[ 230 ][ 293 ],
   alphaCSR[ 230 ][ 294 ],
   alphaCSR[ 230 ][ 295 ],
   alphaCSR[ 230 ][ 296 ],
   alphaCSR[ 230 ][ 297 ],
   alphaCSR[ 230 ][ 298 ],
   alphaCSR[ 230 ][ 299 ],
   alphaCSR[ 230 ][ 300 ],
   alphaCSR[ 230 ][ 301 ],
   alphaCSR[ 230 ][ 302 ],
   alphaCSR[ 230 ][ 303 ],
   alphaCSR[ 230 ][ 304 ],
   alphaCSR[ 230 ][ 305 ],
   alphaCSR[ 230 ][ 306 ],
   alphaCSR[ 230 ][ 307 ],
   alphaCSR[ 230 ][ 308 ],
   alphaCSR[ 230 ][ 309 ],
   alphaCSR[ 230 ][ 310 ],
   alphaCSR[ 230 ][ 311 ],
   alphaCSR[ 230 ][ 312 ],
   alphaCSR[ 230 ][ 313 ],
   alphaCSR[ 230 ][ 314 ],
   alphaCSR[ 230 ][ 315 ],
   alphaCSR[ 230 ][ 316 ],
   alphaCSR[ 230 ][ 317 ],
   alphaCSR[ 230 ][ 318 ],
   alphaCSR[ 230 ][ 319 ],
   alphaCSR[ 230 ][ 320 ],
   alphaCSR[ 230 ][ 321 ],
   alphaCSR[ 230 ][ 322 ],
   alphaCSR[ 230 ][ 323 ],
   alphaCSR[ 230 ][ 324 ],
   alphaCSR[ 230 ][ 325 ],
   alphaCSR[ 230 ][ 326 ],
   alphaCSR[ 230 ][ 327 ],
   alphaCSR[ 230 ][ 328 ],
   alphaCSR[ 230 ][ 329 ],
   alphaCSR[ 230 ][ 330 ],
   alphaCSR[ 230 ][ 331 ],
   alphaCSR[ 230 ][ 332 ],
   alphaCSR[ 230 ][ 333 ],
   alphaCSR[ 230 ][ 334 ],
   alphaCSR[ 230 ][ 335 ],
   alphaCSR[ 230 ][ 336 ],
   alphaCSR[ 230 ][ 337 ],
   alphaCSR[ 230 ][ 338 ],
   alphaCSR[ 230 ][ 339 ],
   alphaCSR[ 230 ][ 340 ],
   alphaCSR[ 230 ][ 341 ],
   alphaCSR[ 230 ][ 342 ],
   alphaCSR[ 230 ][ 343 ],
   alphaCSR[ 230 ][ 344 ],
   alphaCSR[ 230 ][ 345 ],
   alphaCSR[ 230 ][ 346 ],
   alphaCSR[ 230 ][ 347 ],
   alphaCSR[ 230 ][ 348 ],
   alphaCSR[ 230 ][ 349 ],
   alphaCSR[ 230 ][ 350 ],
   alphaCSR[ 230 ][ 351 ],
   alphaCSR[ 230 ][ 352 ],
   alphaCSR[ 230 ][ 353 ],
   alphaCSR[ 230 ][ 354 ],
   alphaCSR[ 230 ][ 355 ],
   alphaCSR[ 230 ][ 356 ],
   alphaCSR[ 230 ][ 357 ],
   alphaCSR[ 230 ][ 358 ],
   alphaCSR[ 230 ][ 359 ],
   alphaCSR[ 230 ][ 360 ],
   alphaCSR[ 230 ][ 361 ],
   alphaCSR[ 230 ][ 362 ],
   alphaCSR[ 230 ][ 363 ],
   alphaCSR[ 230 ][ 364 ],
   alphaCSR[ 230 ][ 365 ],
   alphaCSR[ 230 ][ 366 ],
   alphaCSR[ 230 ][ 367 ],
   alphaCSR[ 230 ][ 368 ],
   alphaCSR[ 230 ][ 369 ],
   alphaCSR[ 230 ][ 370 ],
   alphaCSR[ 230 ][ 371 ],
   alphaCSR[ 230 ][ 372 ],
   alphaCSR[ 230 ][ 373 ],
   alphaCSR[ 230 ][ 374 ],
   alphaCSR[ 230 ][ 375 ],
   alphaCSR[ 230 ][ 376 ],
   alphaCSR[ 230 ][ 377 ],
   alphaCSR[ 230 ][ 378 ],
   alphaCSR[ 230 ][ 379 ],
   alphaCSR[ 230 ][ 380 ],
   alphaCSR[ 230 ][ 381 ],
   alphaCSR[ 230 ][ 382 ],
   alphaCSR[ 230 ][ 383 ],
   alphaCSR[ 231 ][ 0 ],
   alphaCSR[ 231 ][ 1 ],
   alphaCSR[ 231 ][ 2 ],
   alphaCSR[ 231 ][ 3 ],
   alphaCSR[ 231 ][ 4 ],
   alphaCSR[ 231 ][ 5 ],
   alphaCSR[ 231 ][ 6 ],
   alphaCSR[ 231 ][ 7 ],
   alphaCSR[ 231 ][ 8 ],
   alphaCSR[ 231 ][ 9 ],
   alphaCSR[ 231 ][ 10 ],
   alphaCSR[ 231 ][ 11 ],
   alphaCSR[ 231 ][ 12 ],
   alphaCSR[ 231 ][ 13 ],
   alphaCSR[ 231 ][ 14 ],
   alphaCSR[ 231 ][ 15 ],
   alphaCSR[ 231 ][ 16 ],
   alphaCSR[ 231 ][ 17 ],
   alphaCSR[ 231 ][ 18 ],
   alphaCSR[ 231 ][ 19 ],
   alphaCSR[ 231 ][ 20 ],
   alphaCSR[ 231 ][ 21 ],
   alphaCSR[ 231 ][ 22 ],
   alphaCSR[ 231 ][ 23 ],
   alphaCSR[ 231 ][ 24 ],
   alphaCSR[ 231 ][ 25 ],
   alphaCSR[ 231 ][ 26 ],
   alphaCSR[ 231 ][ 27 ],
   alphaCSR[ 231 ][ 28 ],
   alphaCSR[ 231 ][ 29 ],
   alphaCSR[ 231 ][ 30 ],
   alphaCSR[ 231 ][ 31 ],
   alphaCSR[ 231 ][ 32 ],
   alphaCSR[ 231 ][ 33 ],
   alphaCSR[ 231 ][ 34 ],
   alphaCSR[ 231 ][ 35 ],
   alphaCSR[ 231 ][ 36 ],
   alphaCSR[ 231 ][ 37 ],
   alphaCSR[ 231 ][ 38 ],
   alphaCSR[ 231 ][ 39 ],
   alphaCSR[ 231 ][ 40 ],
   alphaCSR[ 231 ][ 41 ],
   alphaCSR[ 231 ][ 42 ],
   alphaCSR[ 231 ][ 43 ],
   alphaCSR[ 231 ][ 44 ],
   alphaCSR[ 231 ][ 45 ],
   alphaCSR[ 231 ][ 46 ],
   alphaCSR[ 231 ][ 47 ],
   alphaCSR[ 231 ][ 48 ],
   alphaCSR[ 231 ][ 49 ],
   alphaCSR[ 231 ][ 50 ],
   alphaCSR[ 231 ][ 51 ],
   alphaCSR[ 231 ][ 52 ],
   alphaCSR[ 231 ][ 53 ],
   alphaCSR[ 231 ][ 54 ],
   alphaCSR[ 231 ][ 55 ],
   alphaCSR[ 231 ][ 56 ],
   alphaCSR[ 231 ][ 57 ],
   alphaCSR[ 231 ][ 58 ],
   alphaCSR[ 231 ][ 59 ],
   alphaCSR[ 231 ][ 60 ],
   alphaCSR[ 231 ][ 61 ],
   alphaCSR[ 231 ][ 62 ],
   alphaCSR[ 231 ][ 63 ],
   alphaCSR[ 231 ][ 64 ],
   alphaCSR[ 231 ][ 65 ],
   alphaCSR[ 231 ][ 66 ],
   alphaCSR[ 231 ][ 67 ],
   alphaCSR[ 231 ][ 68 ],
   alphaCSR[ 231 ][ 69 ],
   alphaCSR[ 231 ][ 70 ],
   alphaCSR[ 231 ][ 71 ],
   alphaCSR[ 231 ][ 72 ],
   alphaCSR[ 231 ][ 73 ],
   alphaCSR[ 231 ][ 74 ],
   alphaCSR[ 231 ][ 75 ],
   alphaCSR[ 231 ][ 76 ],
   alphaCSR[ 231 ][ 77 ],
   alphaCSR[ 231 ][ 78 ],
   alphaCSR[ 231 ][ 79 ],
   alphaCSR[ 231 ][ 80 ],
   alphaCSR[ 231 ][ 81 ],
   alphaCSR[ 231 ][ 82 ],
   alphaCSR[ 231 ][ 83 ],
   alphaCSR[ 231 ][ 84 ],
   alphaCSR[ 231 ][ 85 ],
   alphaCSR[ 231 ][ 86 ],
   alphaCSR[ 231 ][ 87 ],
   alphaCSR[ 231 ][ 88 ],
   alphaCSR[ 231 ][ 89 ],
   alphaCSR[ 231 ][ 90 ],
   alphaCSR[ 231 ][ 91 ],
   alphaCSR[ 231 ][ 92 ],
   alphaCSR[ 231 ][ 93 ],
   alphaCSR[ 231 ][ 94 ],
   alphaCSR[ 231 ][ 95 ],
   alphaCSR[ 231 ][ 96 ],
   alphaCSR[ 231 ][ 97 ],
   alphaCSR[ 231 ][ 98 ],
   alphaCSR[ 231 ][ 99 ],
   alphaCSR[ 231 ][ 100 ],
   alphaCSR[ 231 ][ 101 ],
   alphaCSR[ 231 ][ 102 ],
   alphaCSR[ 231 ][ 103 ],
   alphaCSR[ 231 ][ 104 ],
   alphaCSR[ 231 ][ 105 ],
   alphaCSR[ 231 ][ 106 ],
   alphaCSR[ 231 ][ 107 ],
   alphaCSR[ 231 ][ 108 ],
   alphaCSR[ 231 ][ 109 ],
   alphaCSR[ 231 ][ 110 ],
   alphaCSR[ 231 ][ 111 ],
   alphaCSR[ 231 ][ 112 ],
   alphaCSR[ 231 ][ 113 ],
   alphaCSR[ 231 ][ 114 ],
   alphaCSR[ 231 ][ 115 ],
   alphaCSR[ 231 ][ 116 ],
   alphaCSR[ 231 ][ 117 ],
   alphaCSR[ 231 ][ 118 ],
   alphaCSR[ 231 ][ 119 ],
   alphaCSR[ 231 ][ 120 ],
   alphaCSR[ 231 ][ 121 ],
   alphaCSR[ 231 ][ 122 ],
   alphaCSR[ 231 ][ 123 ],
   alphaCSR[ 231 ][ 124 ],
   alphaCSR[ 231 ][ 125 ],
   alphaCSR[ 231 ][ 126 ],
   alphaCSR[ 231 ][ 127 ],
   alphaCSR[ 231 ][ 128 ],
   alphaCSR[ 231 ][ 129 ],
   alphaCSR[ 231 ][ 130 ],
   alphaCSR[ 231 ][ 131 ],
   alphaCSR[ 231 ][ 132 ],
   alphaCSR[ 231 ][ 133 ],
   alphaCSR[ 231 ][ 134 ],
   alphaCSR[ 231 ][ 135 ],
   alphaCSR[ 231 ][ 136 ],
   alphaCSR[ 231 ][ 137 ],
   alphaCSR[ 231 ][ 138 ],
   alphaCSR[ 231 ][ 139 ],
   alphaCSR[ 231 ][ 140 ],
   alphaCSR[ 231 ][ 141 ],
   alphaCSR[ 231 ][ 142 ],
   alphaCSR[ 231 ][ 143 ],
   alphaCSR[ 231 ][ 144 ],
   alphaCSR[ 231 ][ 145 ],
   alphaCSR[ 231 ][ 146 ],
   alphaCSR[ 231 ][ 147 ],
   alphaCSR[ 231 ][ 148 ],
   alphaCSR[ 231 ][ 149 ],
   alphaCSR[ 231 ][ 150 ],
   alphaCSR[ 231 ][ 151 ],
   alphaCSR[ 231 ][ 152 ],
   alphaCSR[ 231 ][ 153 ],
   alphaCSR[ 231 ][ 154 ],
   alphaCSR[ 231 ][ 155 ],
   alphaCSR[ 231 ][ 156 ],
   alphaCSR[ 231 ][ 157 ],
   alphaCSR[ 231 ][ 158 ],
   alphaCSR[ 231 ][ 159 ],
   alphaCSR[ 231 ][ 160 ],
   alphaCSR[ 231 ][ 161 ],
   alphaCSR[ 231 ][ 162 ],
   alphaCSR[ 231 ][ 163 ],
   alphaCSR[ 231 ][ 164 ],
   alphaCSR[ 231 ][ 165 ],
   alphaCSR[ 231 ][ 166 ],
   alphaCSR[ 231 ][ 167 ],
   alphaCSR[ 231 ][ 168 ],
   alphaCSR[ 231 ][ 169 ],
   alphaCSR[ 231 ][ 170 ],
   alphaCSR[ 231 ][ 171 ],
   alphaCSR[ 231 ][ 172 ],
   alphaCSR[ 231 ][ 173 ],
   alphaCSR[ 231 ][ 174 ],
   alphaCSR[ 231 ][ 175 ],
   alphaCSR[ 231 ][ 176 ],
   alphaCSR[ 231 ][ 177 ],
   alphaCSR[ 231 ][ 178 ],
   alphaCSR[ 231 ][ 179 ],
   alphaCSR[ 231 ][ 180 ],
   alphaCSR[ 231 ][ 181 ],
   alphaCSR[ 231 ][ 182 ],
   alphaCSR[ 231 ][ 183 ],
   alphaCSR[ 231 ][ 184 ],
   alphaCSR[ 231 ][ 185 ],
   alphaCSR[ 231 ][ 186 ],
   alphaCSR[ 231 ][ 187 ],
   alphaCSR[ 231 ][ 188 ],
   alphaCSR[ 231 ][ 189 ],
   alphaCSR[ 231 ][ 190 ],
   alphaCSR[ 231 ][ 191 ],
   alphaCSR[ 231 ][ 192 ],
   alphaCSR[ 231 ][ 193 ],
   alphaCSR[ 231 ][ 194 ],
   alphaCSR[ 231 ][ 195 ],
   alphaCSR[ 231 ][ 196 ],
   alphaCSR[ 231 ][ 197 ],
   alphaCSR[ 231 ][ 198 ],
   alphaCSR[ 231 ][ 199 ],
   alphaCSR[ 231 ][ 200 ],
   alphaCSR[ 231 ][ 201 ],
   alphaCSR[ 231 ][ 202 ],
   alphaCSR[ 231 ][ 203 ],
   alphaCSR[ 231 ][ 204 ],
   alphaCSR[ 231 ][ 205 ],
   alphaCSR[ 231 ][ 206 ],
   alphaCSR[ 231 ][ 207 ],
   alphaCSR[ 231 ][ 208 ],
   alphaCSR[ 231 ][ 209 ],
   alphaCSR[ 231 ][ 210 ],
   alphaCSR[ 231 ][ 211 ],
   alphaCSR[ 231 ][ 212 ],
   alphaCSR[ 231 ][ 213 ],
   alphaCSR[ 231 ][ 214 ],
   alphaCSR[ 231 ][ 215 ],
   alphaCSR[ 231 ][ 216 ],
   alphaCSR[ 231 ][ 217 ],
   alphaCSR[ 231 ][ 218 ],
   alphaCSR[ 231 ][ 219 ],
   alphaCSR[ 231 ][ 220 ],
   alphaCSR[ 231 ][ 221 ],
   alphaCSR[ 231 ][ 222 ],
   alphaCSR[ 231 ][ 223 ],
   alphaCSR[ 231 ][ 224 ],
   alphaCSR[ 231 ][ 225 ],
   alphaCSR[ 231 ][ 226 ],
   alphaCSR[ 231 ][ 227 ],
   alphaCSR[ 231 ][ 228 ],
   alphaCSR[ 231 ][ 229 ],
   alphaCSR[ 231 ][ 230 ],
   alphaCSR[ 231 ][ 231 ],
   alphaCSR[ 231 ][ 232 ],
   alphaCSR[ 231 ][ 233 ],
   alphaCSR[ 231 ][ 234 ],
   alphaCSR[ 231 ][ 235 ],
   alphaCSR[ 231 ][ 236 ],
   alphaCSR[ 231 ][ 237 ],
   alphaCSR[ 231 ][ 238 ],
   alphaCSR[ 231 ][ 239 ],
   alphaCSR[ 231 ][ 240 ],
   alphaCSR[ 231 ][ 241 ],
   alphaCSR[ 231 ][ 242 ],
   alphaCSR[ 231 ][ 243 ],
   alphaCSR[ 231 ][ 244 ],
   alphaCSR[ 231 ][ 245 ],
   alphaCSR[ 231 ][ 246 ],
   alphaCSR[ 231 ][ 247 ],
   alphaCSR[ 231 ][ 248 ],
   alphaCSR[ 231 ][ 249 ],
   alphaCSR[ 231 ][ 250 ],
   alphaCSR[ 231 ][ 251 ],
   alphaCSR[ 231 ][ 252 ],
   alphaCSR[ 231 ][ 253 ],
   alphaCSR[ 231 ][ 254 ],
   alphaCSR[ 231 ][ 255 ],
   alphaCSR[ 231 ][ 256 ],
   alphaCSR[ 231 ][ 257 ],
   alphaCSR[ 231 ][ 258 ],
   alphaCSR[ 231 ][ 259 ],
   alphaCSR[ 231 ][ 260 ],
   alphaCSR[ 231 ][ 261 ],
   alphaCSR[ 231 ][ 262 ],
   alphaCSR[ 231 ][ 263 ],
   alphaCSR[ 231 ][ 264 ],
   alphaCSR[ 231 ][ 265 ],
   alphaCSR[ 231 ][ 266 ],
   alphaCSR[ 231 ][ 267 ],
   alphaCSR[ 231 ][ 268 ],
   alphaCSR[ 231 ][ 269 ],
   alphaCSR[ 231 ][ 270 ],
   alphaCSR[ 231 ][ 271 ],
   alphaCSR[ 231 ][ 272 ],
   alphaCSR[ 231 ][ 273 ],
   alphaCSR[ 231 ][ 274 ],
   alphaCSR[ 231 ][ 275 ],
   alphaCSR[ 231 ][ 276 ],
   alphaCSR[ 231 ][ 277 ],
   alphaCSR[ 231 ][ 278 ],
   alphaCSR[ 231 ][ 279 ],
   alphaCSR[ 231 ][ 280 ],
   alphaCSR[ 231 ][ 281 ],
   alphaCSR[ 231 ][ 282 ],
   alphaCSR[ 231 ][ 283 ],
   alphaCSR[ 231 ][ 284 ],
   alphaCSR[ 231 ][ 285 ],
   alphaCSR[ 231 ][ 286 ],
   alphaCSR[ 231 ][ 287 ],
   alphaCSR[ 231 ][ 288 ],
   alphaCSR[ 231 ][ 289 ],
   alphaCSR[ 231 ][ 290 ],
   alphaCSR[ 231 ][ 291 ],
   alphaCSR[ 231 ][ 292 ],
   alphaCSR[ 231 ][ 293 ],
   alphaCSR[ 231 ][ 294 ],
   alphaCSR[ 231 ][ 295 ],
   alphaCSR[ 231 ][ 296 ],
   alphaCSR[ 231 ][ 297 ],
   alphaCSR[ 231 ][ 298 ],
   alphaCSR[ 231 ][ 299 ],
   alphaCSR[ 231 ][ 300 ],
   alphaCSR[ 231 ][ 301 ],
   alphaCSR[ 231 ][ 302 ],
   alphaCSR[ 231 ][ 303 ],
   alphaCSR[ 231 ][ 304 ],
   alphaCSR[ 231 ][ 305 ],
   alphaCSR[ 231 ][ 306 ],
   alphaCSR[ 231 ][ 307 ],
   alphaCSR[ 231 ][ 308 ],
   alphaCSR[ 231 ][ 309 ],
   alphaCSR[ 231 ][ 310 ],
   alphaCSR[ 231 ][ 311 ],
   alphaCSR[ 231 ][ 312 ],
   alphaCSR[ 231 ][ 313 ],
   alphaCSR[ 231 ][ 314 ],
   alphaCSR[ 231 ][ 315 ],
   alphaCSR[ 231 ][ 316 ],
   alphaCSR[ 231 ][ 317 ],
   alphaCSR[ 231 ][ 318 ],
   alphaCSR[ 231 ][ 319 ],
   alphaCSR[ 231 ][ 320 ],
   alphaCSR[ 231 ][ 321 ],
   alphaCSR[ 231 ][ 322 ],
   alphaCSR[ 231 ][ 323 ],
   alphaCSR[ 231 ][ 324 ],
   alphaCSR[ 231 ][ 325 ],
   alphaCSR[ 231 ][ 326 ],
   alphaCSR[ 231 ][ 327 ],
   alphaCSR[ 231 ][ 328 ],
   alphaCSR[ 231 ][ 329 ],
   alphaCSR[ 231 ][ 330 ],
   alphaCSR[ 231 ][ 331 ],
   alphaCSR[ 231 ][ 332 ],
   alphaCSR[ 231 ][ 333 ],
   alphaCSR[ 231 ][ 334 ],
   alphaCSR[ 231 ][ 335 ],
   alphaCSR[ 231 ][ 336 ],
   alphaCSR[ 231 ][ 337 ],
   alphaCSR[ 231 ][ 338 ],
   alphaCSR[ 231 ][ 339 ],
   alphaCSR[ 231 ][ 340 ],
   alphaCSR[ 231 ][ 341 ],
   alphaCSR[ 231 ][ 342 ],
   alphaCSR[ 231 ][ 343 ],
   alphaCSR[ 231 ][ 344 ],
   alphaCSR[ 231 ][ 345 ],
   alphaCSR[ 231 ][ 346 ],
   alphaCSR[ 231 ][ 347 ],
   alphaCSR[ 231 ][ 348 ],
   alphaCSR[ 231 ][ 349 ],
   alphaCSR[ 231 ][ 350 ],
   alphaCSR[ 231 ][ 351 ],
   alphaCSR[ 231 ][ 352 ],
   alphaCSR[ 231 ][ 353 ],
   alphaCSR[ 231 ][ 354 ],
   alphaCSR[ 231 ][ 355 ],
   alphaCSR[ 231 ][ 356 ],
   alphaCSR[ 231 ][ 357 ],
   alphaCSR[ 231 ][ 358 ],
   alphaCSR[ 231 ][ 359 ],
   alphaCSR[ 231 ][ 360 ],
   alphaCSR[ 231 ][ 361 ],
   alphaCSR[ 231 ][ 362 ],
   alphaCSR[ 231 ][ 363 ],
   alphaCSR[ 231 ][ 364 ],
   alphaCSR[ 231 ][ 365 ],
   alphaCSR[ 231 ][ 366 ],
   alphaCSR[ 231 ][ 367 ],
   alphaCSR[ 231 ][ 368 ],
   alphaCSR[ 231 ][ 369 ],
   alphaCSR[ 231 ][ 370 ],
   alphaCSR[ 231 ][ 371 ],
   alphaCSR[ 231 ][ 372 ],
   alphaCSR[ 231 ][ 373 ],
   alphaCSR[ 231 ][ 374 ],
   alphaCSR[ 231 ][ 375 ],
   alphaCSR[ 231 ][ 376 ],
   alphaCSR[ 231 ][ 377 ],
   alphaCSR[ 231 ][ 378 ],
   alphaCSR[ 231 ][ 379 ],
   alphaCSR[ 231 ][ 380 ],
   alphaCSR[ 231 ][ 381 ],
   alphaCSR[ 231 ][ 382 ],
   alphaCSR[ 231 ][ 383 ],
   alphaCSR[ 232 ][ 0 ],
   alphaCSR[ 232 ][ 1 ],
   alphaCSR[ 232 ][ 2 ],
   alphaCSR[ 232 ][ 3 ],
   alphaCSR[ 232 ][ 4 ],
   alphaCSR[ 232 ][ 5 ],
   alphaCSR[ 232 ][ 6 ],
   alphaCSR[ 232 ][ 7 ],
   alphaCSR[ 232 ][ 8 ],
   alphaCSR[ 232 ][ 9 ],
   alphaCSR[ 232 ][ 10 ],
   alphaCSR[ 232 ][ 11 ],
   alphaCSR[ 232 ][ 12 ],
   alphaCSR[ 232 ][ 13 ],
   alphaCSR[ 232 ][ 14 ],
   alphaCSR[ 232 ][ 15 ],
   alphaCSR[ 232 ][ 16 ],
   alphaCSR[ 232 ][ 17 ],
   alphaCSR[ 232 ][ 18 ],
   alphaCSR[ 232 ][ 19 ],
   alphaCSR[ 232 ][ 20 ],
   alphaCSR[ 232 ][ 21 ],
   alphaCSR[ 232 ][ 22 ],
   alphaCSR[ 232 ][ 23 ],
   alphaCSR[ 232 ][ 24 ],
   alphaCSR[ 232 ][ 25 ],
   alphaCSR[ 232 ][ 26 ],
   alphaCSR[ 232 ][ 27 ],
   alphaCSR[ 232 ][ 28 ],
   alphaCSR[ 232 ][ 29 ],
   alphaCSR[ 232 ][ 30 ],
   alphaCSR[ 232 ][ 31 ],
   alphaCSR[ 232 ][ 32 ],
   alphaCSR[ 232 ][ 33 ],
   alphaCSR[ 232 ][ 34 ],
   alphaCSR[ 232 ][ 35 ],
   alphaCSR[ 232 ][ 36 ],
   alphaCSR[ 232 ][ 37 ],
   alphaCSR[ 232 ][ 38 ],
   alphaCSR[ 232 ][ 39 ],
   alphaCSR[ 232 ][ 40 ],
   alphaCSR[ 232 ][ 41 ],
   alphaCSR[ 232 ][ 42 ],
   alphaCSR[ 232 ][ 43 ],
   alphaCSR[ 232 ][ 44 ],
   alphaCSR[ 232 ][ 45 ],
   alphaCSR[ 232 ][ 46 ],
   alphaCSR[ 232 ][ 47 ],
   alphaCSR[ 232 ][ 48 ],
   alphaCSR[ 232 ][ 49 ],
   alphaCSR[ 232 ][ 50 ],
   alphaCSR[ 232 ][ 51 ],
   alphaCSR[ 232 ][ 52 ],
   alphaCSR[ 232 ][ 53 ],
   alphaCSR[ 232 ][ 54 ],
   alphaCSR[ 232 ][ 55 ],
   alphaCSR[ 232 ][ 56 ],
   alphaCSR[ 232 ][ 57 ],
   alphaCSR[ 232 ][ 58 ],
   alphaCSR[ 232 ][ 59 ],
   alphaCSR[ 232 ][ 60 ],
   alphaCSR[ 232 ][ 61 ],
   alphaCSR[ 232 ][ 62 ],
   alphaCSR[ 232 ][ 63 ],
   alphaCSR[ 232 ][ 64 ],
   alphaCSR[ 232 ][ 65 ],
   alphaCSR[ 232 ][ 66 ],
   alphaCSR[ 232 ][ 67 ],
   alphaCSR[ 232 ][ 68 ],
   alphaCSR[ 232 ][ 69 ],
   alphaCSR[ 232 ][ 70 ],
   alphaCSR[ 232 ][ 71 ],
   alphaCSR[ 232 ][ 72 ],
   alphaCSR[ 232 ][ 73 ],
   alphaCSR[ 232 ][ 74 ],
   alphaCSR[ 232 ][ 75 ],
   alphaCSR[ 232 ][ 76 ],
   alphaCSR[ 232 ][ 77 ],
   alphaCSR[ 232 ][ 78 ],
   alphaCSR[ 232 ][ 79 ],
   alphaCSR[ 232 ][ 80 ],
   alphaCSR[ 232 ][ 81 ],
   alphaCSR[ 232 ][ 82 ],
   alphaCSR[ 232 ][ 83 ],
   alphaCSR[ 232 ][ 84 ],
   alphaCSR[ 232 ][ 85 ],
   alphaCSR[ 232 ][ 86 ],
   alphaCSR[ 232 ][ 87 ],
   alphaCSR[ 232 ][ 88 ],
   alphaCSR[ 232 ][ 89 ],
   alphaCSR[ 232 ][ 90 ],
   alphaCSR[ 232 ][ 91 ],
   alphaCSR[ 232 ][ 92 ],
   alphaCSR[ 232 ][ 93 ],
   alphaCSR[ 232 ][ 94 ],
   alphaCSR[ 232 ][ 95 ],
   alphaCSR[ 232 ][ 96 ],
   alphaCSR[ 232 ][ 97 ],
   alphaCSR[ 232 ][ 98 ],
   alphaCSR[ 232 ][ 99 ],
   alphaCSR[ 232 ][ 100 ],
   alphaCSR[ 232 ][ 101 ],
   alphaCSR[ 232 ][ 102 ],
   alphaCSR[ 232 ][ 103 ],
   alphaCSR[ 232 ][ 104 ],
   alphaCSR[ 232 ][ 105 ],
   alphaCSR[ 232 ][ 106 ],
   alphaCSR[ 232 ][ 107 ],
   alphaCSR[ 232 ][ 108 ],
   alphaCSR[ 232 ][ 109 ],
   alphaCSR[ 232 ][ 110 ],
   alphaCSR[ 232 ][ 111 ],
   alphaCSR[ 232 ][ 112 ],
   alphaCSR[ 232 ][ 113 ],
   alphaCSR[ 232 ][ 114 ],
   alphaCSR[ 232 ][ 115 ],
   alphaCSR[ 232 ][ 116 ],
   alphaCSR[ 232 ][ 117 ],
   alphaCSR[ 232 ][ 118 ],
   alphaCSR[ 232 ][ 119 ],
   alphaCSR[ 232 ][ 120 ],
   alphaCSR[ 232 ][ 121 ],
   alphaCSR[ 232 ][ 122 ],
   alphaCSR[ 232 ][ 123 ],
   alphaCSR[ 232 ][ 124 ],
   alphaCSR[ 232 ][ 125 ],
   alphaCSR[ 232 ][ 126 ],
   alphaCSR[ 232 ][ 127 ],
   alphaCSR[ 232 ][ 128 ],
   alphaCSR[ 232 ][ 129 ],
   alphaCSR[ 232 ][ 130 ],
   alphaCSR[ 232 ][ 131 ],
   alphaCSR[ 232 ][ 132 ],
   alphaCSR[ 232 ][ 133 ],
   alphaCSR[ 232 ][ 134 ],
   alphaCSR[ 232 ][ 135 ],
   alphaCSR[ 232 ][ 136 ],
   alphaCSR[ 232 ][ 137 ],
   alphaCSR[ 232 ][ 138 ],
   alphaCSR[ 232 ][ 139 ],
   alphaCSR[ 232 ][ 140 ],
   alphaCSR[ 232 ][ 141 ],
   alphaCSR[ 232 ][ 142 ],
   alphaCSR[ 232 ][ 143 ],
   alphaCSR[ 232 ][ 144 ],
   alphaCSR[ 232 ][ 145 ],
   alphaCSR[ 232 ][ 146 ],
   alphaCSR[ 232 ][ 147 ],
   alphaCSR[ 232 ][ 148 ],
   alphaCSR[ 232 ][ 149 ],
   alphaCSR[ 232 ][ 150 ],
   alphaCSR[ 232 ][ 151 ],
   alphaCSR[ 232 ][ 152 ],
   alphaCSR[ 232 ][ 153 ],
   alphaCSR[ 232 ][ 154 ],
   alphaCSR[ 232 ][ 155 ],
   alphaCSR[ 232 ][ 156 ],
   alphaCSR[ 232 ][ 157 ],
   alphaCSR[ 232 ][ 158 ],
   alphaCSR[ 232 ][ 159 ],
   alphaCSR[ 232 ][ 160 ],
   alphaCSR[ 232 ][ 161 ],
   alphaCSR[ 232 ][ 162 ],
   alphaCSR[ 232 ][ 163 ],
   alphaCSR[ 232 ][ 164 ],
   alphaCSR[ 232 ][ 165 ],
   alphaCSR[ 232 ][ 166 ],
   alphaCSR[ 232 ][ 167 ],
   alphaCSR[ 232 ][ 168 ],
   alphaCSR[ 232 ][ 169 ],
   alphaCSR[ 232 ][ 170 ],
   alphaCSR[ 232 ][ 171 ],
   alphaCSR[ 232 ][ 172 ],
   alphaCSR[ 232 ][ 173 ],
   alphaCSR[ 232 ][ 174 ],
   alphaCSR[ 232 ][ 175 ],
   alphaCSR[ 232 ][ 176 ],
   alphaCSR[ 232 ][ 177 ],
   alphaCSR[ 232 ][ 178 ],
   alphaCSR[ 232 ][ 179 ],
   alphaCSR[ 232 ][ 180 ],
   alphaCSR[ 232 ][ 181 ],
   alphaCSR[ 232 ][ 182 ],
   alphaCSR[ 232 ][ 183 ],
   alphaCSR[ 232 ][ 184 ],
   alphaCSR[ 232 ][ 185 ],
   alphaCSR[ 232 ][ 186 ],
   alphaCSR[ 232 ][ 187 ],
   alphaCSR[ 232 ][ 188 ],
   alphaCSR[ 232 ][ 189 ],
   alphaCSR[ 232 ][ 190 ],
   alphaCSR[ 232 ][ 191 ],
   alphaCSR[ 232 ][ 192 ],
   alphaCSR[ 232 ][ 193 ],
   alphaCSR[ 232 ][ 194 ],
   alphaCSR[ 232 ][ 195 ],
   alphaCSR[ 232 ][ 196 ],
   alphaCSR[ 232 ][ 197 ],
   alphaCSR[ 232 ][ 198 ],
   alphaCSR[ 232 ][ 199 ],
   alphaCSR[ 232 ][ 200 ],
   alphaCSR[ 232 ][ 201 ],
   alphaCSR[ 232 ][ 202 ],
   alphaCSR[ 232 ][ 203 ],
   alphaCSR[ 232 ][ 204 ],
   alphaCSR[ 232 ][ 205 ],
   alphaCSR[ 232 ][ 206 ],
   alphaCSR[ 232 ][ 207 ],
   alphaCSR[ 232 ][ 208 ],
   alphaCSR[ 232 ][ 209 ],
   alphaCSR[ 232 ][ 210 ],
   alphaCSR[ 232 ][ 211 ],
   alphaCSR[ 232 ][ 212 ],
   alphaCSR[ 232 ][ 213 ],
   alphaCSR[ 232 ][ 214 ],
   alphaCSR[ 232 ][ 215 ],
   alphaCSR[ 232 ][ 216 ],
   alphaCSR[ 232 ][ 217 ],
   alphaCSR[ 232 ][ 218 ],
   alphaCSR[ 232 ][ 219 ],
   alphaCSR[ 232 ][ 220 ],
   alphaCSR[ 232 ][ 221 ],
   alphaCSR[ 232 ][ 222 ],
   alphaCSR[ 232 ][ 223 ],
   alphaCSR[ 232 ][ 224 ],
   alphaCSR[ 232 ][ 225 ],
   alphaCSR[ 232 ][ 226 ],
   alphaCSR[ 232 ][ 227 ],
   alphaCSR[ 232 ][ 228 ],
   alphaCSR[ 232 ][ 229 ],
   alphaCSR[ 232 ][ 230 ],
   alphaCSR[ 232 ][ 231 ],
   alphaCSR[ 232 ][ 232 ],
   alphaCSR[ 232 ][ 233 ],
   alphaCSR[ 232 ][ 234 ],
   alphaCSR[ 232 ][ 235 ],
   alphaCSR[ 232 ][ 236 ],
   alphaCSR[ 232 ][ 237 ],
   alphaCSR[ 232 ][ 238 ],
   alphaCSR[ 232 ][ 239 ],
   alphaCSR[ 232 ][ 240 ],
   alphaCSR[ 232 ][ 241 ],
   alphaCSR[ 232 ][ 242 ],
   alphaCSR[ 232 ][ 243 ],
   alphaCSR[ 232 ][ 244 ],
   alphaCSR[ 232 ][ 245 ],
   alphaCSR[ 232 ][ 246 ],
   alphaCSR[ 232 ][ 247 ],
   alphaCSR[ 232 ][ 248 ],
   alphaCSR[ 232 ][ 249 ],
   alphaCSR[ 232 ][ 250 ],
   alphaCSR[ 232 ][ 251 ],
   alphaCSR[ 232 ][ 252 ],
   alphaCSR[ 232 ][ 253 ],
   alphaCSR[ 232 ][ 254 ],
   alphaCSR[ 232 ][ 255 ],
   alphaCSR[ 232 ][ 256 ],
   alphaCSR[ 232 ][ 257 ],
   alphaCSR[ 232 ][ 258 ],
   alphaCSR[ 232 ][ 259 ],
   alphaCSR[ 232 ][ 260 ],
   alphaCSR[ 232 ][ 261 ],
   alphaCSR[ 232 ][ 262 ],
   alphaCSR[ 232 ][ 263 ],
   alphaCSR[ 232 ][ 264 ],
   alphaCSR[ 232 ][ 265 ],
   alphaCSR[ 232 ][ 266 ],
   alphaCSR[ 232 ][ 267 ],
   alphaCSR[ 232 ][ 268 ],
   alphaCSR[ 232 ][ 269 ],
   alphaCSR[ 232 ][ 270 ],
   alphaCSR[ 232 ][ 271 ],
   alphaCSR[ 232 ][ 272 ],
   alphaCSR[ 232 ][ 273 ],
   alphaCSR[ 232 ][ 274 ],
   alphaCSR[ 232 ][ 275 ],
   alphaCSR[ 232 ][ 276 ],
   alphaCSR[ 232 ][ 277 ],
   alphaCSR[ 232 ][ 278 ],
   alphaCSR[ 232 ][ 279 ],
   alphaCSR[ 232 ][ 280 ],
   alphaCSR[ 232 ][ 281 ],
   alphaCSR[ 232 ][ 282 ],
   alphaCSR[ 232 ][ 283 ],
   alphaCSR[ 232 ][ 284 ],
   alphaCSR[ 232 ][ 285 ],
   alphaCSR[ 232 ][ 286 ],
   alphaCSR[ 232 ][ 287 ],
   alphaCSR[ 232 ][ 288 ],
   alphaCSR[ 232 ][ 289 ],
   alphaCSR[ 232 ][ 290 ],
   alphaCSR[ 232 ][ 291 ],
   alphaCSR[ 232 ][ 292 ],
   alphaCSR[ 232 ][ 293 ],
   alphaCSR[ 232 ][ 294 ],
   alphaCSR[ 232 ][ 295 ],
   alphaCSR[ 232 ][ 296 ],
   alphaCSR[ 232 ][ 297 ],
   alphaCSR[ 232 ][ 298 ],
   alphaCSR[ 232 ][ 299 ],
   alphaCSR[ 232 ][ 300 ],
   alphaCSR[ 232 ][ 301 ],
   alphaCSR[ 232 ][ 302 ],
   alphaCSR[ 232 ][ 303 ],
   alphaCSR[ 232 ][ 304 ],
   alphaCSR[ 232 ][ 305 ],
   alphaCSR[ 232 ][ 306 ],
   alphaCSR[ 232 ][ 307 ],
   alphaCSR[ 232 ][ 308 ],
   alphaCSR[ 232 ][ 309 ],
   alphaCSR[ 232 ][ 310 ],
   alphaCSR[ 232 ][ 311 ],
   alphaCSR[ 232 ][ 312 ],
   alphaCSR[ 232 ][ 313 ],
   alphaCSR[ 232 ][ 314 ],
   alphaCSR[ 232 ][ 315 ],
   alphaCSR[ 232 ][ 316 ],
   alphaCSR[ 232 ][ 317 ],
   alphaCSR[ 232 ][ 318 ],
   alphaCSR[ 232 ][ 319 ],
   alphaCSR[ 232 ][ 320 ],
   alphaCSR[ 232 ][ 321 ],
   alphaCSR[ 232 ][ 322 ],
   alphaCSR[ 232 ][ 323 ],
   alphaCSR[ 232 ][ 324 ],
   alphaCSR[ 232 ][ 325 ],
   alphaCSR[ 232 ][ 326 ],
   alphaCSR[ 232 ][ 327 ],
   alphaCSR[ 232 ][ 328 ],
   alphaCSR[ 232 ][ 329 ],
   alphaCSR[ 232 ][ 330 ],
   alphaCSR[ 232 ][ 331 ],
   alphaCSR[ 232 ][ 332 ],
   alphaCSR[ 232 ][ 333 ],
   alphaCSR[ 232 ][ 334 ],
   alphaCSR[ 232 ][ 335 ],
   alphaCSR[ 232 ][ 336 ],
   alphaCSR[ 232 ][ 337 ],
   alphaCSR[ 232 ][ 338 ],
   alphaCSR[ 232 ][ 339 ],
   alphaCSR[ 232 ][ 340 ],
   alphaCSR[ 232 ][ 341 ],
   alphaCSR[ 232 ][ 342 ],
   alphaCSR[ 232 ][ 343 ],
   alphaCSR[ 232 ][ 344 ],
   alphaCSR[ 232 ][ 345 ],
   alphaCSR[ 232 ][ 346 ],
   alphaCSR[ 232 ][ 347 ],
   alphaCSR[ 232 ][ 348 ],
   alphaCSR[ 232 ][ 349 ],
   alphaCSR[ 232 ][ 350 ],
   alphaCSR[ 232 ][ 351 ],
   alphaCSR[ 232 ][ 352 ],
   alphaCSR[ 232 ][ 353 ],
   alphaCSR[ 232 ][ 354 ],
   alphaCSR[ 232 ][ 355 ],
   alphaCSR[ 232 ][ 356 ],
   alphaCSR[ 232 ][ 357 ],
   alphaCSR[ 232 ][ 358 ],
   alphaCSR[ 232 ][ 359 ],
   alphaCSR[ 232 ][ 360 ],
   alphaCSR[ 232 ][ 361 ],
   alphaCSR[ 232 ][ 362 ],
   alphaCSR[ 232 ][ 363 ],
   alphaCSR[ 232 ][ 364 ],
   alphaCSR[ 232 ][ 365 ],
   alphaCSR[ 232 ][ 366 ],
   alphaCSR[ 232 ][ 367 ],
   alphaCSR[ 232 ][ 368 ],
   alphaCSR[ 232 ][ 369 ],
   alphaCSR[ 232 ][ 370 ],
   alphaCSR[ 232 ][ 371 ],
   alphaCSR[ 232 ][ 372 ],
   alphaCSR[ 232 ][ 373 ],
   alphaCSR[ 232 ][ 374 ],
   alphaCSR[ 232 ][ 375 ],
   alphaCSR[ 232 ][ 376 ],
   alphaCSR[ 232 ][ 377 ],
   alphaCSR[ 232 ][ 378 ],
   alphaCSR[ 232 ][ 379 ],
   alphaCSR[ 232 ][ 380 ],
   alphaCSR[ 232 ][ 381 ],
   alphaCSR[ 232 ][ 382 ],
   alphaCSR[ 232 ][ 383 ],
   alphaCSR[ 233 ][ 0 ],
   alphaCSR[ 233 ][ 1 ],
   alphaCSR[ 233 ][ 2 ],
   alphaCSR[ 233 ][ 3 ],
   alphaCSR[ 233 ][ 4 ],
   alphaCSR[ 233 ][ 5 ],
   alphaCSR[ 233 ][ 6 ],
   alphaCSR[ 233 ][ 7 ],
   alphaCSR[ 233 ][ 8 ],
   alphaCSR[ 233 ][ 9 ],
   alphaCSR[ 233 ][ 10 ],
   alphaCSR[ 233 ][ 11 ],
   alphaCSR[ 233 ][ 12 ],
   alphaCSR[ 233 ][ 13 ],
   alphaCSR[ 233 ][ 14 ],
   alphaCSR[ 233 ][ 15 ],
   alphaCSR[ 233 ][ 16 ],
   alphaCSR[ 233 ][ 17 ],
   alphaCSR[ 233 ][ 18 ],
   alphaCSR[ 233 ][ 19 ],
   alphaCSR[ 233 ][ 20 ],
   alphaCSR[ 233 ][ 21 ],
   alphaCSR[ 233 ][ 22 ],
   alphaCSR[ 233 ][ 23 ],
   alphaCSR[ 233 ][ 24 ],
   alphaCSR[ 233 ][ 25 ],
   alphaCSR[ 233 ][ 26 ],
   alphaCSR[ 233 ][ 27 ],
   alphaCSR[ 233 ][ 28 ],
   alphaCSR[ 233 ][ 29 ],
   alphaCSR[ 233 ][ 30 ],
   alphaCSR[ 233 ][ 31 ],
   alphaCSR[ 233 ][ 32 ],
   alphaCSR[ 233 ][ 33 ],
   alphaCSR[ 233 ][ 34 ],
   alphaCSR[ 233 ][ 35 ],
   alphaCSR[ 233 ][ 36 ],
   alphaCSR[ 233 ][ 37 ],
   alphaCSR[ 233 ][ 38 ],
   alphaCSR[ 233 ][ 39 ],
   alphaCSR[ 233 ][ 40 ],
   alphaCSR[ 233 ][ 41 ],
   alphaCSR[ 233 ][ 42 ],
   alphaCSR[ 233 ][ 43 ],
   alphaCSR[ 233 ][ 44 ],
   alphaCSR[ 233 ][ 45 ],
   alphaCSR[ 233 ][ 46 ],
   alphaCSR[ 233 ][ 47 ],
   alphaCSR[ 233 ][ 48 ],
   alphaCSR[ 233 ][ 49 ],
   alphaCSR[ 233 ][ 50 ],
   alphaCSR[ 233 ][ 51 ],
   alphaCSR[ 233 ][ 52 ],
   alphaCSR[ 233 ][ 53 ],
   alphaCSR[ 233 ][ 54 ],
   alphaCSR[ 233 ][ 55 ],
   alphaCSR[ 233 ][ 56 ],
   alphaCSR[ 233 ][ 57 ],
   alphaCSR[ 233 ][ 58 ],
   alphaCSR[ 233 ][ 59 ],
   alphaCSR[ 233 ][ 60 ],
   alphaCSR[ 233 ][ 61 ],
   alphaCSR[ 233 ][ 62 ],
   alphaCSR[ 233 ][ 63 ],
   alphaCSR[ 233 ][ 64 ],
   alphaCSR[ 233 ][ 65 ],
   alphaCSR[ 233 ][ 66 ],
   alphaCSR[ 233 ][ 67 ],
   alphaCSR[ 233 ][ 68 ],
   alphaCSR[ 233 ][ 69 ],
   alphaCSR[ 233 ][ 70 ],
   alphaCSR[ 233 ][ 71 ],
   alphaCSR[ 233 ][ 72 ],
   alphaCSR[ 233 ][ 73 ],
   alphaCSR[ 233 ][ 74 ],
   alphaCSR[ 233 ][ 75 ],
   alphaCSR[ 233 ][ 76 ],
   alphaCSR[ 233 ][ 77 ],
   alphaCSR[ 233 ][ 78 ],
   alphaCSR[ 233 ][ 79 ],
   alphaCSR[ 233 ][ 80 ],
   alphaCSR[ 233 ][ 81 ],
   alphaCSR[ 233 ][ 82 ],
   alphaCSR[ 233 ][ 83 ],
   alphaCSR[ 233 ][ 84 ],
   alphaCSR[ 233 ][ 85 ],
   alphaCSR[ 233 ][ 86 ],
   alphaCSR[ 233 ][ 87 ],
   alphaCSR[ 233 ][ 88 ],
   alphaCSR[ 233 ][ 89 ],
   alphaCSR[ 233 ][ 90 ],
   alphaCSR[ 233 ][ 91 ],
   alphaCSR[ 233 ][ 92 ],
   alphaCSR[ 233 ][ 93 ],
   alphaCSR[ 233 ][ 94 ],
   alphaCSR[ 233 ][ 95 ],
   alphaCSR[ 233 ][ 96 ],
   alphaCSR[ 233 ][ 97 ],
   alphaCSR[ 233 ][ 98 ],
   alphaCSR[ 233 ][ 99 ],
   alphaCSR[ 233 ][ 100 ],
   alphaCSR[ 233 ][ 101 ],
   alphaCSR[ 233 ][ 102 ],
   alphaCSR[ 233 ][ 103 ],
   alphaCSR[ 233 ][ 104 ],
   alphaCSR[ 233 ][ 105 ],
   alphaCSR[ 233 ][ 106 ],
   alphaCSR[ 233 ][ 107 ],
   alphaCSR[ 233 ][ 108 ],
   alphaCSR[ 233 ][ 109 ],
   alphaCSR[ 233 ][ 110 ],
   alphaCSR[ 233 ][ 111 ],
   alphaCSR[ 233 ][ 112 ],
   alphaCSR[ 233 ][ 113 ],
   alphaCSR[ 233 ][ 114 ],
   alphaCSR[ 233 ][ 115 ],
   alphaCSR[ 233 ][ 116 ],
   alphaCSR[ 233 ][ 117 ],
   alphaCSR[ 233 ][ 118 ],
   alphaCSR[ 233 ][ 119 ],
   alphaCSR[ 233 ][ 120 ],
   alphaCSR[ 233 ][ 121 ],
   alphaCSR[ 233 ][ 122 ],
   alphaCSR[ 233 ][ 123 ],
   alphaCSR[ 233 ][ 124 ],
   alphaCSR[ 233 ][ 125 ],
   alphaCSR[ 233 ][ 126 ],
   alphaCSR[ 233 ][ 127 ],
   alphaCSR[ 233 ][ 128 ],
   alphaCSR[ 233 ][ 129 ],
   alphaCSR[ 233 ][ 130 ],
   alphaCSR[ 233 ][ 131 ],
   alphaCSR[ 233 ][ 132 ],
   alphaCSR[ 233 ][ 133 ],
   alphaCSR[ 233 ][ 134 ],
   alphaCSR[ 233 ][ 135 ],
   alphaCSR[ 233 ][ 136 ],
   alphaCSR[ 233 ][ 137 ],
   alphaCSR[ 233 ][ 138 ],
   alphaCSR[ 233 ][ 139 ],
   alphaCSR[ 233 ][ 140 ],
   alphaCSR[ 233 ][ 141 ],
   alphaCSR[ 233 ][ 142 ],
   alphaCSR[ 233 ][ 143 ],
   alphaCSR[ 233 ][ 144 ],
   alphaCSR[ 233 ][ 145 ],
   alphaCSR[ 233 ][ 146 ],
   alphaCSR[ 233 ][ 147 ],
   alphaCSR[ 233 ][ 148 ],
   alphaCSR[ 233 ][ 149 ],
   alphaCSR[ 233 ][ 150 ],
   alphaCSR[ 233 ][ 151 ],
   alphaCSR[ 233 ][ 152 ],
   alphaCSR[ 233 ][ 153 ],
   alphaCSR[ 233 ][ 154 ],
   alphaCSR[ 233 ][ 155 ],
   alphaCSR[ 233 ][ 156 ],
   alphaCSR[ 233 ][ 157 ],
   alphaCSR[ 233 ][ 158 ],
   alphaCSR[ 233 ][ 159 ],
   alphaCSR[ 233 ][ 160 ],
   alphaCSR[ 233 ][ 161 ],
   alphaCSR[ 233 ][ 162 ],
   alphaCSR[ 233 ][ 163 ],
   alphaCSR[ 233 ][ 164 ],
   alphaCSR[ 233 ][ 165 ],
   alphaCSR[ 233 ][ 166 ],
   alphaCSR[ 233 ][ 167 ],
   alphaCSR[ 233 ][ 168 ],
   alphaCSR[ 233 ][ 169 ],
   alphaCSR[ 233 ][ 170 ],
   alphaCSR[ 233 ][ 171 ],
   alphaCSR[ 233 ][ 172 ],
   alphaCSR[ 233 ][ 173 ],
   alphaCSR[ 233 ][ 174 ],
   alphaCSR[ 233 ][ 175 ],
   alphaCSR[ 233 ][ 176 ],
   alphaCSR[ 233 ][ 177 ],
   alphaCSR[ 233 ][ 178 ],
   alphaCSR[ 233 ][ 179 ],
   alphaCSR[ 233 ][ 180 ],
   alphaCSR[ 233 ][ 181 ],
   alphaCSR[ 233 ][ 182 ],
   alphaCSR[ 233 ][ 183 ],
   alphaCSR[ 233 ][ 184 ],
   alphaCSR[ 233 ][ 185 ],
   alphaCSR[ 233 ][ 186 ],
   alphaCSR[ 233 ][ 187 ],
   alphaCSR[ 233 ][ 188 ],
   alphaCSR[ 233 ][ 189 ],
   alphaCSR[ 233 ][ 190 ],
   alphaCSR[ 233 ][ 191 ],
   alphaCSR[ 233 ][ 192 ],
   alphaCSR[ 233 ][ 193 ],
   alphaCSR[ 233 ][ 194 ],
   alphaCSR[ 233 ][ 195 ],
   alphaCSR[ 233 ][ 196 ],
   alphaCSR[ 233 ][ 197 ],
   alphaCSR[ 233 ][ 198 ],
   alphaCSR[ 233 ][ 199 ],
   alphaCSR[ 233 ][ 200 ],
   alphaCSR[ 233 ][ 201 ],
   alphaCSR[ 233 ][ 202 ],
   alphaCSR[ 233 ][ 203 ],
   alphaCSR[ 233 ][ 204 ],
   alphaCSR[ 233 ][ 205 ],
   alphaCSR[ 233 ][ 206 ],
   alphaCSR[ 233 ][ 207 ],
   alphaCSR[ 233 ][ 208 ],
   alphaCSR[ 233 ][ 209 ],
   alphaCSR[ 233 ][ 210 ],
   alphaCSR[ 233 ][ 211 ],
   alphaCSR[ 233 ][ 212 ],
   alphaCSR[ 233 ][ 213 ],
   alphaCSR[ 233 ][ 214 ],
   alphaCSR[ 233 ][ 215 ],
   alphaCSR[ 233 ][ 216 ],
   alphaCSR[ 233 ][ 217 ],
   alphaCSR[ 233 ][ 218 ],
   alphaCSR[ 233 ][ 219 ],
   alphaCSR[ 233 ][ 220 ],
   alphaCSR[ 233 ][ 221 ],
   alphaCSR[ 233 ][ 222 ],
   alphaCSR[ 233 ][ 223 ],
   alphaCSR[ 233 ][ 224 ],
   alphaCSR[ 233 ][ 225 ],
   alphaCSR[ 233 ][ 226 ],
   alphaCSR[ 233 ][ 227 ],
   alphaCSR[ 233 ][ 228 ],
   alphaCSR[ 233 ][ 229 ],
   alphaCSR[ 233 ][ 230 ],
   alphaCSR[ 233 ][ 231 ],
   alphaCSR[ 233 ][ 232 ],
   alphaCSR[ 233 ][ 233 ],
   alphaCSR[ 233 ][ 234 ],
   alphaCSR[ 233 ][ 235 ],
   alphaCSR[ 233 ][ 236 ],
   alphaCSR[ 233 ][ 237 ],
   alphaCSR[ 233 ][ 238 ],
   alphaCSR[ 233 ][ 239 ],
   alphaCSR[ 233 ][ 240 ],
   alphaCSR[ 233 ][ 241 ],
   alphaCSR[ 233 ][ 242 ],
   alphaCSR[ 233 ][ 243 ],
   alphaCSR[ 233 ][ 244 ],
   alphaCSR[ 233 ][ 245 ],
   alphaCSR[ 233 ][ 246 ],
   alphaCSR[ 233 ][ 247 ],
   alphaCSR[ 233 ][ 248 ],
   alphaCSR[ 233 ][ 249 ],
   alphaCSR[ 233 ][ 250 ],
   alphaCSR[ 233 ][ 251 ],
   alphaCSR[ 233 ][ 252 ],
   alphaCSR[ 233 ][ 253 ],
   alphaCSR[ 233 ][ 254 ],
   alphaCSR[ 233 ][ 255 ],
   alphaCSR[ 233 ][ 256 ],
   alphaCSR[ 233 ][ 257 ],
   alphaCSR[ 233 ][ 258 ],
   alphaCSR[ 233 ][ 259 ],
   alphaCSR[ 233 ][ 260 ],
   alphaCSR[ 233 ][ 261 ],
   alphaCSR[ 233 ][ 262 ],
   alphaCSR[ 233 ][ 263 ],
   alphaCSR[ 233 ][ 264 ],
   alphaCSR[ 233 ][ 265 ],
   alphaCSR[ 233 ][ 266 ],
   alphaCSR[ 233 ][ 267 ],
   alphaCSR[ 233 ][ 268 ],
   alphaCSR[ 233 ][ 269 ],
   alphaCSR[ 233 ][ 270 ],
   alphaCSR[ 233 ][ 271 ],
   alphaCSR[ 233 ][ 272 ],
   alphaCSR[ 233 ][ 273 ],
   alphaCSR[ 233 ][ 274 ],
   alphaCSR[ 233 ][ 275 ],
   alphaCSR[ 233 ][ 276 ],
   alphaCSR[ 233 ][ 277 ],
   alphaCSR[ 233 ][ 278 ],
   alphaCSR[ 233 ][ 279 ],
   alphaCSR[ 233 ][ 280 ],
   alphaCSR[ 233 ][ 281 ],
   alphaCSR[ 233 ][ 282 ],
   alphaCSR[ 233 ][ 283 ],
   alphaCSR[ 233 ][ 284 ],
   alphaCSR[ 233 ][ 285 ],
   alphaCSR[ 233 ][ 286 ],
   alphaCSR[ 233 ][ 287 ],
   alphaCSR[ 233 ][ 288 ],
   alphaCSR[ 233 ][ 289 ],
   alphaCSR[ 233 ][ 290 ],
   alphaCSR[ 233 ][ 291 ],
   alphaCSR[ 233 ][ 292 ],
   alphaCSR[ 233 ][ 293 ],
   alphaCSR[ 233 ][ 294 ],
   alphaCSR[ 233 ][ 295 ],
   alphaCSR[ 233 ][ 296 ],
   alphaCSR[ 233 ][ 297 ],
   alphaCSR[ 233 ][ 298 ],
   alphaCSR[ 233 ][ 299 ],
   alphaCSR[ 233 ][ 300 ],
   alphaCSR[ 233 ][ 301 ],
   alphaCSR[ 233 ][ 302 ],
   alphaCSR[ 233 ][ 303 ],
   alphaCSR[ 233 ][ 304 ],
   alphaCSR[ 233 ][ 305 ],
   alphaCSR[ 233 ][ 306 ],
   alphaCSR[ 233 ][ 307 ],
   alphaCSR[ 233 ][ 308 ],
   alphaCSR[ 233 ][ 309 ],
   alphaCSR[ 233 ][ 310 ],
   alphaCSR[ 233 ][ 311 ],
   alphaCSR[ 233 ][ 312 ],
   alphaCSR[ 233 ][ 313 ],
   alphaCSR[ 233 ][ 314 ],
   alphaCSR[ 233 ][ 315 ],
   alphaCSR[ 233 ][ 316 ],
   alphaCSR[ 233 ][ 317 ],
   alphaCSR[ 233 ][ 318 ],
   alphaCSR[ 233 ][ 319 ],
   alphaCSR[ 233 ][ 320 ],
   alphaCSR[ 233 ][ 321 ],
   alphaCSR[ 233 ][ 322 ],
   alphaCSR[ 233 ][ 323 ],
   alphaCSR[ 233 ][ 324 ],
   alphaCSR[ 233 ][ 325 ],
   alphaCSR[ 233 ][ 326 ],
   alphaCSR[ 233 ][ 327 ],
   alphaCSR[ 233 ][ 328 ],
   alphaCSR[ 233 ][ 329 ],
   alphaCSR[ 233 ][ 330 ],
   alphaCSR[ 233 ][ 331 ],
   alphaCSR[ 233 ][ 332 ],
   alphaCSR[ 233 ][ 333 ],
   alphaCSR[ 233 ][ 334 ],
   alphaCSR[ 233 ][ 335 ],
   alphaCSR[ 233 ][ 336 ],
   alphaCSR[ 233 ][ 337 ],
   alphaCSR[ 233 ][ 338 ],
   alphaCSR[ 233 ][ 339 ],
   alphaCSR[ 233 ][ 340 ],
   alphaCSR[ 233 ][ 341 ],
   alphaCSR[ 233 ][ 342 ],
   alphaCSR[ 233 ][ 343 ],
   alphaCSR[ 233 ][ 344 ],
   alphaCSR[ 233 ][ 345 ],
   alphaCSR[ 233 ][ 346 ],
   alphaCSR[ 233 ][ 347 ],
   alphaCSR[ 233 ][ 348 ],
   alphaCSR[ 233 ][ 349 ],
   alphaCSR[ 233 ][ 350 ],
   alphaCSR[ 233 ][ 351 ],
   alphaCSR[ 233 ][ 352 ],
   alphaCSR[ 233 ][ 353 ],
   alphaCSR[ 233 ][ 354 ],
   alphaCSR[ 233 ][ 355 ],
   alphaCSR[ 233 ][ 356 ],
   alphaCSR[ 233 ][ 357 ],
   alphaCSR[ 233 ][ 358 ],
   alphaCSR[ 233 ][ 359 ],
   alphaCSR[ 233 ][ 360 ],
   alphaCSR[ 233 ][ 361 ],
   alphaCSR[ 233 ][ 362 ],
   alphaCSR[ 233 ][ 363 ],
   alphaCSR[ 233 ][ 364 ],
   alphaCSR[ 233 ][ 365 ],
   alphaCSR[ 233 ][ 366 ],
   alphaCSR[ 233 ][ 367 ],
   alphaCSR[ 233 ][ 368 ],
   alphaCSR[ 233 ][ 369 ],
   alphaCSR[ 233 ][ 370 ],
   alphaCSR[ 233 ][ 371 ],
   alphaCSR[ 233 ][ 372 ],
   alphaCSR[ 233 ][ 373 ],
   alphaCSR[ 233 ][ 374 ],
   alphaCSR[ 233 ][ 375 ],
   alphaCSR[ 233 ][ 376 ],
   alphaCSR[ 233 ][ 377 ],
   alphaCSR[ 233 ][ 378 ],
   alphaCSR[ 233 ][ 379 ],
   alphaCSR[ 233 ][ 380 ],
   alphaCSR[ 233 ][ 381 ],
   alphaCSR[ 233 ][ 382 ],
   alphaCSR[ 233 ][ 383 ],
   alphaCSR[ 234 ][ 0 ],
   alphaCSR[ 234 ][ 1 ],
   alphaCSR[ 234 ][ 2 ],
   alphaCSR[ 234 ][ 3 ],
   alphaCSR[ 234 ][ 4 ],
   alphaCSR[ 234 ][ 5 ],
   alphaCSR[ 234 ][ 6 ],
   alphaCSR[ 234 ][ 7 ],
   alphaCSR[ 234 ][ 8 ],
   alphaCSR[ 234 ][ 9 ],
   alphaCSR[ 234 ][ 10 ],
   alphaCSR[ 234 ][ 11 ],
   alphaCSR[ 234 ][ 12 ],
   alphaCSR[ 234 ][ 13 ],
   alphaCSR[ 234 ][ 14 ],
   alphaCSR[ 234 ][ 15 ],
   alphaCSR[ 234 ][ 16 ],
   alphaCSR[ 234 ][ 17 ],
   alphaCSR[ 234 ][ 18 ],
   alphaCSR[ 234 ][ 19 ],
   alphaCSR[ 234 ][ 20 ],
   alphaCSR[ 234 ][ 21 ],
   alphaCSR[ 234 ][ 22 ],
   alphaCSR[ 234 ][ 23 ],
   alphaCSR[ 234 ][ 24 ],
   alphaCSR[ 234 ][ 25 ],
   alphaCSR[ 234 ][ 26 ],
   alphaCSR[ 234 ][ 27 ],
   alphaCSR[ 234 ][ 28 ],
   alphaCSR[ 234 ][ 29 ],
   alphaCSR[ 234 ][ 30 ],
   alphaCSR[ 234 ][ 31 ],
   alphaCSR[ 234 ][ 32 ],
   alphaCSR[ 234 ][ 33 ],
   alphaCSR[ 234 ][ 34 ],
   alphaCSR[ 234 ][ 35 ],
   alphaCSR[ 234 ][ 36 ],
   alphaCSR[ 234 ][ 37 ],
   alphaCSR[ 234 ][ 38 ],
   alphaCSR[ 234 ][ 39 ],
   alphaCSR[ 234 ][ 40 ],
   alphaCSR[ 234 ][ 41 ],
   alphaCSR[ 234 ][ 42 ],
   alphaCSR[ 234 ][ 43 ],
   alphaCSR[ 234 ][ 44 ],
   alphaCSR[ 234 ][ 45 ],
   alphaCSR[ 234 ][ 46 ],
   alphaCSR[ 234 ][ 47 ],
   alphaCSR[ 234 ][ 48 ],
   alphaCSR[ 234 ][ 49 ],
   alphaCSR[ 234 ][ 50 ],
   alphaCSR[ 234 ][ 51 ],
   alphaCSR[ 234 ][ 52 ],
   alphaCSR[ 234 ][ 53 ],
   alphaCSR[ 234 ][ 54 ],
   alphaCSR[ 234 ][ 55 ],
   alphaCSR[ 234 ][ 56 ],
   alphaCSR[ 234 ][ 57 ],
   alphaCSR[ 234 ][ 58 ],
   alphaCSR[ 234 ][ 59 ],
   alphaCSR[ 234 ][ 60 ],
   alphaCSR[ 234 ][ 61 ],
   alphaCSR[ 234 ][ 62 ],
   alphaCSR[ 234 ][ 63 ],
   alphaCSR[ 234 ][ 64 ],
   alphaCSR[ 234 ][ 65 ],
   alphaCSR[ 234 ][ 66 ],
   alphaCSR[ 234 ][ 67 ],
   alphaCSR[ 234 ][ 68 ],
   alphaCSR[ 234 ][ 69 ],
   alphaCSR[ 234 ][ 70 ],
   alphaCSR[ 234 ][ 71 ],
   alphaCSR[ 234 ][ 72 ],
   alphaCSR[ 234 ][ 73 ],
   alphaCSR[ 234 ][ 74 ],
   alphaCSR[ 234 ][ 75 ],
   alphaCSR[ 234 ][ 76 ],
   alphaCSR[ 234 ][ 77 ],
   alphaCSR[ 234 ][ 78 ],
   alphaCSR[ 234 ][ 79 ],
   alphaCSR[ 234 ][ 80 ],
   alphaCSR[ 234 ][ 81 ],
   alphaCSR[ 234 ][ 82 ],
   alphaCSR[ 234 ][ 83 ],
   alphaCSR[ 234 ][ 84 ],
   alphaCSR[ 234 ][ 85 ],
   alphaCSR[ 234 ][ 86 ],
   alphaCSR[ 234 ][ 87 ],
   alphaCSR[ 234 ][ 88 ],
   alphaCSR[ 234 ][ 89 ],
   alphaCSR[ 234 ][ 90 ],
   alphaCSR[ 234 ][ 91 ],
   alphaCSR[ 234 ][ 92 ],
   alphaCSR[ 234 ][ 93 ],
   alphaCSR[ 234 ][ 94 ],
   alphaCSR[ 234 ][ 95 ],
   alphaCSR[ 234 ][ 96 ],
   alphaCSR[ 234 ][ 97 ],
   alphaCSR[ 234 ][ 98 ],
   alphaCSR[ 234 ][ 99 ],
   alphaCSR[ 234 ][ 100 ],
   alphaCSR[ 234 ][ 101 ],
   alphaCSR[ 234 ][ 102 ],
   alphaCSR[ 234 ][ 103 ],
   alphaCSR[ 234 ][ 104 ],
   alphaCSR[ 234 ][ 105 ],
   alphaCSR[ 234 ][ 106 ],
   alphaCSR[ 234 ][ 107 ],
   alphaCSR[ 234 ][ 108 ],
   alphaCSR[ 234 ][ 109 ],
   alphaCSR[ 234 ][ 110 ],
   alphaCSR[ 234 ][ 111 ],
   alphaCSR[ 234 ][ 112 ],
   alphaCSR[ 234 ][ 113 ],
   alphaCSR[ 234 ][ 114 ],
   alphaCSR[ 234 ][ 115 ],
   alphaCSR[ 234 ][ 116 ],
   alphaCSR[ 234 ][ 117 ],
   alphaCSR[ 234 ][ 118 ],
   alphaCSR[ 234 ][ 119 ],
   alphaCSR[ 234 ][ 120 ],
   alphaCSR[ 234 ][ 121 ],
   alphaCSR[ 234 ][ 122 ],
   alphaCSR[ 234 ][ 123 ],
   alphaCSR[ 234 ][ 124 ],
   alphaCSR[ 234 ][ 125 ],
   alphaCSR[ 234 ][ 126 ],
   alphaCSR[ 234 ][ 127 ],
   alphaCSR[ 234 ][ 128 ],
   alphaCSR[ 234 ][ 129 ],
   alphaCSR[ 234 ][ 130 ],
   alphaCSR[ 234 ][ 131 ],
   alphaCSR[ 234 ][ 132 ],
   alphaCSR[ 234 ][ 133 ],
   alphaCSR[ 234 ][ 134 ],
   alphaCSR[ 234 ][ 135 ],
   alphaCSR[ 234 ][ 136 ],
   alphaCSR[ 234 ][ 137 ],
   alphaCSR[ 234 ][ 138 ],
   alphaCSR[ 234 ][ 139 ],
   alphaCSR[ 234 ][ 140 ],
   alphaCSR[ 234 ][ 141 ],
   alphaCSR[ 234 ][ 142 ],
   alphaCSR[ 234 ][ 143 ],
   alphaCSR[ 234 ][ 144 ],
   alphaCSR[ 234 ][ 145 ],
   alphaCSR[ 234 ][ 146 ],
   alphaCSR[ 234 ][ 147 ],
   alphaCSR[ 234 ][ 148 ],
   alphaCSR[ 234 ][ 149 ],
   alphaCSR[ 234 ][ 150 ],
   alphaCSR[ 234 ][ 151 ],
   alphaCSR[ 234 ][ 152 ],
   alphaCSR[ 234 ][ 153 ],
   alphaCSR[ 234 ][ 154 ],
   alphaCSR[ 234 ][ 155 ],
   alphaCSR[ 234 ][ 156 ],
   alphaCSR[ 234 ][ 157 ],
   alphaCSR[ 234 ][ 158 ],
   alphaCSR[ 234 ][ 159 ],
   alphaCSR[ 234 ][ 160 ],
   alphaCSR[ 234 ][ 161 ],
   alphaCSR[ 234 ][ 162 ],
   alphaCSR[ 234 ][ 163 ],
   alphaCSR[ 234 ][ 164 ],
   alphaCSR[ 234 ][ 165 ],
   alphaCSR[ 234 ][ 166 ],
   alphaCSR[ 234 ][ 167 ],
   alphaCSR[ 234 ][ 168 ],
   alphaCSR[ 234 ][ 169 ],
   alphaCSR[ 234 ][ 170 ],
   alphaCSR[ 234 ][ 171 ],
   alphaCSR[ 234 ][ 172 ],
   alphaCSR[ 234 ][ 173 ],
   alphaCSR[ 234 ][ 174 ],
   alphaCSR[ 234 ][ 175 ],
   alphaCSR[ 234 ][ 176 ],
   alphaCSR[ 234 ][ 177 ],
   alphaCSR[ 234 ][ 178 ],
   alphaCSR[ 234 ][ 179 ],
   alphaCSR[ 234 ][ 180 ],
   alphaCSR[ 234 ][ 181 ],
   alphaCSR[ 234 ][ 182 ],
   alphaCSR[ 234 ][ 183 ],
   alphaCSR[ 234 ][ 184 ],
   alphaCSR[ 234 ][ 185 ],
   alphaCSR[ 234 ][ 186 ],
   alphaCSR[ 234 ][ 187 ],
   alphaCSR[ 234 ][ 188 ],
   alphaCSR[ 234 ][ 189 ],
   alphaCSR[ 234 ][ 190 ],
   alphaCSR[ 234 ][ 191 ],
   alphaCSR[ 234 ][ 192 ],
   alphaCSR[ 234 ][ 193 ],
   alphaCSR[ 234 ][ 194 ],
   alphaCSR[ 234 ][ 195 ],
   alphaCSR[ 234 ][ 196 ],
   alphaCSR[ 234 ][ 197 ],
   alphaCSR[ 234 ][ 198 ],
   alphaCSR[ 234 ][ 199 ],
   alphaCSR[ 234 ][ 200 ],
   alphaCSR[ 234 ][ 201 ],
   alphaCSR[ 234 ][ 202 ],
   alphaCSR[ 234 ][ 203 ],
   alphaCSR[ 234 ][ 204 ],
   alphaCSR[ 234 ][ 205 ],
   alphaCSR[ 234 ][ 206 ],
   alphaCSR[ 234 ][ 207 ],
   alphaCSR[ 234 ][ 208 ],
   alphaCSR[ 234 ][ 209 ],
   alphaCSR[ 234 ][ 210 ],
   alphaCSR[ 234 ][ 211 ],
   alphaCSR[ 234 ][ 212 ],
   alphaCSR[ 234 ][ 213 ],
   alphaCSR[ 234 ][ 214 ],
   alphaCSR[ 234 ][ 215 ],
   alphaCSR[ 234 ][ 216 ],
   alphaCSR[ 234 ][ 217 ],
   alphaCSR[ 234 ][ 218 ],
   alphaCSR[ 234 ][ 219 ],
   alphaCSR[ 234 ][ 220 ],
   alphaCSR[ 234 ][ 221 ],
   alphaCSR[ 234 ][ 222 ],
   alphaCSR[ 234 ][ 223 ],
   alphaCSR[ 234 ][ 224 ],
   alphaCSR[ 234 ][ 225 ],
   alphaCSR[ 234 ][ 226 ],
   alphaCSR[ 234 ][ 227 ],
   alphaCSR[ 234 ][ 228 ],
   alphaCSR[ 234 ][ 229 ],
   alphaCSR[ 234 ][ 230 ],
   alphaCSR[ 234 ][ 231 ],
   alphaCSR[ 234 ][ 232 ],
   alphaCSR[ 234 ][ 233 ],
   alphaCSR[ 234 ][ 234 ],
   alphaCSR[ 234 ][ 235 ],
   alphaCSR[ 234 ][ 236 ],
   alphaCSR[ 234 ][ 237 ],
   alphaCSR[ 234 ][ 238 ],
   alphaCSR[ 234 ][ 239 ],
   alphaCSR[ 234 ][ 240 ],
   alphaCSR[ 234 ][ 241 ],
   alphaCSR[ 234 ][ 242 ],
   alphaCSR[ 234 ][ 243 ],
   alphaCSR[ 234 ][ 244 ],
   alphaCSR[ 234 ][ 245 ],
   alphaCSR[ 234 ][ 246 ],
   alphaCSR[ 234 ][ 247 ],
   alphaCSR[ 234 ][ 248 ],
   alphaCSR[ 234 ][ 249 ],
   alphaCSR[ 234 ][ 250 ],
   alphaCSR[ 234 ][ 251 ],
   alphaCSR[ 234 ][ 252 ],
   alphaCSR[ 234 ][ 253 ],
   alphaCSR[ 234 ][ 254 ],
   alphaCSR[ 234 ][ 255 ],
   alphaCSR[ 234 ][ 256 ],
   alphaCSR[ 234 ][ 257 ],
   alphaCSR[ 234 ][ 258 ],
   alphaCSR[ 234 ][ 259 ],
   alphaCSR[ 234 ][ 260 ],
   alphaCSR[ 234 ][ 261 ],
   alphaCSR[ 234 ][ 262 ],
   alphaCSR[ 234 ][ 263 ],
   alphaCSR[ 234 ][ 264 ],
   alphaCSR[ 234 ][ 265 ],
   alphaCSR[ 234 ][ 266 ],
   alphaCSR[ 234 ][ 267 ],
   alphaCSR[ 234 ][ 268 ],
   alphaCSR[ 234 ][ 269 ],
   alphaCSR[ 234 ][ 270 ],
   alphaCSR[ 234 ][ 271 ],
   alphaCSR[ 234 ][ 272 ],
   alphaCSR[ 234 ][ 273 ],
   alphaCSR[ 234 ][ 274 ],
   alphaCSR[ 234 ][ 275 ],
   alphaCSR[ 234 ][ 276 ],
   alphaCSR[ 234 ][ 277 ],
   alphaCSR[ 234 ][ 278 ],
   alphaCSR[ 234 ][ 279 ],
   alphaCSR[ 234 ][ 280 ],
   alphaCSR[ 234 ][ 281 ],
   alphaCSR[ 234 ][ 282 ],
   alphaCSR[ 234 ][ 283 ],
   alphaCSR[ 234 ][ 284 ],
   alphaCSR[ 234 ][ 285 ],
   alphaCSR[ 234 ][ 286 ],
   alphaCSR[ 234 ][ 287 ],
   alphaCSR[ 234 ][ 288 ],
   alphaCSR[ 234 ][ 289 ],
   alphaCSR[ 234 ][ 290 ],
   alphaCSR[ 234 ][ 291 ],
   alphaCSR[ 234 ][ 292 ],
   alphaCSR[ 234 ][ 293 ],
   alphaCSR[ 234 ][ 294 ],
   alphaCSR[ 234 ][ 295 ],
   alphaCSR[ 234 ][ 296 ],
   alphaCSR[ 234 ][ 297 ],
   alphaCSR[ 234 ][ 298 ],
   alphaCSR[ 234 ][ 299 ],
   alphaCSR[ 234 ][ 300 ],
   alphaCSR[ 234 ][ 301 ],
   alphaCSR[ 234 ][ 302 ],
   alphaCSR[ 234 ][ 303 ],
   alphaCSR[ 234 ][ 304 ],
   alphaCSR[ 234 ][ 305 ],
   alphaCSR[ 234 ][ 306 ],
   alphaCSR[ 234 ][ 307 ],
   alphaCSR[ 234 ][ 308 ],
   alphaCSR[ 234 ][ 309 ],
   alphaCSR[ 234 ][ 310 ],
   alphaCSR[ 234 ][ 311 ],
   alphaCSR[ 234 ][ 312 ],
   alphaCSR[ 234 ][ 313 ],
   alphaCSR[ 234 ][ 314 ],
   alphaCSR[ 234 ][ 315 ],
   alphaCSR[ 234 ][ 316 ],
   alphaCSR[ 234 ][ 317 ],
   alphaCSR[ 234 ][ 318 ],
   alphaCSR[ 234 ][ 319 ],
   alphaCSR[ 234 ][ 320 ],
   alphaCSR[ 234 ][ 321 ],
   alphaCSR[ 234 ][ 322 ],
   alphaCSR[ 234 ][ 323 ],
   alphaCSR[ 234 ][ 324 ],
   alphaCSR[ 234 ][ 325 ],
   alphaCSR[ 234 ][ 326 ],
   alphaCSR[ 234 ][ 327 ],
   alphaCSR[ 234 ][ 328 ],
   alphaCSR[ 234 ][ 329 ],
   alphaCSR[ 234 ][ 330 ],
   alphaCSR[ 234 ][ 331 ],
   alphaCSR[ 234 ][ 332 ],
   alphaCSR[ 234 ][ 333 ],
   alphaCSR[ 234 ][ 334 ],
   alphaCSR[ 234 ][ 335 ],
   alphaCSR[ 234 ][ 336 ],
   alphaCSR[ 234 ][ 337 ],
   alphaCSR[ 234 ][ 338 ],
   alphaCSR[ 234 ][ 339 ],
   alphaCSR[ 234 ][ 340 ],
   alphaCSR[ 234 ][ 341 ],
   alphaCSR[ 234 ][ 342 ],
   alphaCSR[ 234 ][ 343 ],
   alphaCSR[ 234 ][ 344 ],
   alphaCSR[ 234 ][ 345 ],
   alphaCSR[ 234 ][ 346 ],
   alphaCSR[ 234 ][ 347 ],
   alphaCSR[ 234 ][ 348 ],
   alphaCSR[ 234 ][ 349 ],
   alphaCSR[ 234 ][ 350 ],
   alphaCSR[ 234 ][ 351 ],
   alphaCSR[ 234 ][ 352 ],
   alphaCSR[ 234 ][ 353 ],
   alphaCSR[ 234 ][ 354 ],
   alphaCSR[ 234 ][ 355 ],
   alphaCSR[ 234 ][ 356 ],
   alphaCSR[ 234 ][ 357 ],
   alphaCSR[ 234 ][ 358 ],
   alphaCSR[ 234 ][ 359 ],
   alphaCSR[ 234 ][ 360 ],
   alphaCSR[ 234 ][ 361 ],
   alphaCSR[ 234 ][ 362 ],
   alphaCSR[ 234 ][ 363 ],
   alphaCSR[ 234 ][ 364 ],
   alphaCSR[ 234 ][ 365 ],
   alphaCSR[ 234 ][ 366 ],
   alphaCSR[ 234 ][ 367 ],
   alphaCSR[ 234 ][ 368 ],
   alphaCSR[ 234 ][ 369 ],
   alphaCSR[ 234 ][ 370 ],
   alphaCSR[ 234 ][ 371 ],
   alphaCSR[ 234 ][ 372 ],
   alphaCSR[ 234 ][ 373 ],
   alphaCSR[ 234 ][ 374 ],
   alphaCSR[ 234 ][ 375 ],
   alphaCSR[ 234 ][ 376 ],
   alphaCSR[ 234 ][ 377 ],
   alphaCSR[ 234 ][ 378 ],
   alphaCSR[ 234 ][ 379 ],
   alphaCSR[ 234 ][ 380 ],
   alphaCSR[ 234 ][ 381 ],
   alphaCSR[ 234 ][ 382 ],
   alphaCSR[ 234 ][ 383 ],
   alphaCSR[ 235 ][ 0 ],
   alphaCSR[ 235 ][ 1 ],
   alphaCSR[ 235 ][ 2 ],
   alphaCSR[ 235 ][ 3 ],
   alphaCSR[ 235 ][ 4 ],
   alphaCSR[ 235 ][ 5 ],
   alphaCSR[ 235 ][ 6 ],
   alphaCSR[ 235 ][ 7 ],
   alphaCSR[ 235 ][ 8 ],
   alphaCSR[ 235 ][ 9 ],
   alphaCSR[ 235 ][ 10 ],
   alphaCSR[ 235 ][ 11 ],
   alphaCSR[ 235 ][ 12 ],
   alphaCSR[ 235 ][ 13 ],
   alphaCSR[ 235 ][ 14 ],
   alphaCSR[ 235 ][ 15 ],
   alphaCSR[ 235 ][ 16 ],
   alphaCSR[ 235 ][ 17 ],
   alphaCSR[ 235 ][ 18 ],
   alphaCSR[ 235 ][ 19 ],
   alphaCSR[ 235 ][ 20 ],
   alphaCSR[ 235 ][ 21 ],
   alphaCSR[ 235 ][ 22 ],
   alphaCSR[ 235 ][ 23 ],
   alphaCSR[ 235 ][ 24 ],
   alphaCSR[ 235 ][ 25 ],
   alphaCSR[ 235 ][ 26 ],
   alphaCSR[ 235 ][ 27 ],
   alphaCSR[ 235 ][ 28 ],
   alphaCSR[ 235 ][ 29 ],
   alphaCSR[ 235 ][ 30 ],
   alphaCSR[ 235 ][ 31 ],
   alphaCSR[ 235 ][ 32 ],
   alphaCSR[ 235 ][ 33 ],
   alphaCSR[ 235 ][ 34 ],
   alphaCSR[ 235 ][ 35 ],
   alphaCSR[ 235 ][ 36 ],
   alphaCSR[ 235 ][ 37 ],
   alphaCSR[ 235 ][ 38 ],
   alphaCSR[ 235 ][ 39 ],
   alphaCSR[ 235 ][ 40 ],
   alphaCSR[ 235 ][ 41 ],
   alphaCSR[ 235 ][ 42 ],
   alphaCSR[ 235 ][ 43 ],
   alphaCSR[ 235 ][ 44 ],
   alphaCSR[ 235 ][ 45 ],
   alphaCSR[ 235 ][ 46 ],
   alphaCSR[ 235 ][ 47 ],
   alphaCSR[ 235 ][ 48 ],
   alphaCSR[ 235 ][ 49 ],
   alphaCSR[ 235 ][ 50 ],
   alphaCSR[ 235 ][ 51 ],
   alphaCSR[ 235 ][ 52 ],
   alphaCSR[ 235 ][ 53 ],
   alphaCSR[ 235 ][ 54 ],
   alphaCSR[ 235 ][ 55 ],
   alphaCSR[ 235 ][ 56 ],
   alphaCSR[ 235 ][ 57 ],
   alphaCSR[ 235 ][ 58 ],
   alphaCSR[ 235 ][ 59 ],
   alphaCSR[ 235 ][ 60 ],
   alphaCSR[ 235 ][ 61 ],
   alphaCSR[ 235 ][ 62 ],
   alphaCSR[ 235 ][ 63 ],
   alphaCSR[ 235 ][ 64 ],
   alphaCSR[ 235 ][ 65 ],
   alphaCSR[ 235 ][ 66 ],
   alphaCSR[ 235 ][ 67 ],
   alphaCSR[ 235 ][ 68 ],
   alphaCSR[ 235 ][ 69 ],
   alphaCSR[ 235 ][ 70 ],
   alphaCSR[ 235 ][ 71 ],
   alphaCSR[ 235 ][ 72 ],
   alphaCSR[ 235 ][ 73 ],
   alphaCSR[ 235 ][ 74 ],
   alphaCSR[ 235 ][ 75 ],
   alphaCSR[ 235 ][ 76 ],
   alphaCSR[ 235 ][ 77 ],
   alphaCSR[ 235 ][ 78 ],
   alphaCSR[ 235 ][ 79 ],
   alphaCSR[ 235 ][ 80 ],
   alphaCSR[ 235 ][ 81 ],
   alphaCSR[ 235 ][ 82 ],
   alphaCSR[ 235 ][ 83 ],
   alphaCSR[ 235 ][ 84 ],
   alphaCSR[ 235 ][ 85 ],
   alphaCSR[ 235 ][ 86 ],
   alphaCSR[ 235 ][ 87 ],
   alphaCSR[ 235 ][ 88 ],
   alphaCSR[ 235 ][ 89 ],
   alphaCSR[ 235 ][ 90 ],
   alphaCSR[ 235 ][ 91 ],
   alphaCSR[ 235 ][ 92 ],
   alphaCSR[ 235 ][ 93 ],
   alphaCSR[ 235 ][ 94 ],
   alphaCSR[ 235 ][ 95 ],
   alphaCSR[ 235 ][ 96 ],
   alphaCSR[ 235 ][ 97 ],
   alphaCSR[ 235 ][ 98 ],
   alphaCSR[ 235 ][ 99 ],
   alphaCSR[ 235 ][ 100 ],
   alphaCSR[ 235 ][ 101 ],
   alphaCSR[ 235 ][ 102 ],
   alphaCSR[ 235 ][ 103 ],
   alphaCSR[ 235 ][ 104 ],
   alphaCSR[ 235 ][ 105 ],
   alphaCSR[ 235 ][ 106 ],
   alphaCSR[ 235 ][ 107 ],
   alphaCSR[ 235 ][ 108 ],
   alphaCSR[ 235 ][ 109 ],
   alphaCSR[ 235 ][ 110 ],
   alphaCSR[ 235 ][ 111 ],
   alphaCSR[ 235 ][ 112 ],
   alphaCSR[ 235 ][ 113 ],
   alphaCSR[ 235 ][ 114 ],
   alphaCSR[ 235 ][ 115 ],
   alphaCSR[ 235 ][ 116 ],
   alphaCSR[ 235 ][ 117 ],
   alphaCSR[ 235 ][ 118 ],
   alphaCSR[ 235 ][ 119 ],
   alphaCSR[ 235 ][ 120 ],
   alphaCSR[ 235 ][ 121 ],
   alphaCSR[ 235 ][ 122 ],
   alphaCSR[ 235 ][ 123 ],
   alphaCSR[ 235 ][ 124 ],
   alphaCSR[ 235 ][ 125 ],
   alphaCSR[ 235 ][ 126 ],
   alphaCSR[ 235 ][ 127 ],
   alphaCSR[ 235 ][ 128 ],
   alphaCSR[ 235 ][ 129 ],
   alphaCSR[ 235 ][ 130 ],
   alphaCSR[ 235 ][ 131 ],
   alphaCSR[ 235 ][ 132 ],
   alphaCSR[ 235 ][ 133 ],
   alphaCSR[ 235 ][ 134 ],
   alphaCSR[ 235 ][ 135 ],
   alphaCSR[ 235 ][ 136 ],
   alphaCSR[ 235 ][ 137 ],
   alphaCSR[ 235 ][ 138 ],
   alphaCSR[ 235 ][ 139 ],
   alphaCSR[ 235 ][ 140 ],
   alphaCSR[ 235 ][ 141 ],
   alphaCSR[ 235 ][ 142 ],
   alphaCSR[ 235 ][ 143 ],
   alphaCSR[ 235 ][ 144 ],
   alphaCSR[ 235 ][ 145 ],
   alphaCSR[ 235 ][ 146 ],
   alphaCSR[ 235 ][ 147 ],
   alphaCSR[ 235 ][ 148 ],
   alphaCSR[ 235 ][ 149 ],
   alphaCSR[ 235 ][ 150 ],
   alphaCSR[ 235 ][ 151 ],
   alphaCSR[ 235 ][ 152 ],
   alphaCSR[ 235 ][ 153 ],
   alphaCSR[ 235 ][ 154 ],
   alphaCSR[ 235 ][ 155 ],
   alphaCSR[ 235 ][ 156 ],
   alphaCSR[ 235 ][ 157 ],
   alphaCSR[ 235 ][ 158 ],
   alphaCSR[ 235 ][ 159 ],
   alphaCSR[ 235 ][ 160 ],
   alphaCSR[ 235 ][ 161 ],
   alphaCSR[ 235 ][ 162 ],
   alphaCSR[ 235 ][ 163 ],
   alphaCSR[ 235 ][ 164 ],
   alphaCSR[ 235 ][ 165 ],
   alphaCSR[ 235 ][ 166 ],
   alphaCSR[ 235 ][ 167 ],
   alphaCSR[ 235 ][ 168 ],
   alphaCSR[ 235 ][ 169 ],
   alphaCSR[ 235 ][ 170 ],
   alphaCSR[ 235 ][ 171 ],
   alphaCSR[ 235 ][ 172 ],
   alphaCSR[ 235 ][ 173 ],
   alphaCSR[ 235 ][ 174 ],
   alphaCSR[ 235 ][ 175 ],
   alphaCSR[ 235 ][ 176 ],
   alphaCSR[ 235 ][ 177 ],
   alphaCSR[ 235 ][ 178 ],
   alphaCSR[ 235 ][ 179 ],
   alphaCSR[ 235 ][ 180 ],
   alphaCSR[ 235 ][ 181 ],
   alphaCSR[ 235 ][ 182 ],
   alphaCSR[ 235 ][ 183 ],
   alphaCSR[ 235 ][ 184 ],
   alphaCSR[ 235 ][ 185 ],
   alphaCSR[ 235 ][ 186 ],
   alphaCSR[ 235 ][ 187 ],
   alphaCSR[ 235 ][ 188 ],
   alphaCSR[ 235 ][ 189 ],
   alphaCSR[ 235 ][ 190 ],
   alphaCSR[ 235 ][ 191 ],
   alphaCSR[ 235 ][ 192 ],
   alphaCSR[ 235 ][ 193 ],
   alphaCSR[ 235 ][ 194 ],
   alphaCSR[ 235 ][ 195 ],
   alphaCSR[ 235 ][ 196 ],
   alphaCSR[ 235 ][ 197 ],
   alphaCSR[ 235 ][ 198 ],
   alphaCSR[ 235 ][ 199 ],
   alphaCSR[ 235 ][ 200 ],
   alphaCSR[ 235 ][ 201 ],
   alphaCSR[ 235 ][ 202 ],
   alphaCSR[ 235 ][ 203 ],
   alphaCSR[ 235 ][ 204 ],
   alphaCSR[ 235 ][ 205 ],
   alphaCSR[ 235 ][ 206 ],
   alphaCSR[ 235 ][ 207 ],
   alphaCSR[ 235 ][ 208 ],
   alphaCSR[ 235 ][ 209 ],
   alphaCSR[ 235 ][ 210 ],
   alphaCSR[ 235 ][ 211 ],
   alphaCSR[ 235 ][ 212 ],
   alphaCSR[ 235 ][ 213 ],
   alphaCSR[ 235 ][ 214 ],
   alphaCSR[ 235 ][ 215 ],
   alphaCSR[ 235 ][ 216 ],
   alphaCSR[ 235 ][ 217 ],
   alphaCSR[ 235 ][ 218 ],
   alphaCSR[ 235 ][ 219 ],
   alphaCSR[ 235 ][ 220 ],
   alphaCSR[ 235 ][ 221 ],
   alphaCSR[ 235 ][ 222 ],
   alphaCSR[ 235 ][ 223 ],
   alphaCSR[ 235 ][ 224 ],
   alphaCSR[ 235 ][ 225 ],
   alphaCSR[ 235 ][ 226 ],
   alphaCSR[ 235 ][ 227 ],
   alphaCSR[ 235 ][ 228 ],
   alphaCSR[ 235 ][ 229 ],
   alphaCSR[ 235 ][ 230 ],
   alphaCSR[ 235 ][ 231 ],
   alphaCSR[ 235 ][ 232 ],
   alphaCSR[ 235 ][ 233 ],
   alphaCSR[ 235 ][ 234 ],
   alphaCSR[ 235 ][ 235 ],
   alphaCSR[ 235 ][ 236 ],
   alphaCSR[ 235 ][ 237 ],
   alphaCSR[ 235 ][ 238 ],
   alphaCSR[ 235 ][ 239 ],
   alphaCSR[ 235 ][ 240 ],
   alphaCSR[ 235 ][ 241 ],
   alphaCSR[ 235 ][ 242 ],
   alphaCSR[ 235 ][ 243 ],
   alphaCSR[ 235 ][ 244 ],
   alphaCSR[ 235 ][ 245 ],
   alphaCSR[ 235 ][ 246 ],
   alphaCSR[ 235 ][ 247 ],
   alphaCSR[ 235 ][ 248 ],
   alphaCSR[ 235 ][ 249 ],
   alphaCSR[ 235 ][ 250 ],
   alphaCSR[ 235 ][ 251 ],
   alphaCSR[ 235 ][ 252 ],
   alphaCSR[ 235 ][ 253 ],
   alphaCSR[ 235 ][ 254 ],
   alphaCSR[ 235 ][ 255 ],
   alphaCSR[ 235 ][ 256 ],
   alphaCSR[ 235 ][ 257 ],
   alphaCSR[ 235 ][ 258 ],
   alphaCSR[ 235 ][ 259 ],
   alphaCSR[ 235 ][ 260 ],
   alphaCSR[ 235 ][ 261 ],
   alphaCSR[ 235 ][ 262 ],
   alphaCSR[ 235 ][ 263 ],
   alphaCSR[ 235 ][ 264 ],
   alphaCSR[ 235 ][ 265 ],
   alphaCSR[ 235 ][ 266 ],
   alphaCSR[ 235 ][ 267 ],
   alphaCSR[ 235 ][ 268 ],
   alphaCSR[ 235 ][ 269 ],
   alphaCSR[ 235 ][ 270 ],
   alphaCSR[ 235 ][ 271 ],
   alphaCSR[ 235 ][ 272 ],
   alphaCSR[ 235 ][ 273 ],
   alphaCSR[ 235 ][ 274 ],
   alphaCSR[ 235 ][ 275 ],
   alphaCSR[ 235 ][ 276 ],
   alphaCSR[ 235 ][ 277 ],
   alphaCSR[ 235 ][ 278 ],
   alphaCSR[ 235 ][ 279 ],
   alphaCSR[ 235 ][ 280 ],
   alphaCSR[ 235 ][ 281 ],
   alphaCSR[ 235 ][ 282 ],
   alphaCSR[ 235 ][ 283 ],
   alphaCSR[ 235 ][ 284 ],
   alphaCSR[ 235 ][ 285 ],
   alphaCSR[ 235 ][ 286 ],
   alphaCSR[ 235 ][ 287 ],
   alphaCSR[ 235 ][ 288 ],
   alphaCSR[ 235 ][ 289 ],
   alphaCSR[ 235 ][ 290 ],
   alphaCSR[ 235 ][ 291 ],
   alphaCSR[ 235 ][ 292 ],
   alphaCSR[ 235 ][ 293 ],
   alphaCSR[ 235 ][ 294 ],
   alphaCSR[ 235 ][ 295 ],
   alphaCSR[ 235 ][ 296 ],
   alphaCSR[ 235 ][ 297 ],
   alphaCSR[ 235 ][ 298 ],
   alphaCSR[ 235 ][ 299 ],
   alphaCSR[ 235 ][ 300 ],
   alphaCSR[ 235 ][ 301 ],
   alphaCSR[ 235 ][ 302 ],
   alphaCSR[ 235 ][ 303 ],
   alphaCSR[ 235 ][ 304 ],
   alphaCSR[ 235 ][ 305 ],
   alphaCSR[ 235 ][ 306 ],
   alphaCSR[ 235 ][ 307 ],
   alphaCSR[ 235 ][ 308 ],
   alphaCSR[ 235 ][ 309 ],
   alphaCSR[ 235 ][ 310 ],
   alphaCSR[ 235 ][ 311 ],
   alphaCSR[ 235 ][ 312 ],
   alphaCSR[ 235 ][ 313 ],
   alphaCSR[ 235 ][ 314 ],
   alphaCSR[ 235 ][ 315 ],
   alphaCSR[ 235 ][ 316 ],
   alphaCSR[ 235 ][ 317 ],
   alphaCSR[ 235 ][ 318 ],
   alphaCSR[ 235 ][ 319 ],
   alphaCSR[ 235 ][ 320 ],
   alphaCSR[ 235 ][ 321 ],
   alphaCSR[ 235 ][ 322 ],
   alphaCSR[ 235 ][ 323 ],
   alphaCSR[ 235 ][ 324 ],
   alphaCSR[ 235 ][ 325 ],
   alphaCSR[ 235 ][ 326 ],
   alphaCSR[ 235 ][ 327 ],
   alphaCSR[ 235 ][ 328 ],
   alphaCSR[ 235 ][ 329 ],
   alphaCSR[ 235 ][ 330 ],
   alphaCSR[ 235 ][ 331 ],
   alphaCSR[ 235 ][ 332 ],
   alphaCSR[ 235 ][ 333 ],
   alphaCSR[ 235 ][ 334 ],
   alphaCSR[ 235 ][ 335 ],
   alphaCSR[ 235 ][ 336 ],
   alphaCSR[ 235 ][ 337 ],
   alphaCSR[ 235 ][ 338 ],
   alphaCSR[ 235 ][ 339 ],
   alphaCSR[ 235 ][ 340 ],
   alphaCSR[ 235 ][ 341 ],
   alphaCSR[ 235 ][ 342 ],
   alphaCSR[ 235 ][ 343 ],
   alphaCSR[ 235 ][ 344 ],
   alphaCSR[ 235 ][ 345 ],
   alphaCSR[ 235 ][ 346 ],
   alphaCSR[ 235 ][ 347 ],
   alphaCSR[ 235 ][ 348 ],
   alphaCSR[ 235 ][ 349 ],
   alphaCSR[ 235 ][ 350 ],
   alphaCSR[ 235 ][ 351 ],
   alphaCSR[ 235 ][ 352 ],
   alphaCSR[ 235 ][ 353 ],
   alphaCSR[ 235 ][ 354 ],
   alphaCSR[ 235 ][ 355 ],
   alphaCSR[ 235 ][ 356 ],
   alphaCSR[ 235 ][ 357 ],
   alphaCSR[ 235 ][ 358 ],
   alphaCSR[ 235 ][ 359 ],
   alphaCSR[ 235 ][ 360 ],
   alphaCSR[ 235 ][ 361 ],
   alphaCSR[ 235 ][ 362 ],
   alphaCSR[ 235 ][ 363 ],
   alphaCSR[ 235 ][ 364 ],
   alphaCSR[ 235 ][ 365 ],
   alphaCSR[ 235 ][ 366 ],
   alphaCSR[ 235 ][ 367 ],
   alphaCSR[ 235 ][ 368 ],
   alphaCSR[ 235 ][ 369 ],
   alphaCSR[ 235 ][ 370 ],
   alphaCSR[ 235 ][ 371 ],
   alphaCSR[ 235 ][ 372 ],
   alphaCSR[ 235 ][ 373 ],
   alphaCSR[ 235 ][ 374 ],
   alphaCSR[ 235 ][ 375 ],
   alphaCSR[ 235 ][ 376 ],
   alphaCSR[ 235 ][ 377 ],
   alphaCSR[ 235 ][ 378 ],
   alphaCSR[ 235 ][ 379 ],
   alphaCSR[ 235 ][ 380 ],
   alphaCSR[ 235 ][ 381 ],
   alphaCSR[ 235 ][ 382 ],
   alphaCSR[ 235 ][ 383 ],
   alphaCSR[ 236 ][ 0 ],
   alphaCSR[ 236 ][ 1 ],
   alphaCSR[ 236 ][ 2 ],
   alphaCSR[ 236 ][ 3 ],
   alphaCSR[ 236 ][ 4 ],
   alphaCSR[ 236 ][ 5 ],
   alphaCSR[ 236 ][ 6 ],
   alphaCSR[ 236 ][ 7 ],
   alphaCSR[ 236 ][ 8 ],
   alphaCSR[ 236 ][ 9 ],
   alphaCSR[ 236 ][ 10 ],
   alphaCSR[ 236 ][ 11 ],
   alphaCSR[ 236 ][ 12 ],
   alphaCSR[ 236 ][ 13 ],
   alphaCSR[ 236 ][ 14 ],
   alphaCSR[ 236 ][ 15 ],
   alphaCSR[ 236 ][ 16 ],
   alphaCSR[ 236 ][ 17 ],
   alphaCSR[ 236 ][ 18 ],
   alphaCSR[ 236 ][ 19 ],
   alphaCSR[ 236 ][ 20 ],
   alphaCSR[ 236 ][ 21 ],
   alphaCSR[ 236 ][ 22 ],
   alphaCSR[ 236 ][ 23 ],
   alphaCSR[ 236 ][ 24 ],
   alphaCSR[ 236 ][ 25 ],
   alphaCSR[ 236 ][ 26 ],
   alphaCSR[ 236 ][ 27 ],
   alphaCSR[ 236 ][ 28 ],
   alphaCSR[ 236 ][ 29 ],
   alphaCSR[ 236 ][ 30 ],
   alphaCSR[ 236 ][ 31 ],
   alphaCSR[ 236 ][ 32 ],
   alphaCSR[ 236 ][ 33 ],
   alphaCSR[ 236 ][ 34 ],
   alphaCSR[ 236 ][ 35 ],
   alphaCSR[ 236 ][ 36 ],
   alphaCSR[ 236 ][ 37 ],
   alphaCSR[ 236 ][ 38 ],
   alphaCSR[ 236 ][ 39 ],
   alphaCSR[ 236 ][ 40 ],
   alphaCSR[ 236 ][ 41 ],
   alphaCSR[ 236 ][ 42 ],
   alphaCSR[ 236 ][ 43 ],
   alphaCSR[ 236 ][ 44 ],
   alphaCSR[ 236 ][ 45 ],
   alphaCSR[ 236 ][ 46 ],
   alphaCSR[ 236 ][ 47 ],
   alphaCSR[ 236 ][ 48 ],
   alphaCSR[ 236 ][ 49 ],
   alphaCSR[ 236 ][ 50 ],
   alphaCSR[ 236 ][ 51 ],
   alphaCSR[ 236 ][ 52 ],
   alphaCSR[ 236 ][ 53 ],
   alphaCSR[ 236 ][ 54 ],
   alphaCSR[ 236 ][ 55 ],
   alphaCSR[ 236 ][ 56 ],
   alphaCSR[ 236 ][ 57 ],
   alphaCSR[ 236 ][ 58 ],
   alphaCSR[ 236 ][ 59 ],
   alphaCSR[ 236 ][ 60 ],
   alphaCSR[ 236 ][ 61 ],
   alphaCSR[ 236 ][ 62 ],
   alphaCSR[ 236 ][ 63 ],
   alphaCSR[ 236 ][ 64 ],
   alphaCSR[ 236 ][ 65 ],
   alphaCSR[ 236 ][ 66 ],
   alphaCSR[ 236 ][ 67 ],
   alphaCSR[ 236 ][ 68 ],
   alphaCSR[ 236 ][ 69 ],
   alphaCSR[ 236 ][ 70 ],
   alphaCSR[ 236 ][ 71 ],
   alphaCSR[ 236 ][ 72 ],
   alphaCSR[ 236 ][ 73 ],
   alphaCSR[ 236 ][ 74 ],
   alphaCSR[ 236 ][ 75 ],
   alphaCSR[ 236 ][ 76 ],
   alphaCSR[ 236 ][ 77 ],
   alphaCSR[ 236 ][ 78 ],
   alphaCSR[ 236 ][ 79 ],
   alphaCSR[ 236 ][ 80 ],
   alphaCSR[ 236 ][ 81 ],
   alphaCSR[ 236 ][ 82 ],
   alphaCSR[ 236 ][ 83 ],
   alphaCSR[ 236 ][ 84 ],
   alphaCSR[ 236 ][ 85 ],
   alphaCSR[ 236 ][ 86 ],
   alphaCSR[ 236 ][ 87 ],
   alphaCSR[ 236 ][ 88 ],
   alphaCSR[ 236 ][ 89 ],
   alphaCSR[ 236 ][ 90 ],
   alphaCSR[ 236 ][ 91 ],
   alphaCSR[ 236 ][ 92 ],
   alphaCSR[ 236 ][ 93 ],
   alphaCSR[ 236 ][ 94 ],
   alphaCSR[ 236 ][ 95 ],
   alphaCSR[ 236 ][ 96 ],
   alphaCSR[ 236 ][ 97 ],
   alphaCSR[ 236 ][ 98 ],
   alphaCSR[ 236 ][ 99 ],
   alphaCSR[ 236 ][ 100 ],
   alphaCSR[ 236 ][ 101 ],
   alphaCSR[ 236 ][ 102 ],
   alphaCSR[ 236 ][ 103 ],
   alphaCSR[ 236 ][ 104 ],
   alphaCSR[ 236 ][ 105 ],
   alphaCSR[ 236 ][ 106 ],
   alphaCSR[ 236 ][ 107 ],
   alphaCSR[ 236 ][ 108 ],
   alphaCSR[ 236 ][ 109 ],
   alphaCSR[ 236 ][ 110 ],
   alphaCSR[ 236 ][ 111 ],
   alphaCSR[ 236 ][ 112 ],
   alphaCSR[ 236 ][ 113 ],
   alphaCSR[ 236 ][ 114 ],
   alphaCSR[ 236 ][ 115 ],
   alphaCSR[ 236 ][ 116 ],
   alphaCSR[ 236 ][ 117 ],
   alphaCSR[ 236 ][ 118 ],
   alphaCSR[ 236 ][ 119 ],
   alphaCSR[ 236 ][ 120 ],
   alphaCSR[ 236 ][ 121 ],
   alphaCSR[ 236 ][ 122 ],
   alphaCSR[ 236 ][ 123 ],
   alphaCSR[ 236 ][ 124 ],
   alphaCSR[ 236 ][ 125 ],
   alphaCSR[ 236 ][ 126 ],
   alphaCSR[ 236 ][ 127 ],
   alphaCSR[ 236 ][ 128 ],
   alphaCSR[ 236 ][ 129 ],
   alphaCSR[ 236 ][ 130 ],
   alphaCSR[ 236 ][ 131 ],
   alphaCSR[ 236 ][ 132 ],
   alphaCSR[ 236 ][ 133 ],
   alphaCSR[ 236 ][ 134 ],
   alphaCSR[ 236 ][ 135 ],
   alphaCSR[ 236 ][ 136 ],
   alphaCSR[ 236 ][ 137 ],
   alphaCSR[ 236 ][ 138 ],
   alphaCSR[ 236 ][ 139 ],
   alphaCSR[ 236 ][ 140 ],
   alphaCSR[ 236 ][ 141 ],
   alphaCSR[ 236 ][ 142 ],
   alphaCSR[ 236 ][ 143 ],
   alphaCSR[ 236 ][ 144 ],
   alphaCSR[ 236 ][ 145 ],
   alphaCSR[ 236 ][ 146 ],
   alphaCSR[ 236 ][ 147 ],
   alphaCSR[ 236 ][ 148 ],
   alphaCSR[ 236 ][ 149 ],
   alphaCSR[ 236 ][ 150 ],
   alphaCSR[ 236 ][ 151 ],
   alphaCSR[ 236 ][ 152 ],
   alphaCSR[ 236 ][ 153 ],
   alphaCSR[ 236 ][ 154 ],
   alphaCSR[ 236 ][ 155 ],
   alphaCSR[ 236 ][ 156 ],
   alphaCSR[ 236 ][ 157 ],
   alphaCSR[ 236 ][ 158 ],
   alphaCSR[ 236 ][ 159 ],
   alphaCSR[ 236 ][ 160 ],
   alphaCSR[ 236 ][ 161 ],
   alphaCSR[ 236 ][ 162 ],
   alphaCSR[ 236 ][ 163 ],
   alphaCSR[ 236 ][ 164 ],
   alphaCSR[ 236 ][ 165 ],
   alphaCSR[ 236 ][ 166 ],
   alphaCSR[ 236 ][ 167 ],
   alphaCSR[ 236 ][ 168 ],
   alphaCSR[ 236 ][ 169 ],
   alphaCSR[ 236 ][ 170 ],
   alphaCSR[ 236 ][ 171 ],
   alphaCSR[ 236 ][ 172 ],
   alphaCSR[ 236 ][ 173 ],
   alphaCSR[ 236 ][ 174 ],
   alphaCSR[ 236 ][ 175 ],
   alphaCSR[ 236 ][ 176 ],
   alphaCSR[ 236 ][ 177 ],
   alphaCSR[ 236 ][ 178 ],
   alphaCSR[ 236 ][ 179 ],
   alphaCSR[ 236 ][ 180 ],
   alphaCSR[ 236 ][ 181 ],
   alphaCSR[ 236 ][ 182 ],
   alphaCSR[ 236 ][ 183 ],
   alphaCSR[ 236 ][ 184 ],
   alphaCSR[ 236 ][ 185 ],
   alphaCSR[ 236 ][ 186 ],
   alphaCSR[ 236 ][ 187 ],
   alphaCSR[ 236 ][ 188 ],
   alphaCSR[ 236 ][ 189 ],
   alphaCSR[ 236 ][ 190 ],
   alphaCSR[ 236 ][ 191 ],
   alphaCSR[ 236 ][ 192 ],
   alphaCSR[ 236 ][ 193 ],
   alphaCSR[ 236 ][ 194 ],
   alphaCSR[ 236 ][ 195 ],
   alphaCSR[ 236 ][ 196 ],
   alphaCSR[ 236 ][ 197 ],
   alphaCSR[ 236 ][ 198 ],
   alphaCSR[ 236 ][ 199 ],
   alphaCSR[ 236 ][ 200 ],
   alphaCSR[ 236 ][ 201 ],
   alphaCSR[ 236 ][ 202 ],
   alphaCSR[ 236 ][ 203 ],
   alphaCSR[ 236 ][ 204 ],
   alphaCSR[ 236 ][ 205 ],
   alphaCSR[ 236 ][ 206 ],
   alphaCSR[ 236 ][ 207 ],
   alphaCSR[ 236 ][ 208 ],
   alphaCSR[ 236 ][ 209 ],
   alphaCSR[ 236 ][ 210 ],
   alphaCSR[ 236 ][ 211 ],
   alphaCSR[ 236 ][ 212 ],
   alphaCSR[ 236 ][ 213 ],
   alphaCSR[ 236 ][ 214 ],
   alphaCSR[ 236 ][ 215 ],
   alphaCSR[ 236 ][ 216 ],
   alphaCSR[ 236 ][ 217 ],
   alphaCSR[ 236 ][ 218 ],
   alphaCSR[ 236 ][ 219 ],
   alphaCSR[ 236 ][ 220 ],
   alphaCSR[ 236 ][ 221 ],
   alphaCSR[ 236 ][ 222 ],
   alphaCSR[ 236 ][ 223 ],
   alphaCSR[ 236 ][ 224 ],
   alphaCSR[ 236 ][ 225 ],
   alphaCSR[ 236 ][ 226 ],
   alphaCSR[ 236 ][ 227 ],
   alphaCSR[ 236 ][ 228 ],
   alphaCSR[ 236 ][ 229 ],
   alphaCSR[ 236 ][ 230 ],
   alphaCSR[ 236 ][ 231 ],
   alphaCSR[ 236 ][ 232 ],
   alphaCSR[ 236 ][ 233 ],
   alphaCSR[ 236 ][ 234 ],
   alphaCSR[ 236 ][ 235 ],
   alphaCSR[ 236 ][ 236 ],
   alphaCSR[ 236 ][ 237 ],
   alphaCSR[ 236 ][ 238 ],
   alphaCSR[ 236 ][ 239 ],
   alphaCSR[ 236 ][ 240 ],
   alphaCSR[ 236 ][ 241 ],
   alphaCSR[ 236 ][ 242 ],
   alphaCSR[ 236 ][ 243 ],
   alphaCSR[ 236 ][ 244 ],
   alphaCSR[ 236 ][ 245 ],
   alphaCSR[ 236 ][ 246 ],
   alphaCSR[ 236 ][ 247 ],
   alphaCSR[ 236 ][ 248 ],
   alphaCSR[ 236 ][ 249 ],
   alphaCSR[ 236 ][ 250 ],
   alphaCSR[ 236 ][ 251 ],
   alphaCSR[ 236 ][ 252 ],
   alphaCSR[ 236 ][ 253 ],
   alphaCSR[ 236 ][ 254 ],
   alphaCSR[ 236 ][ 255 ],
   alphaCSR[ 236 ][ 256 ],
   alphaCSR[ 236 ][ 257 ],
   alphaCSR[ 236 ][ 258 ],
   alphaCSR[ 236 ][ 259 ],
   alphaCSR[ 236 ][ 260 ],
   alphaCSR[ 236 ][ 261 ],
   alphaCSR[ 236 ][ 262 ],
   alphaCSR[ 236 ][ 263 ],
   alphaCSR[ 236 ][ 264 ],
   alphaCSR[ 236 ][ 265 ],
   alphaCSR[ 236 ][ 266 ],
   alphaCSR[ 236 ][ 267 ],
   alphaCSR[ 236 ][ 268 ],
   alphaCSR[ 236 ][ 269 ],
   alphaCSR[ 236 ][ 270 ],
   alphaCSR[ 236 ][ 271 ],
   alphaCSR[ 236 ][ 272 ],
   alphaCSR[ 236 ][ 273 ],
   alphaCSR[ 236 ][ 274 ],
   alphaCSR[ 236 ][ 275 ],
   alphaCSR[ 236 ][ 276 ],
   alphaCSR[ 236 ][ 277 ],
   alphaCSR[ 236 ][ 278 ],
   alphaCSR[ 236 ][ 279 ],
   alphaCSR[ 236 ][ 280 ],
   alphaCSR[ 236 ][ 281 ],
   alphaCSR[ 236 ][ 282 ],
   alphaCSR[ 236 ][ 283 ],
   alphaCSR[ 236 ][ 284 ],
   alphaCSR[ 236 ][ 285 ],
   alphaCSR[ 236 ][ 286 ],
   alphaCSR[ 236 ][ 287 ],
   alphaCSR[ 236 ][ 288 ],
   alphaCSR[ 236 ][ 289 ],
   alphaCSR[ 236 ][ 290 ],
   alphaCSR[ 236 ][ 291 ],
   alphaCSR[ 236 ][ 292 ],
   alphaCSR[ 236 ][ 293 ],
   alphaCSR[ 236 ][ 294 ],
   alphaCSR[ 236 ][ 295 ],
   alphaCSR[ 236 ][ 296 ],
   alphaCSR[ 236 ][ 297 ],
   alphaCSR[ 236 ][ 298 ],
   alphaCSR[ 236 ][ 299 ],
   alphaCSR[ 236 ][ 300 ],
   alphaCSR[ 236 ][ 301 ],
   alphaCSR[ 236 ][ 302 ],
   alphaCSR[ 236 ][ 303 ],
   alphaCSR[ 236 ][ 304 ],
   alphaCSR[ 236 ][ 305 ],
   alphaCSR[ 236 ][ 306 ],
   alphaCSR[ 236 ][ 307 ],
   alphaCSR[ 236 ][ 308 ],
   alphaCSR[ 236 ][ 309 ],
   alphaCSR[ 236 ][ 310 ],
   alphaCSR[ 236 ][ 311 ],
   alphaCSR[ 236 ][ 312 ],
   alphaCSR[ 236 ][ 313 ],
   alphaCSR[ 236 ][ 314 ],
   alphaCSR[ 236 ][ 315 ],
   alphaCSR[ 236 ][ 316 ],
   alphaCSR[ 236 ][ 317 ],
   alphaCSR[ 236 ][ 318 ],
   alphaCSR[ 236 ][ 319 ],
   alphaCSR[ 236 ][ 320 ],
   alphaCSR[ 236 ][ 321 ],
   alphaCSR[ 236 ][ 322 ],
   alphaCSR[ 236 ][ 323 ],
   alphaCSR[ 236 ][ 324 ],
   alphaCSR[ 236 ][ 325 ],
   alphaCSR[ 236 ][ 326 ],
   alphaCSR[ 236 ][ 327 ],
   alphaCSR[ 236 ][ 328 ],
   alphaCSR[ 236 ][ 329 ],
   alphaCSR[ 236 ][ 330 ],
   alphaCSR[ 236 ][ 331 ],
   alphaCSR[ 236 ][ 332 ],
   alphaCSR[ 236 ][ 333 ],
   alphaCSR[ 236 ][ 334 ],
   alphaCSR[ 236 ][ 335 ],
   alphaCSR[ 236 ][ 336 ],
   alphaCSR[ 236 ][ 337 ],
   alphaCSR[ 236 ][ 338 ],
   alphaCSR[ 236 ][ 339 ],
   alphaCSR[ 236 ][ 340 ],
   alphaCSR[ 236 ][ 341 ],
   alphaCSR[ 236 ][ 342 ],
   alphaCSR[ 236 ][ 343 ],
   alphaCSR[ 236 ][ 344 ],
   alphaCSR[ 236 ][ 345 ],
   alphaCSR[ 236 ][ 346 ],
   alphaCSR[ 236 ][ 347 ],
   alphaCSR[ 236 ][ 348 ],
   alphaCSR[ 236 ][ 349 ],
   alphaCSR[ 236 ][ 350 ],
   alphaCSR[ 236 ][ 351 ],
   alphaCSR[ 236 ][ 352 ],
   alphaCSR[ 236 ][ 353 ],
   alphaCSR[ 236 ][ 354 ],
   alphaCSR[ 236 ][ 355 ],
   alphaCSR[ 236 ][ 356 ],
   alphaCSR[ 236 ][ 357 ],
   alphaCSR[ 236 ][ 358 ],
   alphaCSR[ 236 ][ 359 ],
   alphaCSR[ 236 ][ 360 ],
   alphaCSR[ 236 ][ 361 ],
   alphaCSR[ 236 ][ 362 ],
   alphaCSR[ 236 ][ 363 ],
   alphaCSR[ 236 ][ 364 ],
   alphaCSR[ 236 ][ 365 ],
   alphaCSR[ 236 ][ 366 ],
   alphaCSR[ 236 ][ 367 ],
   alphaCSR[ 236 ][ 368 ],
   alphaCSR[ 236 ][ 369 ],
   alphaCSR[ 236 ][ 370 ],
   alphaCSR[ 236 ][ 371 ],
   alphaCSR[ 236 ][ 372 ],
   alphaCSR[ 236 ][ 373 ],
   alphaCSR[ 236 ][ 374 ],
   alphaCSR[ 236 ][ 375 ],
   alphaCSR[ 236 ][ 376 ],
   alphaCSR[ 236 ][ 377 ],
   alphaCSR[ 236 ][ 378 ],
   alphaCSR[ 236 ][ 379 ],
   alphaCSR[ 236 ][ 380 ],
   alphaCSR[ 236 ][ 381 ],
   alphaCSR[ 236 ][ 382 ],
   alphaCSR[ 236 ][ 383 ],
   alphaCSR[ 237 ][ 0 ],
   alphaCSR[ 237 ][ 1 ],
   alphaCSR[ 237 ][ 2 ],
   alphaCSR[ 237 ][ 3 ],
   alphaCSR[ 237 ][ 4 ],
   alphaCSR[ 237 ][ 5 ],
   alphaCSR[ 237 ][ 6 ],
   alphaCSR[ 237 ][ 7 ],
   alphaCSR[ 237 ][ 8 ],
   alphaCSR[ 237 ][ 9 ],
   alphaCSR[ 237 ][ 10 ],
   alphaCSR[ 237 ][ 11 ],
   alphaCSR[ 237 ][ 12 ],
   alphaCSR[ 237 ][ 13 ],
   alphaCSR[ 237 ][ 14 ],
   alphaCSR[ 237 ][ 15 ],
   alphaCSR[ 237 ][ 16 ],
   alphaCSR[ 237 ][ 17 ],
   alphaCSR[ 237 ][ 18 ],
   alphaCSR[ 237 ][ 19 ],
   alphaCSR[ 237 ][ 20 ],
   alphaCSR[ 237 ][ 21 ],
   alphaCSR[ 237 ][ 22 ],
   alphaCSR[ 237 ][ 23 ],
   alphaCSR[ 237 ][ 24 ],
   alphaCSR[ 237 ][ 25 ],
   alphaCSR[ 237 ][ 26 ],
   alphaCSR[ 237 ][ 27 ],
   alphaCSR[ 237 ][ 28 ],
   alphaCSR[ 237 ][ 29 ],
   alphaCSR[ 237 ][ 30 ],
   alphaCSR[ 237 ][ 31 ],
   alphaCSR[ 237 ][ 32 ],
   alphaCSR[ 237 ][ 33 ],
   alphaCSR[ 237 ][ 34 ],
   alphaCSR[ 237 ][ 35 ],
   alphaCSR[ 237 ][ 36 ],
   alphaCSR[ 237 ][ 37 ],
   alphaCSR[ 237 ][ 38 ],
   alphaCSR[ 237 ][ 39 ],
   alphaCSR[ 237 ][ 40 ],
   alphaCSR[ 237 ][ 41 ],
   alphaCSR[ 237 ][ 42 ],
   alphaCSR[ 237 ][ 43 ],
   alphaCSR[ 237 ][ 44 ],
   alphaCSR[ 237 ][ 45 ],
   alphaCSR[ 237 ][ 46 ],
   alphaCSR[ 237 ][ 47 ],
   alphaCSR[ 237 ][ 48 ],
   alphaCSR[ 237 ][ 49 ],
   alphaCSR[ 237 ][ 50 ],
   alphaCSR[ 237 ][ 51 ],
   alphaCSR[ 237 ][ 52 ],
   alphaCSR[ 237 ][ 53 ],
   alphaCSR[ 237 ][ 54 ],
   alphaCSR[ 237 ][ 55 ],
   alphaCSR[ 237 ][ 56 ],
   alphaCSR[ 237 ][ 57 ],
   alphaCSR[ 237 ][ 58 ],
   alphaCSR[ 237 ][ 59 ],
   alphaCSR[ 237 ][ 60 ],
   alphaCSR[ 237 ][ 61 ],
   alphaCSR[ 237 ][ 62 ],
   alphaCSR[ 237 ][ 63 ],
   alphaCSR[ 237 ][ 64 ],
   alphaCSR[ 237 ][ 65 ],
   alphaCSR[ 237 ][ 66 ],
   alphaCSR[ 237 ][ 67 ],
   alphaCSR[ 237 ][ 68 ],
   alphaCSR[ 237 ][ 69 ],
   alphaCSR[ 237 ][ 70 ],
   alphaCSR[ 237 ][ 71 ],
   alphaCSR[ 237 ][ 72 ],
   alphaCSR[ 237 ][ 73 ],
   alphaCSR[ 237 ][ 74 ],
   alphaCSR[ 237 ][ 75 ],
   alphaCSR[ 237 ][ 76 ],
   alphaCSR[ 237 ][ 77 ],
   alphaCSR[ 237 ][ 78 ],
   alphaCSR[ 237 ][ 79 ],
   alphaCSR[ 237 ][ 80 ],
   alphaCSR[ 237 ][ 81 ],
   alphaCSR[ 237 ][ 82 ],
   alphaCSR[ 237 ][ 83 ],
   alphaCSR[ 237 ][ 84 ],
   alphaCSR[ 237 ][ 85 ],
   alphaCSR[ 237 ][ 86 ],
   alphaCSR[ 237 ][ 87 ],
   alphaCSR[ 237 ][ 88 ],
   alphaCSR[ 237 ][ 89 ],
   alphaCSR[ 237 ][ 90 ],
   alphaCSR[ 237 ][ 91 ],
   alphaCSR[ 237 ][ 92 ],
   alphaCSR[ 237 ][ 93 ],
   alphaCSR[ 237 ][ 94 ],
   alphaCSR[ 237 ][ 95 ],
   alphaCSR[ 237 ][ 96 ],
   alphaCSR[ 237 ][ 97 ],
   alphaCSR[ 237 ][ 98 ],
   alphaCSR[ 237 ][ 99 ],
   alphaCSR[ 237 ][ 100 ],
   alphaCSR[ 237 ][ 101 ],
   alphaCSR[ 237 ][ 102 ],
   alphaCSR[ 237 ][ 103 ],
   alphaCSR[ 237 ][ 104 ],
   alphaCSR[ 237 ][ 105 ],
   alphaCSR[ 237 ][ 106 ],
   alphaCSR[ 237 ][ 107 ],
   alphaCSR[ 237 ][ 108 ],
   alphaCSR[ 237 ][ 109 ],
   alphaCSR[ 237 ][ 110 ],
   alphaCSR[ 237 ][ 111 ],
   alphaCSR[ 237 ][ 112 ],
   alphaCSR[ 237 ][ 113 ],
   alphaCSR[ 237 ][ 114 ],
   alphaCSR[ 237 ][ 115 ],
   alphaCSR[ 237 ][ 116 ],
   alphaCSR[ 237 ][ 117 ],
   alphaCSR[ 237 ][ 118 ],
   alphaCSR[ 237 ][ 119 ],
   alphaCSR[ 237 ][ 120 ],
   alphaCSR[ 237 ][ 121 ],
   alphaCSR[ 237 ][ 122 ],
   alphaCSR[ 237 ][ 123 ],
   alphaCSR[ 237 ][ 124 ],
   alphaCSR[ 237 ][ 125 ],
   alphaCSR[ 237 ][ 126 ],
   alphaCSR[ 237 ][ 127 ],
   alphaCSR[ 237 ][ 128 ],
   alphaCSR[ 237 ][ 129 ],
   alphaCSR[ 237 ][ 130 ],
   alphaCSR[ 237 ][ 131 ],
   alphaCSR[ 237 ][ 132 ],
   alphaCSR[ 237 ][ 133 ],
   alphaCSR[ 237 ][ 134 ],
   alphaCSR[ 237 ][ 135 ],
   alphaCSR[ 237 ][ 136 ],
   alphaCSR[ 237 ][ 137 ],
   alphaCSR[ 237 ][ 138 ],
   alphaCSR[ 237 ][ 139 ],
   alphaCSR[ 237 ][ 140 ],
   alphaCSR[ 237 ][ 141 ],
   alphaCSR[ 237 ][ 142 ],
   alphaCSR[ 237 ][ 143 ],
   alphaCSR[ 237 ][ 144 ],
   alphaCSR[ 237 ][ 145 ],
   alphaCSR[ 237 ][ 146 ],
   alphaCSR[ 237 ][ 147 ],
   alphaCSR[ 237 ][ 148 ],
   alphaCSR[ 237 ][ 149 ],
   alphaCSR[ 237 ][ 150 ],
   alphaCSR[ 237 ][ 151 ],
   alphaCSR[ 237 ][ 152 ],
   alphaCSR[ 237 ][ 153 ],
   alphaCSR[ 237 ][ 154 ],
   alphaCSR[ 237 ][ 155 ],
   alphaCSR[ 237 ][ 156 ],
   alphaCSR[ 237 ][ 157 ],
   alphaCSR[ 237 ][ 158 ],
   alphaCSR[ 237 ][ 159 ],
   alphaCSR[ 237 ][ 160 ],
   alphaCSR[ 237 ][ 161 ],
   alphaCSR[ 237 ][ 162 ],
   alphaCSR[ 237 ][ 163 ],
   alphaCSR[ 237 ][ 164 ],
   alphaCSR[ 237 ][ 165 ],
   alphaCSR[ 237 ][ 166 ],
   alphaCSR[ 237 ][ 167 ],
   alphaCSR[ 237 ][ 168 ],
   alphaCSR[ 237 ][ 169 ],
   alphaCSR[ 237 ][ 170 ],
   alphaCSR[ 237 ][ 171 ],
   alphaCSR[ 237 ][ 172 ],
   alphaCSR[ 237 ][ 173 ],
   alphaCSR[ 237 ][ 174 ],
   alphaCSR[ 237 ][ 175 ],
   alphaCSR[ 237 ][ 176 ],
   alphaCSR[ 237 ][ 177 ],
   alphaCSR[ 237 ][ 178 ],
   alphaCSR[ 237 ][ 179 ],
   alphaCSR[ 237 ][ 180 ],
   alphaCSR[ 237 ][ 181 ],
   alphaCSR[ 237 ][ 182 ],
   alphaCSR[ 237 ][ 183 ],
   alphaCSR[ 237 ][ 184 ],
   alphaCSR[ 237 ][ 185 ],
   alphaCSR[ 237 ][ 186 ],
   alphaCSR[ 237 ][ 187 ],
   alphaCSR[ 237 ][ 188 ],
   alphaCSR[ 237 ][ 189 ],
   alphaCSR[ 237 ][ 190 ],
   alphaCSR[ 237 ][ 191 ],
   alphaCSR[ 237 ][ 192 ],
   alphaCSR[ 237 ][ 193 ],
   alphaCSR[ 237 ][ 194 ],
   alphaCSR[ 237 ][ 195 ],
   alphaCSR[ 237 ][ 196 ],
   alphaCSR[ 237 ][ 197 ],
   alphaCSR[ 237 ][ 198 ],
   alphaCSR[ 237 ][ 199 ],
   alphaCSR[ 237 ][ 200 ],
   alphaCSR[ 237 ][ 201 ],
   alphaCSR[ 237 ][ 202 ],
   alphaCSR[ 237 ][ 203 ],
   alphaCSR[ 237 ][ 204 ],
   alphaCSR[ 237 ][ 205 ],
   alphaCSR[ 237 ][ 206 ],
   alphaCSR[ 237 ][ 207 ],
   alphaCSR[ 237 ][ 208 ],
   alphaCSR[ 237 ][ 209 ],
   alphaCSR[ 237 ][ 210 ],
   alphaCSR[ 237 ][ 211 ],
   alphaCSR[ 237 ][ 212 ],
   alphaCSR[ 237 ][ 213 ],
   alphaCSR[ 237 ][ 214 ],
   alphaCSR[ 237 ][ 215 ],
   alphaCSR[ 237 ][ 216 ],
   alphaCSR[ 237 ][ 217 ],
   alphaCSR[ 237 ][ 218 ],
   alphaCSR[ 237 ][ 219 ],
   alphaCSR[ 237 ][ 220 ],
   alphaCSR[ 237 ][ 221 ],
   alphaCSR[ 237 ][ 222 ],
   alphaCSR[ 237 ][ 223 ],
   alphaCSR[ 237 ][ 224 ],
   alphaCSR[ 237 ][ 225 ],
   alphaCSR[ 237 ][ 226 ],
   alphaCSR[ 237 ][ 227 ],
   alphaCSR[ 237 ][ 228 ],
   alphaCSR[ 237 ][ 229 ],
   alphaCSR[ 237 ][ 230 ],
   alphaCSR[ 237 ][ 231 ],
   alphaCSR[ 237 ][ 232 ],
   alphaCSR[ 237 ][ 233 ],
   alphaCSR[ 237 ][ 234 ],
   alphaCSR[ 237 ][ 235 ],
   alphaCSR[ 237 ][ 236 ],
   alphaCSR[ 237 ][ 237 ],
   alphaCSR[ 237 ][ 238 ],
   alphaCSR[ 237 ][ 239 ],
   alphaCSR[ 237 ][ 240 ],
   alphaCSR[ 237 ][ 241 ],
   alphaCSR[ 237 ][ 242 ],
   alphaCSR[ 237 ][ 243 ],
   alphaCSR[ 237 ][ 244 ],
   alphaCSR[ 237 ][ 245 ],
   alphaCSR[ 237 ][ 246 ],
   alphaCSR[ 237 ][ 247 ],
   alphaCSR[ 237 ][ 248 ],
   alphaCSR[ 237 ][ 249 ],
   alphaCSR[ 237 ][ 250 ],
   alphaCSR[ 237 ][ 251 ],
   alphaCSR[ 237 ][ 252 ],
   alphaCSR[ 237 ][ 253 ],
   alphaCSR[ 237 ][ 254 ],
   alphaCSR[ 237 ][ 255 ],
   alphaCSR[ 237 ][ 256 ],
   alphaCSR[ 237 ][ 257 ],
   alphaCSR[ 237 ][ 258 ],
   alphaCSR[ 237 ][ 259 ],
   alphaCSR[ 237 ][ 260 ],
   alphaCSR[ 237 ][ 261 ],
   alphaCSR[ 237 ][ 262 ],
   alphaCSR[ 237 ][ 263 ],
   alphaCSR[ 237 ][ 264 ],
   alphaCSR[ 237 ][ 265 ],
   alphaCSR[ 237 ][ 266 ],
   alphaCSR[ 237 ][ 267 ],
   alphaCSR[ 237 ][ 268 ],
   alphaCSR[ 237 ][ 269 ],
   alphaCSR[ 237 ][ 270 ],
   alphaCSR[ 237 ][ 271 ],
   alphaCSR[ 237 ][ 272 ],
   alphaCSR[ 237 ][ 273 ],
   alphaCSR[ 237 ][ 274 ],
   alphaCSR[ 237 ][ 275 ],
   alphaCSR[ 237 ][ 276 ],
   alphaCSR[ 237 ][ 277 ],
   alphaCSR[ 237 ][ 278 ],
   alphaCSR[ 237 ][ 279 ],
   alphaCSR[ 237 ][ 280 ],
   alphaCSR[ 237 ][ 281 ],
   alphaCSR[ 237 ][ 282 ],
   alphaCSR[ 237 ][ 283 ],
   alphaCSR[ 237 ][ 284 ],
   alphaCSR[ 237 ][ 285 ],
   alphaCSR[ 237 ][ 286 ],
   alphaCSR[ 237 ][ 287 ],
   alphaCSR[ 237 ][ 288 ],
   alphaCSR[ 237 ][ 289 ],
   alphaCSR[ 237 ][ 290 ],
   alphaCSR[ 237 ][ 291 ],
   alphaCSR[ 237 ][ 292 ],
   alphaCSR[ 237 ][ 293 ],
   alphaCSR[ 237 ][ 294 ],
   alphaCSR[ 237 ][ 295 ],
   alphaCSR[ 237 ][ 296 ],
   alphaCSR[ 237 ][ 297 ],
   alphaCSR[ 237 ][ 298 ],
   alphaCSR[ 237 ][ 299 ],
   alphaCSR[ 237 ][ 300 ],
   alphaCSR[ 237 ][ 301 ],
   alphaCSR[ 237 ][ 302 ],
   alphaCSR[ 237 ][ 303 ],
   alphaCSR[ 237 ][ 304 ],
   alphaCSR[ 237 ][ 305 ],
   alphaCSR[ 237 ][ 306 ],
   alphaCSR[ 237 ][ 307 ],
   alphaCSR[ 237 ][ 308 ],
   alphaCSR[ 237 ][ 309 ],
   alphaCSR[ 237 ][ 310 ],
   alphaCSR[ 237 ][ 311 ],
   alphaCSR[ 237 ][ 312 ],
   alphaCSR[ 237 ][ 313 ],
   alphaCSR[ 237 ][ 314 ],
   alphaCSR[ 237 ][ 315 ],
   alphaCSR[ 237 ][ 316 ],
   alphaCSR[ 237 ][ 317 ],
   alphaCSR[ 237 ][ 318 ],
   alphaCSR[ 237 ][ 319 ],
   alphaCSR[ 237 ][ 320 ],
   alphaCSR[ 237 ][ 321 ],
   alphaCSR[ 237 ][ 322 ],
   alphaCSR[ 237 ][ 323 ],
   alphaCSR[ 237 ][ 324 ],
   alphaCSR[ 237 ][ 325 ],
   alphaCSR[ 237 ][ 326 ],
   alphaCSR[ 237 ][ 327 ],
   alphaCSR[ 237 ][ 328 ],
   alphaCSR[ 237 ][ 329 ],
   alphaCSR[ 237 ][ 330 ],
   alphaCSR[ 237 ][ 331 ],
   alphaCSR[ 237 ][ 332 ],
   alphaCSR[ 237 ][ 333 ],
   alphaCSR[ 237 ][ 334 ],
   alphaCSR[ 237 ][ 335 ],
   alphaCSR[ 237 ][ 336 ],
   alphaCSR[ 237 ][ 337 ],
   alphaCSR[ 237 ][ 338 ],
   alphaCSR[ 237 ][ 339 ],
   alphaCSR[ 237 ][ 340 ],
   alphaCSR[ 237 ][ 341 ],
   alphaCSR[ 237 ][ 342 ],
   alphaCSR[ 237 ][ 343 ],
   alphaCSR[ 237 ][ 344 ],
   alphaCSR[ 237 ][ 345 ],
   alphaCSR[ 237 ][ 346 ],
   alphaCSR[ 237 ][ 347 ],
   alphaCSR[ 237 ][ 348 ],
   alphaCSR[ 237 ][ 349 ],
   alphaCSR[ 237 ][ 350 ],
   alphaCSR[ 237 ][ 351 ],
   alphaCSR[ 237 ][ 352 ],
   alphaCSR[ 237 ][ 353 ],
   alphaCSR[ 237 ][ 354 ],
   alphaCSR[ 237 ][ 355 ],
   alphaCSR[ 237 ][ 356 ],
   alphaCSR[ 237 ][ 357 ],
   alphaCSR[ 237 ][ 358 ],
   alphaCSR[ 237 ][ 359 ],
   alphaCSR[ 237 ][ 360 ],
   alphaCSR[ 237 ][ 361 ],
   alphaCSR[ 237 ][ 362 ],
   alphaCSR[ 237 ][ 363 ],
   alphaCSR[ 237 ][ 364 ],
   alphaCSR[ 237 ][ 365 ],
   alphaCSR[ 237 ][ 366 ],
   alphaCSR[ 237 ][ 367 ],
   alphaCSR[ 237 ][ 368 ],
   alphaCSR[ 237 ][ 369 ],
   alphaCSR[ 237 ][ 370 ],
   alphaCSR[ 237 ][ 371 ],
   alphaCSR[ 237 ][ 372 ],
   alphaCSR[ 237 ][ 373 ],
   alphaCSR[ 237 ][ 374 ],
   alphaCSR[ 237 ][ 375 ],
   alphaCSR[ 237 ][ 376 ],
   alphaCSR[ 237 ][ 377 ],
   alphaCSR[ 237 ][ 378 ],
   alphaCSR[ 237 ][ 379 ],
   alphaCSR[ 237 ][ 380 ],
   alphaCSR[ 237 ][ 381 ],
   alphaCSR[ 237 ][ 382 ],
   alphaCSR[ 237 ][ 383 ],
   alphaCSR[ 238 ][ 0 ],
   alphaCSR[ 238 ][ 1 ],
   alphaCSR[ 238 ][ 2 ],
   alphaCSR[ 238 ][ 3 ],
   alphaCSR[ 238 ][ 4 ],
   alphaCSR[ 238 ][ 5 ],
   alphaCSR[ 238 ][ 6 ],
   alphaCSR[ 238 ][ 7 ],
   alphaCSR[ 238 ][ 8 ],
   alphaCSR[ 238 ][ 9 ],
   alphaCSR[ 238 ][ 10 ],
   alphaCSR[ 238 ][ 11 ],
   alphaCSR[ 238 ][ 12 ],
   alphaCSR[ 238 ][ 13 ],
   alphaCSR[ 238 ][ 14 ],
   alphaCSR[ 238 ][ 15 ],
   alphaCSR[ 238 ][ 16 ],
   alphaCSR[ 238 ][ 17 ],
   alphaCSR[ 238 ][ 18 ],
   alphaCSR[ 238 ][ 19 ],
   alphaCSR[ 238 ][ 20 ],
   alphaCSR[ 238 ][ 21 ],
   alphaCSR[ 238 ][ 22 ],
   alphaCSR[ 238 ][ 23 ],
   alphaCSR[ 238 ][ 24 ],
   alphaCSR[ 238 ][ 25 ],
   alphaCSR[ 238 ][ 26 ],
   alphaCSR[ 238 ][ 27 ],
   alphaCSR[ 238 ][ 28 ],
   alphaCSR[ 238 ][ 29 ],
   alphaCSR[ 238 ][ 30 ],
   alphaCSR[ 238 ][ 31 ],
   alphaCSR[ 238 ][ 32 ],
   alphaCSR[ 238 ][ 33 ],
   alphaCSR[ 238 ][ 34 ],
   alphaCSR[ 238 ][ 35 ],
   alphaCSR[ 238 ][ 36 ],
   alphaCSR[ 238 ][ 37 ],
   alphaCSR[ 238 ][ 38 ],
   alphaCSR[ 238 ][ 39 ],
   alphaCSR[ 238 ][ 40 ],
   alphaCSR[ 238 ][ 41 ],
   alphaCSR[ 238 ][ 42 ],
   alphaCSR[ 238 ][ 43 ],
   alphaCSR[ 238 ][ 44 ],
   alphaCSR[ 238 ][ 45 ],
   alphaCSR[ 238 ][ 46 ],
   alphaCSR[ 238 ][ 47 ],
   alphaCSR[ 238 ][ 48 ],
   alphaCSR[ 238 ][ 49 ],
   alphaCSR[ 238 ][ 50 ],
   alphaCSR[ 238 ][ 51 ],
   alphaCSR[ 238 ][ 52 ],
   alphaCSR[ 238 ][ 53 ],
   alphaCSR[ 238 ][ 54 ],
   alphaCSR[ 238 ][ 55 ],
   alphaCSR[ 238 ][ 56 ],
   alphaCSR[ 238 ][ 57 ],
   alphaCSR[ 238 ][ 58 ],
   alphaCSR[ 238 ][ 59 ],
   alphaCSR[ 238 ][ 60 ],
   alphaCSR[ 238 ][ 61 ],
   alphaCSR[ 238 ][ 62 ],
   alphaCSR[ 238 ][ 63 ],
   alphaCSR[ 238 ][ 64 ],
   alphaCSR[ 238 ][ 65 ],
   alphaCSR[ 238 ][ 66 ],
   alphaCSR[ 238 ][ 67 ],
   alphaCSR[ 238 ][ 68 ],
   alphaCSR[ 238 ][ 69 ],
   alphaCSR[ 238 ][ 70 ],
   alphaCSR[ 238 ][ 71 ],
   alphaCSR[ 238 ][ 72 ],
   alphaCSR[ 238 ][ 73 ],
   alphaCSR[ 238 ][ 74 ],
   alphaCSR[ 238 ][ 75 ],
   alphaCSR[ 238 ][ 76 ],
   alphaCSR[ 238 ][ 77 ],
   alphaCSR[ 238 ][ 78 ],
   alphaCSR[ 238 ][ 79 ],
   alphaCSR[ 238 ][ 80 ],
   alphaCSR[ 238 ][ 81 ],
   alphaCSR[ 238 ][ 82 ],
   alphaCSR[ 238 ][ 83 ],
   alphaCSR[ 238 ][ 84 ],
   alphaCSR[ 238 ][ 85 ],
   alphaCSR[ 238 ][ 86 ],
   alphaCSR[ 238 ][ 87 ],
   alphaCSR[ 238 ][ 88 ],
   alphaCSR[ 238 ][ 89 ],
   alphaCSR[ 238 ][ 90 ],
   alphaCSR[ 238 ][ 91 ],
   alphaCSR[ 238 ][ 92 ],
   alphaCSR[ 238 ][ 93 ],
   alphaCSR[ 238 ][ 94 ],
   alphaCSR[ 238 ][ 95 ],
   alphaCSR[ 238 ][ 96 ],
   alphaCSR[ 238 ][ 97 ],
   alphaCSR[ 238 ][ 98 ],
   alphaCSR[ 238 ][ 99 ],
   alphaCSR[ 238 ][ 100 ],
   alphaCSR[ 238 ][ 101 ],
   alphaCSR[ 238 ][ 102 ],
   alphaCSR[ 238 ][ 103 ],
   alphaCSR[ 238 ][ 104 ],
   alphaCSR[ 238 ][ 105 ],
   alphaCSR[ 238 ][ 106 ],
   alphaCSR[ 238 ][ 107 ],
   alphaCSR[ 238 ][ 108 ],
   alphaCSR[ 238 ][ 109 ],
   alphaCSR[ 238 ][ 110 ],
   alphaCSR[ 238 ][ 111 ],
   alphaCSR[ 238 ][ 112 ],
   alphaCSR[ 238 ][ 113 ],
   alphaCSR[ 238 ][ 114 ],
   alphaCSR[ 238 ][ 115 ],
   alphaCSR[ 238 ][ 116 ],
   alphaCSR[ 238 ][ 117 ],
   alphaCSR[ 238 ][ 118 ],
   alphaCSR[ 238 ][ 119 ],
   alphaCSR[ 238 ][ 120 ],
   alphaCSR[ 238 ][ 121 ],
   alphaCSR[ 238 ][ 122 ],
   alphaCSR[ 238 ][ 123 ],
   alphaCSR[ 238 ][ 124 ],
   alphaCSR[ 238 ][ 125 ],
   alphaCSR[ 238 ][ 126 ],
   alphaCSR[ 238 ][ 127 ],
   alphaCSR[ 238 ][ 128 ],
   alphaCSR[ 238 ][ 129 ],
   alphaCSR[ 238 ][ 130 ],
   alphaCSR[ 238 ][ 131 ],
   alphaCSR[ 238 ][ 132 ],
   alphaCSR[ 238 ][ 133 ],
   alphaCSR[ 238 ][ 134 ],
   alphaCSR[ 238 ][ 135 ],
   alphaCSR[ 238 ][ 136 ],
   alphaCSR[ 238 ][ 137 ],
   alphaCSR[ 238 ][ 138 ],
   alphaCSR[ 238 ][ 139 ],
   alphaCSR[ 238 ][ 140 ],
   alphaCSR[ 238 ][ 141 ],
   alphaCSR[ 238 ][ 142 ],
   alphaCSR[ 238 ][ 143 ],
   alphaCSR[ 238 ][ 144 ],
   alphaCSR[ 238 ][ 145 ],
   alphaCSR[ 238 ][ 146 ],
   alphaCSR[ 238 ][ 147 ],
   alphaCSR[ 238 ][ 148 ],
   alphaCSR[ 238 ][ 149 ],
   alphaCSR[ 238 ][ 150 ],
   alphaCSR[ 238 ][ 151 ],
   alphaCSR[ 238 ][ 152 ],
   alphaCSR[ 238 ][ 153 ],
   alphaCSR[ 238 ][ 154 ],
   alphaCSR[ 238 ][ 155 ],
   alphaCSR[ 238 ][ 156 ],
   alphaCSR[ 238 ][ 157 ],
   alphaCSR[ 238 ][ 158 ],
   alphaCSR[ 238 ][ 159 ],
   alphaCSR[ 238 ][ 160 ],
   alphaCSR[ 238 ][ 161 ],
   alphaCSR[ 238 ][ 162 ],
   alphaCSR[ 238 ][ 163 ],
   alphaCSR[ 238 ][ 164 ],
   alphaCSR[ 238 ][ 165 ],
   alphaCSR[ 238 ][ 166 ],
   alphaCSR[ 238 ][ 167 ],
   alphaCSR[ 238 ][ 168 ],
   alphaCSR[ 238 ][ 169 ],
   alphaCSR[ 238 ][ 170 ],
   alphaCSR[ 238 ][ 171 ],
   alphaCSR[ 238 ][ 172 ],
   alphaCSR[ 238 ][ 173 ],
   alphaCSR[ 238 ][ 174 ],
   alphaCSR[ 238 ][ 175 ],
   alphaCSR[ 238 ][ 176 ],
   alphaCSR[ 238 ][ 177 ],
   alphaCSR[ 238 ][ 178 ],
   alphaCSR[ 238 ][ 179 ],
   alphaCSR[ 238 ][ 180 ],
   alphaCSR[ 238 ][ 181 ],
   alphaCSR[ 238 ][ 182 ],
   alphaCSR[ 238 ][ 183 ],
   alphaCSR[ 238 ][ 184 ],
   alphaCSR[ 238 ][ 185 ],
   alphaCSR[ 238 ][ 186 ],
   alphaCSR[ 238 ][ 187 ],
   alphaCSR[ 238 ][ 188 ],
   alphaCSR[ 238 ][ 189 ],
   alphaCSR[ 238 ][ 190 ],
   alphaCSR[ 238 ][ 191 ],
   alphaCSR[ 238 ][ 192 ],
   alphaCSR[ 238 ][ 193 ],
   alphaCSR[ 238 ][ 194 ],
   alphaCSR[ 238 ][ 195 ],
   alphaCSR[ 238 ][ 196 ],
   alphaCSR[ 238 ][ 197 ],
   alphaCSR[ 238 ][ 198 ],
   alphaCSR[ 238 ][ 199 ],
   alphaCSR[ 238 ][ 200 ],
   alphaCSR[ 238 ][ 201 ],
   alphaCSR[ 238 ][ 202 ],
   alphaCSR[ 238 ][ 203 ],
   alphaCSR[ 238 ][ 204 ],
   alphaCSR[ 238 ][ 205 ],
   alphaCSR[ 238 ][ 206 ],
   alphaCSR[ 238 ][ 207 ],
   alphaCSR[ 238 ][ 208 ],
   alphaCSR[ 238 ][ 209 ],
   alphaCSR[ 238 ][ 210 ],
   alphaCSR[ 238 ][ 211 ],
   alphaCSR[ 238 ][ 212 ],
   alphaCSR[ 238 ][ 213 ],
   alphaCSR[ 238 ][ 214 ],
   alphaCSR[ 238 ][ 215 ],
   alphaCSR[ 238 ][ 216 ],
   alphaCSR[ 238 ][ 217 ],
   alphaCSR[ 238 ][ 218 ],
   alphaCSR[ 238 ][ 219 ],
   alphaCSR[ 238 ][ 220 ],
   alphaCSR[ 238 ][ 221 ],
   alphaCSR[ 238 ][ 222 ],
   alphaCSR[ 238 ][ 223 ],
   alphaCSR[ 238 ][ 224 ],
   alphaCSR[ 238 ][ 225 ],
   alphaCSR[ 238 ][ 226 ],
   alphaCSR[ 238 ][ 227 ],
   alphaCSR[ 238 ][ 228 ],
   alphaCSR[ 238 ][ 229 ],
   alphaCSR[ 238 ][ 230 ],
   alphaCSR[ 238 ][ 231 ],
   alphaCSR[ 238 ][ 232 ],
   alphaCSR[ 238 ][ 233 ],
   alphaCSR[ 238 ][ 234 ],
   alphaCSR[ 238 ][ 235 ],
   alphaCSR[ 238 ][ 236 ],
   alphaCSR[ 238 ][ 237 ],
   alphaCSR[ 238 ][ 238 ],
   alphaCSR[ 238 ][ 239 ],
   alphaCSR[ 238 ][ 240 ],
   alphaCSR[ 238 ][ 241 ],
   alphaCSR[ 238 ][ 242 ],
   alphaCSR[ 238 ][ 243 ],
   alphaCSR[ 238 ][ 244 ],
   alphaCSR[ 238 ][ 245 ],
   alphaCSR[ 238 ][ 246 ],
   alphaCSR[ 238 ][ 247 ],
   alphaCSR[ 238 ][ 248 ],
   alphaCSR[ 238 ][ 249 ],
   alphaCSR[ 238 ][ 250 ],
   alphaCSR[ 238 ][ 251 ],
   alphaCSR[ 238 ][ 252 ],
   alphaCSR[ 238 ][ 253 ],
   alphaCSR[ 238 ][ 254 ],
   alphaCSR[ 238 ][ 255 ],
   alphaCSR[ 238 ][ 256 ],
   alphaCSR[ 238 ][ 257 ],
   alphaCSR[ 238 ][ 258 ],
   alphaCSR[ 238 ][ 259 ],
   alphaCSR[ 238 ][ 260 ],
   alphaCSR[ 238 ][ 261 ],
   alphaCSR[ 238 ][ 262 ],
   alphaCSR[ 238 ][ 263 ],
   alphaCSR[ 238 ][ 264 ],
   alphaCSR[ 238 ][ 265 ],
   alphaCSR[ 238 ][ 266 ],
   alphaCSR[ 238 ][ 267 ],
   alphaCSR[ 238 ][ 268 ],
   alphaCSR[ 238 ][ 269 ],
   alphaCSR[ 238 ][ 270 ],
   alphaCSR[ 238 ][ 271 ],
   alphaCSR[ 238 ][ 272 ],
   alphaCSR[ 238 ][ 273 ],
   alphaCSR[ 238 ][ 274 ],
   alphaCSR[ 238 ][ 275 ],
   alphaCSR[ 238 ][ 276 ],
   alphaCSR[ 238 ][ 277 ],
   alphaCSR[ 238 ][ 278 ],
   alphaCSR[ 238 ][ 279 ],
   alphaCSR[ 238 ][ 280 ],
   alphaCSR[ 238 ][ 281 ],
   alphaCSR[ 238 ][ 282 ],
   alphaCSR[ 238 ][ 283 ],
   alphaCSR[ 238 ][ 284 ],
   alphaCSR[ 238 ][ 285 ],
   alphaCSR[ 238 ][ 286 ],
   alphaCSR[ 238 ][ 287 ],
   alphaCSR[ 238 ][ 288 ],
   alphaCSR[ 238 ][ 289 ],
   alphaCSR[ 238 ][ 290 ],
   alphaCSR[ 238 ][ 291 ],
   alphaCSR[ 238 ][ 292 ],
   alphaCSR[ 238 ][ 293 ],
   alphaCSR[ 238 ][ 294 ],
   alphaCSR[ 238 ][ 295 ],
   alphaCSR[ 238 ][ 296 ],
   alphaCSR[ 238 ][ 297 ],
   alphaCSR[ 238 ][ 298 ],
   alphaCSR[ 238 ][ 299 ],
   alphaCSR[ 238 ][ 300 ],
   alphaCSR[ 238 ][ 301 ],
   alphaCSR[ 238 ][ 302 ],
   alphaCSR[ 238 ][ 303 ],
   alphaCSR[ 238 ][ 304 ],
   alphaCSR[ 238 ][ 305 ],
   alphaCSR[ 238 ][ 306 ],
   alphaCSR[ 238 ][ 307 ],
   alphaCSR[ 238 ][ 308 ],
   alphaCSR[ 238 ][ 309 ],
   alphaCSR[ 238 ][ 310 ],
   alphaCSR[ 238 ][ 311 ],
   alphaCSR[ 238 ][ 312 ],
   alphaCSR[ 238 ][ 313 ],
   alphaCSR[ 238 ][ 314 ],
   alphaCSR[ 238 ][ 315 ],
   alphaCSR[ 238 ][ 316 ],
   alphaCSR[ 238 ][ 317 ],
   alphaCSR[ 238 ][ 318 ],
   alphaCSR[ 238 ][ 319 ],
   alphaCSR[ 238 ][ 320 ],
   alphaCSR[ 238 ][ 321 ],
   alphaCSR[ 238 ][ 322 ],
   alphaCSR[ 238 ][ 323 ],
   alphaCSR[ 238 ][ 324 ],
   alphaCSR[ 238 ][ 325 ],
   alphaCSR[ 238 ][ 326 ],
   alphaCSR[ 238 ][ 327 ],
   alphaCSR[ 238 ][ 328 ],
   alphaCSR[ 238 ][ 329 ],
   alphaCSR[ 238 ][ 330 ],
   alphaCSR[ 238 ][ 331 ],
   alphaCSR[ 238 ][ 332 ],
   alphaCSR[ 238 ][ 333 ],
   alphaCSR[ 238 ][ 334 ],
   alphaCSR[ 238 ][ 335 ],
   alphaCSR[ 238 ][ 336 ],
   alphaCSR[ 238 ][ 337 ],
   alphaCSR[ 238 ][ 338 ],
   alphaCSR[ 238 ][ 339 ],
   alphaCSR[ 238 ][ 340 ],
   alphaCSR[ 238 ][ 341 ],
   alphaCSR[ 238 ][ 342 ],
   alphaCSR[ 238 ][ 343 ],
   alphaCSR[ 238 ][ 344 ],
   alphaCSR[ 238 ][ 345 ],
   alphaCSR[ 238 ][ 346 ],
   alphaCSR[ 238 ][ 347 ],
   alphaCSR[ 238 ][ 348 ],
   alphaCSR[ 238 ][ 349 ],
   alphaCSR[ 238 ][ 350 ],
   alphaCSR[ 238 ][ 351 ],
   alphaCSR[ 238 ][ 352 ],
   alphaCSR[ 238 ][ 353 ],
   alphaCSR[ 238 ][ 354 ],
   alphaCSR[ 238 ][ 355 ],
   alphaCSR[ 238 ][ 356 ],
   alphaCSR[ 238 ][ 357 ],
   alphaCSR[ 238 ][ 358 ],
   alphaCSR[ 238 ][ 359 ],
   alphaCSR[ 238 ][ 360 ],
   alphaCSR[ 238 ][ 361 ],
   alphaCSR[ 238 ][ 362 ],
   alphaCSR[ 238 ][ 363 ],
   alphaCSR[ 238 ][ 364 ],
   alphaCSR[ 238 ][ 365 ],
   alphaCSR[ 238 ][ 366 ],
   alphaCSR[ 238 ][ 367 ],
   alphaCSR[ 238 ][ 368 ],
   alphaCSR[ 238 ][ 369 ],
   alphaCSR[ 238 ][ 370 ],
   alphaCSR[ 238 ][ 371 ],
   alphaCSR[ 238 ][ 372 ],
   alphaCSR[ 238 ][ 373 ],
   alphaCSR[ 238 ][ 374 ],
   alphaCSR[ 238 ][ 375 ],
   alphaCSR[ 238 ][ 376 ],
   alphaCSR[ 238 ][ 377 ],
   alphaCSR[ 238 ][ 378 ],
   alphaCSR[ 238 ][ 379 ],
   alphaCSR[ 238 ][ 380 ],
   alphaCSR[ 238 ][ 381 ],
   alphaCSR[ 238 ][ 382 ],
   alphaCSR[ 238 ][ 383 ],
   alphaCSR[ 239 ][ 0 ],
   alphaCSR[ 239 ][ 1 ],
   alphaCSR[ 239 ][ 2 ],
   alphaCSR[ 239 ][ 3 ],
   alphaCSR[ 239 ][ 4 ],
   alphaCSR[ 239 ][ 5 ],
   alphaCSR[ 239 ][ 6 ],
   alphaCSR[ 239 ][ 7 ],
   alphaCSR[ 239 ][ 8 ],
   alphaCSR[ 239 ][ 9 ],
   alphaCSR[ 239 ][ 10 ],
   alphaCSR[ 239 ][ 11 ],
   alphaCSR[ 239 ][ 12 ],
   alphaCSR[ 239 ][ 13 ],
   alphaCSR[ 239 ][ 14 ],
   alphaCSR[ 239 ][ 15 ],
   alphaCSR[ 239 ][ 16 ],
   alphaCSR[ 239 ][ 17 ],
   alphaCSR[ 239 ][ 18 ],
   alphaCSR[ 239 ][ 19 ],
   alphaCSR[ 239 ][ 20 ],
   alphaCSR[ 239 ][ 21 ],
   alphaCSR[ 239 ][ 22 ],
   alphaCSR[ 239 ][ 23 ],
   alphaCSR[ 239 ][ 24 ],
   alphaCSR[ 239 ][ 25 ],
   alphaCSR[ 239 ][ 26 ],
   alphaCSR[ 239 ][ 27 ],
   alphaCSR[ 239 ][ 28 ],
   alphaCSR[ 239 ][ 29 ],
   alphaCSR[ 239 ][ 30 ],
   alphaCSR[ 239 ][ 31 ],
   alphaCSR[ 239 ][ 32 ],
   alphaCSR[ 239 ][ 33 ],
   alphaCSR[ 239 ][ 34 ],
   alphaCSR[ 239 ][ 35 ],
   alphaCSR[ 239 ][ 36 ],
   alphaCSR[ 239 ][ 37 ],
   alphaCSR[ 239 ][ 38 ],
   alphaCSR[ 239 ][ 39 ],
   alphaCSR[ 239 ][ 40 ],
   alphaCSR[ 239 ][ 41 ],
   alphaCSR[ 239 ][ 42 ],
   alphaCSR[ 239 ][ 43 ],
   alphaCSR[ 239 ][ 44 ],
   alphaCSR[ 239 ][ 45 ],
   alphaCSR[ 239 ][ 46 ],
   alphaCSR[ 239 ][ 47 ],
   alphaCSR[ 239 ][ 48 ],
   alphaCSR[ 239 ][ 49 ],
   alphaCSR[ 239 ][ 50 ],
   alphaCSR[ 239 ][ 51 ],
   alphaCSR[ 239 ][ 52 ],
   alphaCSR[ 239 ][ 53 ],
   alphaCSR[ 239 ][ 54 ],
   alphaCSR[ 239 ][ 55 ],
   alphaCSR[ 239 ][ 56 ],
   alphaCSR[ 239 ][ 57 ],
   alphaCSR[ 239 ][ 58 ],
   alphaCSR[ 239 ][ 59 ],
   alphaCSR[ 239 ][ 60 ],
   alphaCSR[ 239 ][ 61 ],
   alphaCSR[ 239 ][ 62 ],
   alphaCSR[ 239 ][ 63 ],
   alphaCSR[ 239 ][ 64 ],
   alphaCSR[ 239 ][ 65 ],
   alphaCSR[ 239 ][ 66 ],
   alphaCSR[ 239 ][ 67 ],
   alphaCSR[ 239 ][ 68 ],
   alphaCSR[ 239 ][ 69 ],
   alphaCSR[ 239 ][ 70 ],
   alphaCSR[ 239 ][ 71 ],
   alphaCSR[ 239 ][ 72 ],
   alphaCSR[ 239 ][ 73 ],
   alphaCSR[ 239 ][ 74 ],
   alphaCSR[ 239 ][ 75 ],
   alphaCSR[ 239 ][ 76 ],
   alphaCSR[ 239 ][ 77 ],
   alphaCSR[ 239 ][ 78 ],
   alphaCSR[ 239 ][ 79 ],
   alphaCSR[ 239 ][ 80 ],
   alphaCSR[ 239 ][ 81 ],
   alphaCSR[ 239 ][ 82 ],
   alphaCSR[ 239 ][ 83 ],
   alphaCSR[ 239 ][ 84 ],
   alphaCSR[ 239 ][ 85 ],
   alphaCSR[ 239 ][ 86 ],
   alphaCSR[ 239 ][ 87 ],
   alphaCSR[ 239 ][ 88 ],
   alphaCSR[ 239 ][ 89 ],
   alphaCSR[ 239 ][ 90 ],
   alphaCSR[ 239 ][ 91 ],
   alphaCSR[ 239 ][ 92 ],
   alphaCSR[ 239 ][ 93 ],
   alphaCSR[ 239 ][ 94 ],
   alphaCSR[ 239 ][ 95 ],
   alphaCSR[ 239 ][ 96 ],
   alphaCSR[ 239 ][ 97 ],
   alphaCSR[ 239 ][ 98 ],
   alphaCSR[ 239 ][ 99 ],
   alphaCSR[ 239 ][ 100 ],
   alphaCSR[ 239 ][ 101 ],
   alphaCSR[ 239 ][ 102 ],
   alphaCSR[ 239 ][ 103 ],
   alphaCSR[ 239 ][ 104 ],
   alphaCSR[ 239 ][ 105 ],
   alphaCSR[ 239 ][ 106 ],
   alphaCSR[ 239 ][ 107 ],
   alphaCSR[ 239 ][ 108 ],
   alphaCSR[ 239 ][ 109 ],
   alphaCSR[ 239 ][ 110 ],
   alphaCSR[ 239 ][ 111 ],
   alphaCSR[ 239 ][ 112 ],
   alphaCSR[ 239 ][ 113 ],
   alphaCSR[ 239 ][ 114 ],
   alphaCSR[ 239 ][ 115 ],
   alphaCSR[ 239 ][ 116 ],
   alphaCSR[ 239 ][ 117 ],
   alphaCSR[ 239 ][ 118 ],
   alphaCSR[ 239 ][ 119 ],
   alphaCSR[ 239 ][ 120 ],
   alphaCSR[ 239 ][ 121 ],
   alphaCSR[ 239 ][ 122 ],
   alphaCSR[ 239 ][ 123 ],
   alphaCSR[ 239 ][ 124 ],
   alphaCSR[ 239 ][ 125 ],
   alphaCSR[ 239 ][ 126 ],
   alphaCSR[ 239 ][ 127 ],
   alphaCSR[ 239 ][ 128 ],
   alphaCSR[ 239 ][ 129 ],
   alphaCSR[ 239 ][ 130 ],
   alphaCSR[ 239 ][ 131 ],
   alphaCSR[ 239 ][ 132 ],
   alphaCSR[ 239 ][ 133 ],
   alphaCSR[ 239 ][ 134 ],
   alphaCSR[ 239 ][ 135 ],
   alphaCSR[ 239 ][ 136 ],
   alphaCSR[ 239 ][ 137 ],
   alphaCSR[ 239 ][ 138 ],
   alphaCSR[ 239 ][ 139 ],
   alphaCSR[ 239 ][ 140 ],
   alphaCSR[ 239 ][ 141 ],
   alphaCSR[ 239 ][ 142 ],
   alphaCSR[ 239 ][ 143 ],
   alphaCSR[ 239 ][ 144 ],
   alphaCSR[ 239 ][ 145 ],
   alphaCSR[ 239 ][ 146 ],
   alphaCSR[ 239 ][ 147 ],
   alphaCSR[ 239 ][ 148 ],
   alphaCSR[ 239 ][ 149 ],
   alphaCSR[ 239 ][ 150 ],
   alphaCSR[ 239 ][ 151 ],
   alphaCSR[ 239 ][ 152 ],
   alphaCSR[ 239 ][ 153 ],
   alphaCSR[ 239 ][ 154 ],
   alphaCSR[ 239 ][ 155 ],
   alphaCSR[ 239 ][ 156 ],
   alphaCSR[ 239 ][ 157 ],
   alphaCSR[ 239 ][ 158 ],
   alphaCSR[ 239 ][ 159 ],
   alphaCSR[ 239 ][ 160 ],
   alphaCSR[ 239 ][ 161 ],
   alphaCSR[ 239 ][ 162 ],
   alphaCSR[ 239 ][ 163 ],
   alphaCSR[ 239 ][ 164 ],
   alphaCSR[ 239 ][ 165 ],
   alphaCSR[ 239 ][ 166 ],
   alphaCSR[ 239 ][ 167 ],
   alphaCSR[ 239 ][ 168 ],
   alphaCSR[ 239 ][ 169 ],
   alphaCSR[ 239 ][ 170 ],
   alphaCSR[ 239 ][ 171 ],
   alphaCSR[ 239 ][ 172 ],
   alphaCSR[ 239 ][ 173 ],
   alphaCSR[ 239 ][ 174 ],
   alphaCSR[ 239 ][ 175 ],
   alphaCSR[ 239 ][ 176 ],
   alphaCSR[ 239 ][ 177 ],
   alphaCSR[ 239 ][ 178 ],
   alphaCSR[ 239 ][ 179 ],
   alphaCSR[ 239 ][ 180 ],
   alphaCSR[ 239 ][ 181 ],
   alphaCSR[ 239 ][ 182 ],
   alphaCSR[ 239 ][ 183 ],
   alphaCSR[ 239 ][ 184 ],
   alphaCSR[ 239 ][ 185 ],
   alphaCSR[ 239 ][ 186 ],
   alphaCSR[ 239 ][ 187 ],
   alphaCSR[ 239 ][ 188 ],
   alphaCSR[ 239 ][ 189 ],
   alphaCSR[ 239 ][ 190 ],
   alphaCSR[ 239 ][ 191 ],
   alphaCSR[ 239 ][ 192 ],
   alphaCSR[ 239 ][ 193 ],
   alphaCSR[ 239 ][ 194 ],
   alphaCSR[ 239 ][ 195 ],
   alphaCSR[ 239 ][ 196 ],
   alphaCSR[ 239 ][ 197 ],
   alphaCSR[ 239 ][ 198 ],
   alphaCSR[ 239 ][ 199 ],
   alphaCSR[ 239 ][ 200 ],
   alphaCSR[ 239 ][ 201 ],
   alphaCSR[ 239 ][ 202 ],
   alphaCSR[ 239 ][ 203 ],
   alphaCSR[ 239 ][ 204 ],
   alphaCSR[ 239 ][ 205 ],
   alphaCSR[ 239 ][ 206 ],
   alphaCSR[ 239 ][ 207 ],
   alphaCSR[ 239 ][ 208 ],
   alphaCSR[ 239 ][ 209 ],
   alphaCSR[ 239 ][ 210 ],
   alphaCSR[ 239 ][ 211 ],
   alphaCSR[ 239 ][ 212 ],
   alphaCSR[ 239 ][ 213 ],
   alphaCSR[ 239 ][ 214 ],
   alphaCSR[ 239 ][ 215 ],
   alphaCSR[ 239 ][ 216 ],
   alphaCSR[ 239 ][ 217 ],
   alphaCSR[ 239 ][ 218 ],
   alphaCSR[ 239 ][ 219 ],
   alphaCSR[ 239 ][ 220 ],
   alphaCSR[ 239 ][ 221 ],
   alphaCSR[ 239 ][ 222 ],
   alphaCSR[ 239 ][ 223 ],
   alphaCSR[ 239 ][ 224 ],
   alphaCSR[ 239 ][ 225 ],
   alphaCSR[ 239 ][ 226 ],
   alphaCSR[ 239 ][ 227 ],
   alphaCSR[ 239 ][ 228 ],
   alphaCSR[ 239 ][ 229 ],
   alphaCSR[ 239 ][ 230 ],
   alphaCSR[ 239 ][ 231 ],
   alphaCSR[ 239 ][ 232 ],
   alphaCSR[ 239 ][ 233 ],
   alphaCSR[ 239 ][ 234 ],
   alphaCSR[ 239 ][ 235 ],
   alphaCSR[ 239 ][ 236 ],
   alphaCSR[ 239 ][ 237 ],
   alphaCSR[ 239 ][ 238 ],
   alphaCSR[ 239 ][ 239 ],
   alphaCSR[ 239 ][ 240 ],
   alphaCSR[ 239 ][ 241 ],
   alphaCSR[ 239 ][ 242 ],
   alphaCSR[ 239 ][ 243 ],
   alphaCSR[ 239 ][ 244 ],
   alphaCSR[ 239 ][ 245 ],
   alphaCSR[ 239 ][ 246 ],
   alphaCSR[ 239 ][ 247 ],
   alphaCSR[ 239 ][ 248 ],
   alphaCSR[ 239 ][ 249 ],
   alphaCSR[ 239 ][ 250 ],
   alphaCSR[ 239 ][ 251 ],
   alphaCSR[ 239 ][ 252 ],
   alphaCSR[ 239 ][ 253 ],
   alphaCSR[ 239 ][ 254 ],
   alphaCSR[ 239 ][ 255 ],
   alphaCSR[ 239 ][ 256 ],
   alphaCSR[ 239 ][ 257 ],
   alphaCSR[ 239 ][ 258 ],
   alphaCSR[ 239 ][ 259 ],
   alphaCSR[ 239 ][ 260 ],
   alphaCSR[ 239 ][ 261 ],
   alphaCSR[ 239 ][ 262 ],
   alphaCSR[ 239 ][ 263 ],
   alphaCSR[ 239 ][ 264 ],
   alphaCSR[ 239 ][ 265 ],
   alphaCSR[ 239 ][ 266 ],
   alphaCSR[ 239 ][ 267 ],
   alphaCSR[ 239 ][ 268 ],
   alphaCSR[ 239 ][ 269 ],
   alphaCSR[ 239 ][ 270 ],
   alphaCSR[ 239 ][ 271 ],
   alphaCSR[ 239 ][ 272 ],
   alphaCSR[ 239 ][ 273 ],
   alphaCSR[ 239 ][ 274 ],
   alphaCSR[ 239 ][ 275 ],
   alphaCSR[ 239 ][ 276 ],
   alphaCSR[ 239 ][ 277 ],
   alphaCSR[ 239 ][ 278 ],
   alphaCSR[ 239 ][ 279 ],
   alphaCSR[ 239 ][ 280 ],
   alphaCSR[ 239 ][ 281 ],
   alphaCSR[ 239 ][ 282 ],
   alphaCSR[ 239 ][ 283 ],
   alphaCSR[ 239 ][ 284 ],
   alphaCSR[ 239 ][ 285 ],
   alphaCSR[ 239 ][ 286 ],
   alphaCSR[ 239 ][ 287 ],
   alphaCSR[ 239 ][ 288 ],
   alphaCSR[ 239 ][ 289 ],
   alphaCSR[ 239 ][ 290 ],
   alphaCSR[ 239 ][ 291 ],
   alphaCSR[ 239 ][ 292 ],
   alphaCSR[ 239 ][ 293 ],
   alphaCSR[ 239 ][ 294 ],
   alphaCSR[ 239 ][ 295 ],
   alphaCSR[ 239 ][ 296 ],
   alphaCSR[ 239 ][ 297 ],
   alphaCSR[ 239 ][ 298 ],
   alphaCSR[ 239 ][ 299 ],
   alphaCSR[ 239 ][ 300 ],
   alphaCSR[ 239 ][ 301 ],
   alphaCSR[ 239 ][ 302 ],
   alphaCSR[ 239 ][ 303 ],
   alphaCSR[ 239 ][ 304 ],
   alphaCSR[ 239 ][ 305 ],
   alphaCSR[ 239 ][ 306 ],
   alphaCSR[ 239 ][ 307 ],
   alphaCSR[ 239 ][ 308 ],
   alphaCSR[ 239 ][ 309 ],
   alphaCSR[ 239 ][ 310 ],
   alphaCSR[ 239 ][ 311 ],
   alphaCSR[ 239 ][ 312 ],
   alphaCSR[ 239 ][ 313 ],
   alphaCSR[ 239 ][ 314 ],
   alphaCSR[ 239 ][ 315 ],
   alphaCSR[ 239 ][ 316 ],
   alphaCSR[ 239 ][ 317 ],
   alphaCSR[ 239 ][ 318 ],
   alphaCSR[ 239 ][ 319 ],
   alphaCSR[ 239 ][ 320 ],
   alphaCSR[ 239 ][ 321 ],
   alphaCSR[ 239 ][ 322 ],
   alphaCSR[ 239 ][ 323 ],
   alphaCSR[ 239 ][ 324 ],
   alphaCSR[ 239 ][ 325 ],
   alphaCSR[ 239 ][ 326 ],
   alphaCSR[ 239 ][ 327 ],
   alphaCSR[ 239 ][ 328 ],
   alphaCSR[ 239 ][ 329 ],
   alphaCSR[ 239 ][ 330 ],
   alphaCSR[ 239 ][ 331 ],
   alphaCSR[ 239 ][ 332 ],
   alphaCSR[ 239 ][ 333 ],
   alphaCSR[ 239 ][ 334 ],
   alphaCSR[ 239 ][ 335 ],
   alphaCSR[ 239 ][ 336 ],
   alphaCSR[ 239 ][ 337 ],
   alphaCSR[ 239 ][ 338 ],
   alphaCSR[ 239 ][ 339 ],
   alphaCSR[ 239 ][ 340 ],
   alphaCSR[ 239 ][ 341 ],
   alphaCSR[ 239 ][ 342 ],
   alphaCSR[ 239 ][ 343 ],
   alphaCSR[ 239 ][ 344 ],
   alphaCSR[ 239 ][ 345 ],
   alphaCSR[ 239 ][ 346 ],
   alphaCSR[ 239 ][ 347 ],
   alphaCSR[ 239 ][ 348 ],
   alphaCSR[ 239 ][ 349 ],
   alphaCSR[ 239 ][ 350 ],
   alphaCSR[ 239 ][ 351 ],
   alphaCSR[ 239 ][ 352 ],
   alphaCSR[ 239 ][ 353 ],
   alphaCSR[ 239 ][ 354 ],
   alphaCSR[ 239 ][ 355 ],
   alphaCSR[ 239 ][ 356 ],
   alphaCSR[ 239 ][ 357 ],
   alphaCSR[ 239 ][ 358 ],
   alphaCSR[ 239 ][ 359 ],
   alphaCSR[ 239 ][ 360 ],
   alphaCSR[ 239 ][ 361 ],
   alphaCSR[ 239 ][ 362 ],
   alphaCSR[ 239 ][ 363 ],
   alphaCSR[ 239 ][ 364 ],
   alphaCSR[ 239 ][ 365 ],
   alphaCSR[ 239 ][ 366 ],
   alphaCSR[ 239 ][ 367 ],
   alphaCSR[ 239 ][ 368 ],
   alphaCSR[ 239 ][ 369 ],
   alphaCSR[ 239 ][ 370 ],
   alphaCSR[ 239 ][ 371 ],
   alphaCSR[ 239 ][ 372 ],
   alphaCSR[ 239 ][ 373 ],
   alphaCSR[ 239 ][ 374 ],
   alphaCSR[ 239 ][ 375 ],
   alphaCSR[ 239 ][ 376 ],
   alphaCSR[ 239 ][ 377 ],
   alphaCSR[ 239 ][ 378 ],
   alphaCSR[ 239 ][ 379 ],
   alphaCSR[ 239 ][ 380 ],
   alphaCSR[ 239 ][ 381 ],
   alphaCSR[ 239 ][ 382 ],
   alphaCSR[ 239 ][ 383 ],
   alphaCSR[ 240 ][ 0 ],
   alphaCSR[ 240 ][ 1 ],
   alphaCSR[ 240 ][ 2 ],
   alphaCSR[ 240 ][ 3 ],
   alphaCSR[ 240 ][ 4 ],
   alphaCSR[ 240 ][ 5 ],
   alphaCSR[ 240 ][ 6 ],
   alphaCSR[ 240 ][ 7 ],
   alphaCSR[ 240 ][ 8 ],
   alphaCSR[ 240 ][ 9 ],
   alphaCSR[ 240 ][ 10 ],
   alphaCSR[ 240 ][ 11 ],
   alphaCSR[ 240 ][ 12 ],
   alphaCSR[ 240 ][ 13 ],
   alphaCSR[ 240 ][ 14 ],
   alphaCSR[ 240 ][ 15 ],
   alphaCSR[ 240 ][ 16 ],
   alphaCSR[ 240 ][ 17 ],
   alphaCSR[ 240 ][ 18 ],
   alphaCSR[ 240 ][ 19 ],
   alphaCSR[ 240 ][ 20 ],
   alphaCSR[ 240 ][ 21 ],
   alphaCSR[ 240 ][ 22 ],
   alphaCSR[ 240 ][ 23 ],
   alphaCSR[ 240 ][ 24 ],
   alphaCSR[ 240 ][ 25 ],
   alphaCSR[ 240 ][ 26 ],
   alphaCSR[ 240 ][ 27 ],
   alphaCSR[ 240 ][ 28 ],
   alphaCSR[ 240 ][ 29 ],
   alphaCSR[ 240 ][ 30 ],
   alphaCSR[ 240 ][ 31 ],
   alphaCSR[ 240 ][ 32 ],
   alphaCSR[ 240 ][ 33 ],
   alphaCSR[ 240 ][ 34 ],
   alphaCSR[ 240 ][ 35 ],
   alphaCSR[ 240 ][ 36 ],
   alphaCSR[ 240 ][ 37 ],
   alphaCSR[ 240 ][ 38 ],
   alphaCSR[ 240 ][ 39 ],
   alphaCSR[ 240 ][ 40 ],
   alphaCSR[ 240 ][ 41 ],
   alphaCSR[ 240 ][ 42 ],
   alphaCSR[ 240 ][ 43 ],
   alphaCSR[ 240 ][ 44 ],
   alphaCSR[ 240 ][ 45 ],
   alphaCSR[ 240 ][ 46 ],
   alphaCSR[ 240 ][ 47 ],
   alphaCSR[ 240 ][ 48 ],
   alphaCSR[ 240 ][ 49 ],
   alphaCSR[ 240 ][ 50 ],
   alphaCSR[ 240 ][ 51 ],
   alphaCSR[ 240 ][ 52 ],
   alphaCSR[ 240 ][ 53 ],
   alphaCSR[ 240 ][ 54 ],
   alphaCSR[ 240 ][ 55 ],
   alphaCSR[ 240 ][ 56 ],
   alphaCSR[ 240 ][ 57 ],
   alphaCSR[ 240 ][ 58 ],
   alphaCSR[ 240 ][ 59 ],
   alphaCSR[ 240 ][ 60 ],
   alphaCSR[ 240 ][ 61 ],
   alphaCSR[ 240 ][ 62 ],
   alphaCSR[ 240 ][ 63 ],
   alphaCSR[ 240 ][ 64 ],
   alphaCSR[ 240 ][ 65 ],
   alphaCSR[ 240 ][ 66 ],
   alphaCSR[ 240 ][ 67 ],
   alphaCSR[ 240 ][ 68 ],
   alphaCSR[ 240 ][ 69 ],
   alphaCSR[ 240 ][ 70 ],
   alphaCSR[ 240 ][ 71 ],
   alphaCSR[ 240 ][ 72 ],
   alphaCSR[ 240 ][ 73 ],
   alphaCSR[ 240 ][ 74 ],
   alphaCSR[ 240 ][ 75 ],
   alphaCSR[ 240 ][ 76 ],
   alphaCSR[ 240 ][ 77 ],
   alphaCSR[ 240 ][ 78 ],
   alphaCSR[ 240 ][ 79 ],
   alphaCSR[ 240 ][ 80 ],
   alphaCSR[ 240 ][ 81 ],
   alphaCSR[ 240 ][ 82 ],
   alphaCSR[ 240 ][ 83 ],
   alphaCSR[ 240 ][ 84 ],
   alphaCSR[ 240 ][ 85 ],
   alphaCSR[ 240 ][ 86 ],
   alphaCSR[ 240 ][ 87 ],
   alphaCSR[ 240 ][ 88 ],
   alphaCSR[ 240 ][ 89 ],
   alphaCSR[ 240 ][ 90 ],
   alphaCSR[ 240 ][ 91 ],
   alphaCSR[ 240 ][ 92 ],
   alphaCSR[ 240 ][ 93 ],
   alphaCSR[ 240 ][ 94 ],
   alphaCSR[ 240 ][ 95 ],
   alphaCSR[ 240 ][ 96 ],
   alphaCSR[ 240 ][ 97 ],
   alphaCSR[ 240 ][ 98 ],
   alphaCSR[ 240 ][ 99 ],
   alphaCSR[ 240 ][ 100 ],
   alphaCSR[ 240 ][ 101 ],
   alphaCSR[ 240 ][ 102 ],
   alphaCSR[ 240 ][ 103 ],
   alphaCSR[ 240 ][ 104 ],
   alphaCSR[ 240 ][ 105 ],
   alphaCSR[ 240 ][ 106 ],
   alphaCSR[ 240 ][ 107 ],
   alphaCSR[ 240 ][ 108 ],
   alphaCSR[ 240 ][ 109 ],
   alphaCSR[ 240 ][ 110 ],
   alphaCSR[ 240 ][ 111 ],
   alphaCSR[ 240 ][ 112 ],
   alphaCSR[ 240 ][ 113 ],
   alphaCSR[ 240 ][ 114 ],
   alphaCSR[ 240 ][ 115 ],
   alphaCSR[ 240 ][ 116 ],
   alphaCSR[ 240 ][ 117 ],
   alphaCSR[ 240 ][ 118 ],
   alphaCSR[ 240 ][ 119 ],
   alphaCSR[ 240 ][ 120 ],
   alphaCSR[ 240 ][ 121 ],
   alphaCSR[ 240 ][ 122 ],
   alphaCSR[ 240 ][ 123 ],
   alphaCSR[ 240 ][ 124 ],
   alphaCSR[ 240 ][ 125 ],
   alphaCSR[ 240 ][ 126 ],
   alphaCSR[ 240 ][ 127 ],
   alphaCSR[ 240 ][ 128 ],
   alphaCSR[ 240 ][ 129 ],
   alphaCSR[ 240 ][ 130 ],
   alphaCSR[ 240 ][ 131 ],
   alphaCSR[ 240 ][ 132 ],
   alphaCSR[ 240 ][ 133 ],
   alphaCSR[ 240 ][ 134 ],
   alphaCSR[ 240 ][ 135 ],
   alphaCSR[ 240 ][ 136 ],
   alphaCSR[ 240 ][ 137 ],
   alphaCSR[ 240 ][ 138 ],
   alphaCSR[ 240 ][ 139 ],
   alphaCSR[ 240 ][ 140 ],
   alphaCSR[ 240 ][ 141 ],
   alphaCSR[ 240 ][ 142 ],
   alphaCSR[ 240 ][ 143 ],
   alphaCSR[ 240 ][ 144 ],
   alphaCSR[ 240 ][ 145 ],
   alphaCSR[ 240 ][ 146 ],
   alphaCSR[ 240 ][ 147 ],
   alphaCSR[ 240 ][ 148 ],
   alphaCSR[ 240 ][ 149 ],
   alphaCSR[ 240 ][ 150 ],
   alphaCSR[ 240 ][ 151 ],
   alphaCSR[ 240 ][ 152 ],
   alphaCSR[ 240 ][ 153 ],
   alphaCSR[ 240 ][ 154 ],
   alphaCSR[ 240 ][ 155 ],
   alphaCSR[ 240 ][ 156 ],
   alphaCSR[ 240 ][ 157 ],
   alphaCSR[ 240 ][ 158 ],
   alphaCSR[ 240 ][ 159 ],
   alphaCSR[ 240 ][ 160 ],
   alphaCSR[ 240 ][ 161 ],
   alphaCSR[ 240 ][ 162 ],
   alphaCSR[ 240 ][ 163 ],
   alphaCSR[ 240 ][ 164 ],
   alphaCSR[ 240 ][ 165 ],
   alphaCSR[ 240 ][ 166 ],
   alphaCSR[ 240 ][ 167 ],
   alphaCSR[ 240 ][ 168 ],
   alphaCSR[ 240 ][ 169 ],
   alphaCSR[ 240 ][ 170 ],
   alphaCSR[ 240 ][ 171 ],
   alphaCSR[ 240 ][ 172 ],
   alphaCSR[ 240 ][ 173 ],
   alphaCSR[ 240 ][ 174 ],
   alphaCSR[ 240 ][ 175 ],
   alphaCSR[ 240 ][ 176 ],
   alphaCSR[ 240 ][ 177 ],
   alphaCSR[ 240 ][ 178 ],
   alphaCSR[ 240 ][ 179 ],
   alphaCSR[ 240 ][ 180 ],
   alphaCSR[ 240 ][ 181 ],
   alphaCSR[ 240 ][ 182 ],
   alphaCSR[ 240 ][ 183 ],
   alphaCSR[ 240 ][ 184 ],
   alphaCSR[ 240 ][ 185 ],
   alphaCSR[ 240 ][ 186 ],
   alphaCSR[ 240 ][ 187 ],
   alphaCSR[ 240 ][ 188 ],
   alphaCSR[ 240 ][ 189 ],
   alphaCSR[ 240 ][ 190 ],
   alphaCSR[ 240 ][ 191 ],
   alphaCSR[ 240 ][ 192 ],
   alphaCSR[ 240 ][ 193 ],
   alphaCSR[ 240 ][ 194 ],
   alphaCSR[ 240 ][ 195 ],
   alphaCSR[ 240 ][ 196 ],
   alphaCSR[ 240 ][ 197 ],
   alphaCSR[ 240 ][ 198 ],
   alphaCSR[ 240 ][ 199 ],
   alphaCSR[ 240 ][ 200 ],
   alphaCSR[ 240 ][ 201 ],
   alphaCSR[ 240 ][ 202 ],
   alphaCSR[ 240 ][ 203 ],
   alphaCSR[ 240 ][ 204 ],
   alphaCSR[ 240 ][ 205 ],
   alphaCSR[ 240 ][ 206 ],
   alphaCSR[ 240 ][ 207 ],
   alphaCSR[ 240 ][ 208 ],
   alphaCSR[ 240 ][ 209 ],
   alphaCSR[ 240 ][ 210 ],
   alphaCSR[ 240 ][ 211 ],
   alphaCSR[ 240 ][ 212 ],
   alphaCSR[ 240 ][ 213 ],
   alphaCSR[ 240 ][ 214 ],
   alphaCSR[ 240 ][ 215 ],
   alphaCSR[ 240 ][ 216 ],
   alphaCSR[ 240 ][ 217 ],
   alphaCSR[ 240 ][ 218 ],
   alphaCSR[ 240 ][ 219 ],
   alphaCSR[ 240 ][ 220 ],
   alphaCSR[ 240 ][ 221 ],
   alphaCSR[ 240 ][ 222 ],
   alphaCSR[ 240 ][ 223 ],
   alphaCSR[ 240 ][ 224 ],
   alphaCSR[ 240 ][ 225 ],
   alphaCSR[ 240 ][ 226 ],
   alphaCSR[ 240 ][ 227 ],
   alphaCSR[ 240 ][ 228 ],
   alphaCSR[ 240 ][ 229 ],
   alphaCSR[ 240 ][ 230 ],
   alphaCSR[ 240 ][ 231 ],
   alphaCSR[ 240 ][ 232 ],
   alphaCSR[ 240 ][ 233 ],
   alphaCSR[ 240 ][ 234 ],
   alphaCSR[ 240 ][ 235 ],
   alphaCSR[ 240 ][ 236 ],
   alphaCSR[ 240 ][ 237 ],
   alphaCSR[ 240 ][ 238 ],
   alphaCSR[ 240 ][ 239 ],
   alphaCSR[ 240 ][ 240 ],
   alphaCSR[ 240 ][ 241 ],
   alphaCSR[ 240 ][ 242 ],
   alphaCSR[ 240 ][ 243 ],
   alphaCSR[ 240 ][ 244 ],
   alphaCSR[ 240 ][ 245 ],
   alphaCSR[ 240 ][ 246 ],
   alphaCSR[ 240 ][ 247 ],
   alphaCSR[ 240 ][ 248 ],
   alphaCSR[ 240 ][ 249 ],
   alphaCSR[ 240 ][ 250 ],
   alphaCSR[ 240 ][ 251 ],
   alphaCSR[ 240 ][ 252 ],
   alphaCSR[ 240 ][ 253 ],
   alphaCSR[ 240 ][ 254 ],
   alphaCSR[ 240 ][ 255 ],
   alphaCSR[ 240 ][ 256 ],
   alphaCSR[ 240 ][ 257 ],
   alphaCSR[ 240 ][ 258 ],
   alphaCSR[ 240 ][ 259 ],
   alphaCSR[ 240 ][ 260 ],
   alphaCSR[ 240 ][ 261 ],
   alphaCSR[ 240 ][ 262 ],
   alphaCSR[ 240 ][ 263 ],
   alphaCSR[ 240 ][ 264 ],
   alphaCSR[ 240 ][ 265 ],
   alphaCSR[ 240 ][ 266 ],
   alphaCSR[ 240 ][ 267 ],
   alphaCSR[ 240 ][ 268 ],
   alphaCSR[ 240 ][ 269 ],
   alphaCSR[ 240 ][ 270 ],
   alphaCSR[ 240 ][ 271 ],
   alphaCSR[ 240 ][ 272 ],
   alphaCSR[ 240 ][ 273 ],
   alphaCSR[ 240 ][ 274 ],
   alphaCSR[ 240 ][ 275 ],
   alphaCSR[ 240 ][ 276 ],
   alphaCSR[ 240 ][ 277 ],
   alphaCSR[ 240 ][ 278 ],
   alphaCSR[ 240 ][ 279 ],
   alphaCSR[ 240 ][ 280 ],
   alphaCSR[ 240 ][ 281 ],
   alphaCSR[ 240 ][ 282 ],
   alphaCSR[ 240 ][ 283 ],
   alphaCSR[ 240 ][ 284 ],
   alphaCSR[ 240 ][ 285 ],
   alphaCSR[ 240 ][ 286 ],
   alphaCSR[ 240 ][ 287 ],
   alphaCSR[ 240 ][ 288 ],
   alphaCSR[ 240 ][ 289 ],
   alphaCSR[ 240 ][ 290 ],
   alphaCSR[ 240 ][ 291 ],
   alphaCSR[ 240 ][ 292 ],
   alphaCSR[ 240 ][ 293 ],
   alphaCSR[ 240 ][ 294 ],
   alphaCSR[ 240 ][ 295 ],
   alphaCSR[ 240 ][ 296 ],
   alphaCSR[ 240 ][ 297 ],
   alphaCSR[ 240 ][ 298 ],
   alphaCSR[ 240 ][ 299 ],
   alphaCSR[ 240 ][ 300 ],
   alphaCSR[ 240 ][ 301 ],
   alphaCSR[ 240 ][ 302 ],
   alphaCSR[ 240 ][ 303 ],
   alphaCSR[ 240 ][ 304 ],
   alphaCSR[ 240 ][ 305 ],
   alphaCSR[ 240 ][ 306 ],
   alphaCSR[ 240 ][ 307 ],
   alphaCSR[ 240 ][ 308 ],
   alphaCSR[ 240 ][ 309 ],
   alphaCSR[ 240 ][ 310 ],
   alphaCSR[ 240 ][ 311 ],
   alphaCSR[ 240 ][ 312 ],
   alphaCSR[ 240 ][ 313 ],
   alphaCSR[ 240 ][ 314 ],
   alphaCSR[ 240 ][ 315 ],
   alphaCSR[ 240 ][ 316 ],
   alphaCSR[ 240 ][ 317 ],
   alphaCSR[ 240 ][ 318 ],
   alphaCSR[ 240 ][ 319 ],
   alphaCSR[ 240 ][ 320 ],
   alphaCSR[ 240 ][ 321 ],
   alphaCSR[ 240 ][ 322 ],
   alphaCSR[ 240 ][ 323 ],
   alphaCSR[ 240 ][ 324 ],
   alphaCSR[ 240 ][ 325 ],
   alphaCSR[ 240 ][ 326 ],
   alphaCSR[ 240 ][ 327 ],
   alphaCSR[ 240 ][ 328 ],
   alphaCSR[ 240 ][ 329 ],
   alphaCSR[ 240 ][ 330 ],
   alphaCSR[ 240 ][ 331 ],
   alphaCSR[ 240 ][ 332 ],
   alphaCSR[ 240 ][ 333 ],
   alphaCSR[ 240 ][ 334 ],
   alphaCSR[ 240 ][ 335 ],
   alphaCSR[ 240 ][ 336 ],
   alphaCSR[ 240 ][ 337 ],
   alphaCSR[ 240 ][ 338 ],
   alphaCSR[ 240 ][ 339 ],
   alphaCSR[ 240 ][ 340 ],
   alphaCSR[ 240 ][ 341 ],
   alphaCSR[ 240 ][ 342 ],
   alphaCSR[ 240 ][ 343 ],
   alphaCSR[ 240 ][ 344 ],
   alphaCSR[ 240 ][ 345 ],
   alphaCSR[ 240 ][ 346 ],
   alphaCSR[ 240 ][ 347 ],
   alphaCSR[ 240 ][ 348 ],
   alphaCSR[ 240 ][ 349 ],
   alphaCSR[ 240 ][ 350 ],
   alphaCSR[ 240 ][ 351 ],
   alphaCSR[ 240 ][ 352 ],
   alphaCSR[ 240 ][ 353 ],
   alphaCSR[ 240 ][ 354 ],
   alphaCSR[ 240 ][ 355 ],
   alphaCSR[ 240 ][ 356 ],
   alphaCSR[ 240 ][ 357 ],
   alphaCSR[ 240 ][ 358 ],
   alphaCSR[ 240 ][ 359 ],
   alphaCSR[ 240 ][ 360 ],
   alphaCSR[ 240 ][ 361 ],
   alphaCSR[ 240 ][ 362 ],
   alphaCSR[ 240 ][ 363 ],
   alphaCSR[ 240 ][ 364 ],
   alphaCSR[ 240 ][ 365 ],
   alphaCSR[ 240 ][ 366 ],
   alphaCSR[ 240 ][ 367 ],
   alphaCSR[ 240 ][ 368 ],
   alphaCSR[ 240 ][ 369 ],
   alphaCSR[ 240 ][ 370 ],
   alphaCSR[ 240 ][ 371 ],
   alphaCSR[ 240 ][ 372 ],
   alphaCSR[ 240 ][ 373 ],
   alphaCSR[ 240 ][ 374 ],
   alphaCSR[ 240 ][ 375 ],
   alphaCSR[ 240 ][ 376 ],
   alphaCSR[ 240 ][ 377 ],
   alphaCSR[ 240 ][ 378 ],
   alphaCSR[ 240 ][ 379 ],
   alphaCSR[ 240 ][ 380 ],
   alphaCSR[ 240 ][ 381 ],
   alphaCSR[ 240 ][ 382 ],
   alphaCSR[ 240 ][ 383 ],
   alphaCSR[ 241 ][ 0 ],
   alphaCSR[ 241 ][ 1 ],
   alphaCSR[ 241 ][ 2 ],
   alphaCSR[ 241 ][ 3 ],
   alphaCSR[ 241 ][ 4 ],
   alphaCSR[ 241 ][ 5 ],
   alphaCSR[ 241 ][ 6 ],
   alphaCSR[ 241 ][ 7 ],
   alphaCSR[ 241 ][ 8 ],
   alphaCSR[ 241 ][ 9 ],
   alphaCSR[ 241 ][ 10 ],
   alphaCSR[ 241 ][ 11 ],
   alphaCSR[ 241 ][ 12 ],
   alphaCSR[ 241 ][ 13 ],
   alphaCSR[ 241 ][ 14 ],
   alphaCSR[ 241 ][ 15 ],
   alphaCSR[ 241 ][ 16 ],
   alphaCSR[ 241 ][ 17 ],
   alphaCSR[ 241 ][ 18 ],
   alphaCSR[ 241 ][ 19 ],
   alphaCSR[ 241 ][ 20 ],
   alphaCSR[ 241 ][ 21 ],
   alphaCSR[ 241 ][ 22 ],
   alphaCSR[ 241 ][ 23 ],
   alphaCSR[ 241 ][ 24 ],
   alphaCSR[ 241 ][ 25 ],
   alphaCSR[ 241 ][ 26 ],
   alphaCSR[ 241 ][ 27 ],
   alphaCSR[ 241 ][ 28 ],
   alphaCSR[ 241 ][ 29 ],
   alphaCSR[ 241 ][ 30 ],
   alphaCSR[ 241 ][ 31 ],
   alphaCSR[ 241 ][ 32 ],
   alphaCSR[ 241 ][ 33 ],
   alphaCSR[ 241 ][ 34 ],
   alphaCSR[ 241 ][ 35 ],
   alphaCSR[ 241 ][ 36 ],
   alphaCSR[ 241 ][ 37 ],
   alphaCSR[ 241 ][ 38 ],
   alphaCSR[ 241 ][ 39 ],
   alphaCSR[ 241 ][ 40 ],
   alphaCSR[ 241 ][ 41 ],
   alphaCSR[ 241 ][ 42 ],
   alphaCSR[ 241 ][ 43 ],
   alphaCSR[ 241 ][ 44 ],
   alphaCSR[ 241 ][ 45 ],
   alphaCSR[ 241 ][ 46 ],
   alphaCSR[ 241 ][ 47 ],
   alphaCSR[ 241 ][ 48 ],
   alphaCSR[ 241 ][ 49 ],
   alphaCSR[ 241 ][ 50 ],
   alphaCSR[ 241 ][ 51 ],
   alphaCSR[ 241 ][ 52 ],
   alphaCSR[ 241 ][ 53 ],
   alphaCSR[ 241 ][ 54 ],
   alphaCSR[ 241 ][ 55 ],
   alphaCSR[ 241 ][ 56 ],
   alphaCSR[ 241 ][ 57 ],
   alphaCSR[ 241 ][ 58 ],
   alphaCSR[ 241 ][ 59 ],
   alphaCSR[ 241 ][ 60 ],
   alphaCSR[ 241 ][ 61 ],
   alphaCSR[ 241 ][ 62 ],
   alphaCSR[ 241 ][ 63 ],
   alphaCSR[ 241 ][ 64 ],
   alphaCSR[ 241 ][ 65 ],
   alphaCSR[ 241 ][ 66 ],
   alphaCSR[ 241 ][ 67 ],
   alphaCSR[ 241 ][ 68 ],
   alphaCSR[ 241 ][ 69 ],
   alphaCSR[ 241 ][ 70 ],
   alphaCSR[ 241 ][ 71 ],
   alphaCSR[ 241 ][ 72 ],
   alphaCSR[ 241 ][ 73 ],
   alphaCSR[ 241 ][ 74 ],
   alphaCSR[ 241 ][ 75 ],
   alphaCSR[ 241 ][ 76 ],
   alphaCSR[ 241 ][ 77 ],
   alphaCSR[ 241 ][ 78 ],
   alphaCSR[ 241 ][ 79 ],
   alphaCSR[ 241 ][ 80 ],
   alphaCSR[ 241 ][ 81 ],
   alphaCSR[ 241 ][ 82 ],
   alphaCSR[ 241 ][ 83 ],
   alphaCSR[ 241 ][ 84 ],
   alphaCSR[ 241 ][ 85 ],
   alphaCSR[ 241 ][ 86 ],
   alphaCSR[ 241 ][ 87 ],
   alphaCSR[ 241 ][ 88 ],
   alphaCSR[ 241 ][ 89 ],
   alphaCSR[ 241 ][ 90 ],
   alphaCSR[ 241 ][ 91 ],
   alphaCSR[ 241 ][ 92 ],
   alphaCSR[ 241 ][ 93 ],
   alphaCSR[ 241 ][ 94 ],
   alphaCSR[ 241 ][ 95 ],
   alphaCSR[ 241 ][ 96 ],
   alphaCSR[ 241 ][ 97 ],
   alphaCSR[ 241 ][ 98 ],
   alphaCSR[ 241 ][ 99 ],
   alphaCSR[ 241 ][ 100 ],
   alphaCSR[ 241 ][ 101 ],
   alphaCSR[ 241 ][ 102 ],
   alphaCSR[ 241 ][ 103 ],
   alphaCSR[ 241 ][ 104 ],
   alphaCSR[ 241 ][ 105 ],
   alphaCSR[ 241 ][ 106 ],
   alphaCSR[ 241 ][ 107 ],
   alphaCSR[ 241 ][ 108 ],
   alphaCSR[ 241 ][ 109 ],
   alphaCSR[ 241 ][ 110 ],
   alphaCSR[ 241 ][ 111 ],
   alphaCSR[ 241 ][ 112 ],
   alphaCSR[ 241 ][ 113 ],
   alphaCSR[ 241 ][ 114 ],
   alphaCSR[ 241 ][ 115 ],
   alphaCSR[ 241 ][ 116 ],
   alphaCSR[ 241 ][ 117 ],
   alphaCSR[ 241 ][ 118 ],
   alphaCSR[ 241 ][ 119 ],
   alphaCSR[ 241 ][ 120 ],
   alphaCSR[ 241 ][ 121 ],
   alphaCSR[ 241 ][ 122 ],
   alphaCSR[ 241 ][ 123 ],
   alphaCSR[ 241 ][ 124 ],
   alphaCSR[ 241 ][ 125 ],
   alphaCSR[ 241 ][ 126 ],
   alphaCSR[ 241 ][ 127 ],
   alphaCSR[ 241 ][ 128 ],
   alphaCSR[ 241 ][ 129 ],
   alphaCSR[ 241 ][ 130 ],
   alphaCSR[ 241 ][ 131 ],
   alphaCSR[ 241 ][ 132 ],
   alphaCSR[ 241 ][ 133 ],
   alphaCSR[ 241 ][ 134 ],
   alphaCSR[ 241 ][ 135 ],
   alphaCSR[ 241 ][ 136 ],
   alphaCSR[ 241 ][ 137 ],
   alphaCSR[ 241 ][ 138 ],
   alphaCSR[ 241 ][ 139 ],
   alphaCSR[ 241 ][ 140 ],
   alphaCSR[ 241 ][ 141 ],
   alphaCSR[ 241 ][ 142 ],
   alphaCSR[ 241 ][ 143 ],
   alphaCSR[ 241 ][ 144 ],
   alphaCSR[ 241 ][ 145 ],
   alphaCSR[ 241 ][ 146 ],
   alphaCSR[ 241 ][ 147 ],
   alphaCSR[ 241 ][ 148 ],
   alphaCSR[ 241 ][ 149 ],
   alphaCSR[ 241 ][ 150 ],
   alphaCSR[ 241 ][ 151 ],
   alphaCSR[ 241 ][ 152 ],
   alphaCSR[ 241 ][ 153 ],
   alphaCSR[ 241 ][ 154 ],
   alphaCSR[ 241 ][ 155 ],
   alphaCSR[ 241 ][ 156 ],
   alphaCSR[ 241 ][ 157 ],
   alphaCSR[ 241 ][ 158 ],
   alphaCSR[ 241 ][ 159 ],
   alphaCSR[ 241 ][ 160 ],
   alphaCSR[ 241 ][ 161 ],
   alphaCSR[ 241 ][ 162 ],
   alphaCSR[ 241 ][ 163 ],
   alphaCSR[ 241 ][ 164 ],
   alphaCSR[ 241 ][ 165 ],
   alphaCSR[ 241 ][ 166 ],
   alphaCSR[ 241 ][ 167 ],
   alphaCSR[ 241 ][ 168 ],
   alphaCSR[ 241 ][ 169 ],
   alphaCSR[ 241 ][ 170 ],
   alphaCSR[ 241 ][ 171 ],
   alphaCSR[ 241 ][ 172 ],
   alphaCSR[ 241 ][ 173 ],
   alphaCSR[ 241 ][ 174 ],
   alphaCSR[ 241 ][ 175 ],
   alphaCSR[ 241 ][ 176 ],
   alphaCSR[ 241 ][ 177 ],
   alphaCSR[ 241 ][ 178 ],
   alphaCSR[ 241 ][ 179 ],
   alphaCSR[ 241 ][ 180 ],
   alphaCSR[ 241 ][ 181 ],
   alphaCSR[ 241 ][ 182 ],
   alphaCSR[ 241 ][ 183 ],
   alphaCSR[ 241 ][ 184 ],
   alphaCSR[ 241 ][ 185 ],
   alphaCSR[ 241 ][ 186 ],
   alphaCSR[ 241 ][ 187 ],
   alphaCSR[ 241 ][ 188 ],
   alphaCSR[ 241 ][ 189 ],
   alphaCSR[ 241 ][ 190 ],
   alphaCSR[ 241 ][ 191 ],
   alphaCSR[ 241 ][ 192 ],
   alphaCSR[ 241 ][ 193 ],
   alphaCSR[ 241 ][ 194 ],
   alphaCSR[ 241 ][ 195 ],
   alphaCSR[ 241 ][ 196 ],
   alphaCSR[ 241 ][ 197 ],
   alphaCSR[ 241 ][ 198 ],
   alphaCSR[ 241 ][ 199 ],
   alphaCSR[ 241 ][ 200 ],
   alphaCSR[ 241 ][ 201 ],
   alphaCSR[ 241 ][ 202 ],
   alphaCSR[ 241 ][ 203 ],
   alphaCSR[ 241 ][ 204 ],
   alphaCSR[ 241 ][ 205 ],
   alphaCSR[ 241 ][ 206 ],
   alphaCSR[ 241 ][ 207 ],
   alphaCSR[ 241 ][ 208 ],
   alphaCSR[ 241 ][ 209 ],
   alphaCSR[ 241 ][ 210 ],
   alphaCSR[ 241 ][ 211 ],
   alphaCSR[ 241 ][ 212 ],
   alphaCSR[ 241 ][ 213 ],
   alphaCSR[ 241 ][ 214 ],
   alphaCSR[ 241 ][ 215 ],
   alphaCSR[ 241 ][ 216 ],
   alphaCSR[ 241 ][ 217 ],
   alphaCSR[ 241 ][ 218 ],
   alphaCSR[ 241 ][ 219 ],
   alphaCSR[ 241 ][ 220 ],
   alphaCSR[ 241 ][ 221 ],
   alphaCSR[ 241 ][ 222 ],
   alphaCSR[ 241 ][ 223 ],
   alphaCSR[ 241 ][ 224 ],
   alphaCSR[ 241 ][ 225 ],
   alphaCSR[ 241 ][ 226 ],
   alphaCSR[ 241 ][ 227 ],
   alphaCSR[ 241 ][ 228 ],
   alphaCSR[ 241 ][ 229 ],
   alphaCSR[ 241 ][ 230 ],
   alphaCSR[ 241 ][ 231 ],
   alphaCSR[ 241 ][ 232 ],
   alphaCSR[ 241 ][ 233 ],
   alphaCSR[ 241 ][ 234 ],
   alphaCSR[ 241 ][ 235 ],
   alphaCSR[ 241 ][ 236 ],
   alphaCSR[ 241 ][ 237 ],
   alphaCSR[ 241 ][ 238 ],
   alphaCSR[ 241 ][ 239 ],
   alphaCSR[ 241 ][ 240 ],
   alphaCSR[ 241 ][ 241 ],
   alphaCSR[ 241 ][ 242 ],
   alphaCSR[ 241 ][ 243 ],
   alphaCSR[ 241 ][ 244 ],
   alphaCSR[ 241 ][ 245 ],
   alphaCSR[ 241 ][ 246 ],
   alphaCSR[ 241 ][ 247 ],
   alphaCSR[ 241 ][ 248 ],
   alphaCSR[ 241 ][ 249 ],
   alphaCSR[ 241 ][ 250 ],
   alphaCSR[ 241 ][ 251 ],
   alphaCSR[ 241 ][ 252 ],
   alphaCSR[ 241 ][ 253 ],
   alphaCSR[ 241 ][ 254 ],
   alphaCSR[ 241 ][ 255 ],
   alphaCSR[ 241 ][ 256 ],
   alphaCSR[ 241 ][ 257 ],
   alphaCSR[ 241 ][ 258 ],
   alphaCSR[ 241 ][ 259 ],
   alphaCSR[ 241 ][ 260 ],
   alphaCSR[ 241 ][ 261 ],
   alphaCSR[ 241 ][ 262 ],
   alphaCSR[ 241 ][ 263 ],
   alphaCSR[ 241 ][ 264 ],
   alphaCSR[ 241 ][ 265 ],
   alphaCSR[ 241 ][ 266 ],
   alphaCSR[ 241 ][ 267 ],
   alphaCSR[ 241 ][ 268 ],
   alphaCSR[ 241 ][ 269 ],
   alphaCSR[ 241 ][ 270 ],
   alphaCSR[ 241 ][ 271 ],
   alphaCSR[ 241 ][ 272 ],
   alphaCSR[ 241 ][ 273 ],
   alphaCSR[ 241 ][ 274 ],
   alphaCSR[ 241 ][ 275 ],
   alphaCSR[ 241 ][ 276 ],
   alphaCSR[ 241 ][ 277 ],
   alphaCSR[ 241 ][ 278 ],
   alphaCSR[ 241 ][ 279 ],
   alphaCSR[ 241 ][ 280 ],
   alphaCSR[ 241 ][ 281 ],
   alphaCSR[ 241 ][ 282 ],
   alphaCSR[ 241 ][ 283 ],
   alphaCSR[ 241 ][ 284 ],
   alphaCSR[ 241 ][ 285 ],
   alphaCSR[ 241 ][ 286 ],
   alphaCSR[ 241 ][ 287 ],
   alphaCSR[ 241 ][ 288 ],
   alphaCSR[ 241 ][ 289 ],
   alphaCSR[ 241 ][ 290 ],
   alphaCSR[ 241 ][ 291 ],
   alphaCSR[ 241 ][ 292 ],
   alphaCSR[ 241 ][ 293 ],
   alphaCSR[ 241 ][ 294 ],
   alphaCSR[ 241 ][ 295 ],
   alphaCSR[ 241 ][ 296 ],
   alphaCSR[ 241 ][ 297 ],
   alphaCSR[ 241 ][ 298 ],
   alphaCSR[ 241 ][ 299 ],
   alphaCSR[ 241 ][ 300 ],
   alphaCSR[ 241 ][ 301 ],
   alphaCSR[ 241 ][ 302 ],
   alphaCSR[ 241 ][ 303 ],
   alphaCSR[ 241 ][ 304 ],
   alphaCSR[ 241 ][ 305 ],
   alphaCSR[ 241 ][ 306 ],
   alphaCSR[ 241 ][ 307 ],
   alphaCSR[ 241 ][ 308 ],
   alphaCSR[ 241 ][ 309 ],
   alphaCSR[ 241 ][ 310 ],
   alphaCSR[ 241 ][ 311 ],
   alphaCSR[ 241 ][ 312 ],
   alphaCSR[ 241 ][ 313 ],
   alphaCSR[ 241 ][ 314 ],
   alphaCSR[ 241 ][ 315 ],
   alphaCSR[ 241 ][ 316 ],
   alphaCSR[ 241 ][ 317 ],
   alphaCSR[ 241 ][ 318 ],
   alphaCSR[ 241 ][ 319 ],
   alphaCSR[ 241 ][ 320 ],
   alphaCSR[ 241 ][ 321 ],
   alphaCSR[ 241 ][ 322 ],
   alphaCSR[ 241 ][ 323 ],
   alphaCSR[ 241 ][ 324 ],
   alphaCSR[ 241 ][ 325 ],
   alphaCSR[ 241 ][ 326 ],
   alphaCSR[ 241 ][ 327 ],
   alphaCSR[ 241 ][ 328 ],
   alphaCSR[ 241 ][ 329 ],
   alphaCSR[ 241 ][ 330 ],
   alphaCSR[ 241 ][ 331 ],
   alphaCSR[ 241 ][ 332 ],
   alphaCSR[ 241 ][ 333 ],
   alphaCSR[ 241 ][ 334 ],
   alphaCSR[ 241 ][ 335 ],
   alphaCSR[ 241 ][ 336 ],
   alphaCSR[ 241 ][ 337 ],
   alphaCSR[ 241 ][ 338 ],
   alphaCSR[ 241 ][ 339 ],
   alphaCSR[ 241 ][ 340 ],
   alphaCSR[ 241 ][ 341 ],
   alphaCSR[ 241 ][ 342 ],
   alphaCSR[ 241 ][ 343 ],
   alphaCSR[ 241 ][ 344 ],
   alphaCSR[ 241 ][ 345 ],
   alphaCSR[ 241 ][ 346 ],
   alphaCSR[ 241 ][ 347 ],
   alphaCSR[ 241 ][ 348 ],
   alphaCSR[ 241 ][ 349 ],
   alphaCSR[ 241 ][ 350 ],
   alphaCSR[ 241 ][ 351 ],
   alphaCSR[ 241 ][ 352 ],
   alphaCSR[ 241 ][ 353 ],
   alphaCSR[ 241 ][ 354 ],
   alphaCSR[ 241 ][ 355 ],
   alphaCSR[ 241 ][ 356 ],
   alphaCSR[ 241 ][ 357 ],
   alphaCSR[ 241 ][ 358 ],
   alphaCSR[ 241 ][ 359 ],
   alphaCSR[ 241 ][ 360 ],
   alphaCSR[ 241 ][ 361 ],
   alphaCSR[ 241 ][ 362 ],
   alphaCSR[ 241 ][ 363 ],
   alphaCSR[ 241 ][ 364 ],
   alphaCSR[ 241 ][ 365 ],
   alphaCSR[ 241 ][ 366 ],
   alphaCSR[ 241 ][ 367 ],
   alphaCSR[ 241 ][ 368 ],
   alphaCSR[ 241 ][ 369 ],
   alphaCSR[ 241 ][ 370 ],
   alphaCSR[ 241 ][ 371 ],
   alphaCSR[ 241 ][ 372 ],
   alphaCSR[ 241 ][ 373 ],
   alphaCSR[ 241 ][ 374 ],
   alphaCSR[ 241 ][ 375 ],
   alphaCSR[ 241 ][ 376 ],
   alphaCSR[ 241 ][ 377 ],
   alphaCSR[ 241 ][ 378 ],
   alphaCSR[ 241 ][ 379 ],
   alphaCSR[ 241 ][ 380 ],
   alphaCSR[ 241 ][ 381 ],
   alphaCSR[ 241 ][ 382 ],
   alphaCSR[ 241 ][ 383 ],
   alphaCSR[ 242 ][ 0 ],
   alphaCSR[ 242 ][ 1 ],
   alphaCSR[ 242 ][ 2 ],
   alphaCSR[ 242 ][ 3 ],
   alphaCSR[ 242 ][ 4 ],
   alphaCSR[ 242 ][ 5 ],
   alphaCSR[ 242 ][ 6 ],
   alphaCSR[ 242 ][ 7 ],
   alphaCSR[ 242 ][ 8 ],
   alphaCSR[ 242 ][ 9 ],
   alphaCSR[ 242 ][ 10 ],
   alphaCSR[ 242 ][ 11 ],
   alphaCSR[ 242 ][ 12 ],
   alphaCSR[ 242 ][ 13 ],
   alphaCSR[ 242 ][ 14 ],
   alphaCSR[ 242 ][ 15 ],
   alphaCSR[ 242 ][ 16 ],
   alphaCSR[ 242 ][ 17 ],
   alphaCSR[ 242 ][ 18 ],
   alphaCSR[ 242 ][ 19 ],
   alphaCSR[ 242 ][ 20 ],
   alphaCSR[ 242 ][ 21 ],
   alphaCSR[ 242 ][ 22 ],
   alphaCSR[ 242 ][ 23 ],
   alphaCSR[ 242 ][ 24 ],
   alphaCSR[ 242 ][ 25 ],
   alphaCSR[ 242 ][ 26 ],
   alphaCSR[ 242 ][ 27 ],
   alphaCSR[ 242 ][ 28 ],
   alphaCSR[ 242 ][ 29 ],
   alphaCSR[ 242 ][ 30 ],
   alphaCSR[ 242 ][ 31 ],
   alphaCSR[ 242 ][ 32 ],
   alphaCSR[ 242 ][ 33 ],
   alphaCSR[ 242 ][ 34 ],
   alphaCSR[ 242 ][ 35 ],
   alphaCSR[ 242 ][ 36 ],
   alphaCSR[ 242 ][ 37 ],
   alphaCSR[ 242 ][ 38 ],
   alphaCSR[ 242 ][ 39 ],
   alphaCSR[ 242 ][ 40 ],
   alphaCSR[ 242 ][ 41 ],
   alphaCSR[ 242 ][ 42 ],
   alphaCSR[ 242 ][ 43 ],
   alphaCSR[ 242 ][ 44 ],
   alphaCSR[ 242 ][ 45 ],
   alphaCSR[ 242 ][ 46 ],
   alphaCSR[ 242 ][ 47 ],
   alphaCSR[ 242 ][ 48 ],
   alphaCSR[ 242 ][ 49 ],
   alphaCSR[ 242 ][ 50 ],
   alphaCSR[ 242 ][ 51 ],
   alphaCSR[ 242 ][ 52 ],
   alphaCSR[ 242 ][ 53 ],
   alphaCSR[ 242 ][ 54 ],
   alphaCSR[ 242 ][ 55 ],
   alphaCSR[ 242 ][ 56 ],
   alphaCSR[ 242 ][ 57 ],
   alphaCSR[ 242 ][ 58 ],
   alphaCSR[ 242 ][ 59 ],
   alphaCSR[ 242 ][ 60 ],
   alphaCSR[ 242 ][ 61 ],
   alphaCSR[ 242 ][ 62 ],
   alphaCSR[ 242 ][ 63 ],
   alphaCSR[ 242 ][ 64 ],
   alphaCSR[ 242 ][ 65 ],
   alphaCSR[ 242 ][ 66 ],
   alphaCSR[ 242 ][ 67 ],
   alphaCSR[ 242 ][ 68 ],
   alphaCSR[ 242 ][ 69 ],
   alphaCSR[ 242 ][ 70 ],
   alphaCSR[ 242 ][ 71 ],
   alphaCSR[ 242 ][ 72 ],
   alphaCSR[ 242 ][ 73 ],
   alphaCSR[ 242 ][ 74 ],
   alphaCSR[ 242 ][ 75 ],
   alphaCSR[ 242 ][ 76 ],
   alphaCSR[ 242 ][ 77 ],
   alphaCSR[ 242 ][ 78 ],
   alphaCSR[ 242 ][ 79 ],
   alphaCSR[ 242 ][ 80 ],
   alphaCSR[ 242 ][ 81 ],
   alphaCSR[ 242 ][ 82 ],
   alphaCSR[ 242 ][ 83 ],
   alphaCSR[ 242 ][ 84 ],
   alphaCSR[ 242 ][ 85 ],
   alphaCSR[ 242 ][ 86 ],
   alphaCSR[ 242 ][ 87 ],
   alphaCSR[ 242 ][ 88 ],
   alphaCSR[ 242 ][ 89 ],
   alphaCSR[ 242 ][ 90 ],
   alphaCSR[ 242 ][ 91 ],
   alphaCSR[ 242 ][ 92 ],
   alphaCSR[ 242 ][ 93 ],
   alphaCSR[ 242 ][ 94 ],
   alphaCSR[ 242 ][ 95 ],
   alphaCSR[ 242 ][ 96 ],
   alphaCSR[ 242 ][ 97 ],
   alphaCSR[ 242 ][ 98 ],
   alphaCSR[ 242 ][ 99 ],
   alphaCSR[ 242 ][ 100 ],
   alphaCSR[ 242 ][ 101 ],
   alphaCSR[ 242 ][ 102 ],
   alphaCSR[ 242 ][ 103 ],
   alphaCSR[ 242 ][ 104 ],
   alphaCSR[ 242 ][ 105 ],
   alphaCSR[ 242 ][ 106 ],
   alphaCSR[ 242 ][ 107 ],
   alphaCSR[ 242 ][ 108 ],
   alphaCSR[ 242 ][ 109 ],
   alphaCSR[ 242 ][ 110 ],
   alphaCSR[ 242 ][ 111 ],
   alphaCSR[ 242 ][ 112 ],
   alphaCSR[ 242 ][ 113 ],
   alphaCSR[ 242 ][ 114 ],
   alphaCSR[ 242 ][ 115 ],
   alphaCSR[ 242 ][ 116 ],
   alphaCSR[ 242 ][ 117 ],
   alphaCSR[ 242 ][ 118 ],
   alphaCSR[ 242 ][ 119 ],
   alphaCSR[ 242 ][ 120 ],
   alphaCSR[ 242 ][ 121 ],
   alphaCSR[ 242 ][ 122 ],
   alphaCSR[ 242 ][ 123 ],
   alphaCSR[ 242 ][ 124 ],
   alphaCSR[ 242 ][ 125 ],
   alphaCSR[ 242 ][ 126 ],
   alphaCSR[ 242 ][ 127 ],
   alphaCSR[ 242 ][ 128 ],
   alphaCSR[ 242 ][ 129 ],
   alphaCSR[ 242 ][ 130 ],
   alphaCSR[ 242 ][ 131 ],
   alphaCSR[ 242 ][ 132 ],
   alphaCSR[ 242 ][ 133 ],
   alphaCSR[ 242 ][ 134 ],
   alphaCSR[ 242 ][ 135 ],
   alphaCSR[ 242 ][ 136 ],
   alphaCSR[ 242 ][ 137 ],
   alphaCSR[ 242 ][ 138 ],
   alphaCSR[ 242 ][ 139 ],
   alphaCSR[ 242 ][ 140 ],
   alphaCSR[ 242 ][ 141 ],
   alphaCSR[ 242 ][ 142 ],
   alphaCSR[ 242 ][ 143 ],
   alphaCSR[ 242 ][ 144 ],
   alphaCSR[ 242 ][ 145 ],
   alphaCSR[ 242 ][ 146 ],
   alphaCSR[ 242 ][ 147 ],
   alphaCSR[ 242 ][ 148 ],
   alphaCSR[ 242 ][ 149 ],
   alphaCSR[ 242 ][ 150 ],
   alphaCSR[ 242 ][ 151 ],
   alphaCSR[ 242 ][ 152 ],
   alphaCSR[ 242 ][ 153 ],
   alphaCSR[ 242 ][ 154 ],
   alphaCSR[ 242 ][ 155 ],
   alphaCSR[ 242 ][ 156 ],
   alphaCSR[ 242 ][ 157 ],
   alphaCSR[ 242 ][ 158 ],
   alphaCSR[ 242 ][ 159 ],
   alphaCSR[ 242 ][ 160 ],
   alphaCSR[ 242 ][ 161 ],
   alphaCSR[ 242 ][ 162 ],
   alphaCSR[ 242 ][ 163 ],
   alphaCSR[ 242 ][ 164 ],
   alphaCSR[ 242 ][ 165 ],
   alphaCSR[ 242 ][ 166 ],
   alphaCSR[ 242 ][ 167 ],
   alphaCSR[ 242 ][ 168 ],
   alphaCSR[ 242 ][ 169 ],
   alphaCSR[ 242 ][ 170 ],
   alphaCSR[ 242 ][ 171 ],
   alphaCSR[ 242 ][ 172 ],
   alphaCSR[ 242 ][ 173 ],
   alphaCSR[ 242 ][ 174 ],
   alphaCSR[ 242 ][ 175 ],
   alphaCSR[ 242 ][ 176 ],
   alphaCSR[ 242 ][ 177 ],
   alphaCSR[ 242 ][ 178 ],
   alphaCSR[ 242 ][ 179 ],
   alphaCSR[ 242 ][ 180 ],
   alphaCSR[ 242 ][ 181 ],
   alphaCSR[ 242 ][ 182 ],
   alphaCSR[ 242 ][ 183 ],
   alphaCSR[ 242 ][ 184 ],
   alphaCSR[ 242 ][ 185 ],
   alphaCSR[ 242 ][ 186 ],
   alphaCSR[ 242 ][ 187 ],
   alphaCSR[ 242 ][ 188 ],
   alphaCSR[ 242 ][ 189 ],
   alphaCSR[ 242 ][ 190 ],
   alphaCSR[ 242 ][ 191 ],
   alphaCSR[ 242 ][ 192 ],
   alphaCSR[ 242 ][ 193 ],
   alphaCSR[ 242 ][ 194 ],
   alphaCSR[ 242 ][ 195 ],
   alphaCSR[ 242 ][ 196 ],
   alphaCSR[ 242 ][ 197 ],
   alphaCSR[ 242 ][ 198 ],
   alphaCSR[ 242 ][ 199 ],
   alphaCSR[ 242 ][ 200 ],
   alphaCSR[ 242 ][ 201 ],
   alphaCSR[ 242 ][ 202 ],
   alphaCSR[ 242 ][ 203 ],
   alphaCSR[ 242 ][ 204 ],
   alphaCSR[ 242 ][ 205 ],
   alphaCSR[ 242 ][ 206 ],
   alphaCSR[ 242 ][ 207 ],
   alphaCSR[ 242 ][ 208 ],
   alphaCSR[ 242 ][ 209 ],
   alphaCSR[ 242 ][ 210 ],
   alphaCSR[ 242 ][ 211 ],
   alphaCSR[ 242 ][ 212 ],
   alphaCSR[ 242 ][ 213 ],
   alphaCSR[ 242 ][ 214 ],
   alphaCSR[ 242 ][ 215 ],
   alphaCSR[ 242 ][ 216 ],
   alphaCSR[ 242 ][ 217 ],
   alphaCSR[ 242 ][ 218 ],
   alphaCSR[ 242 ][ 219 ],
   alphaCSR[ 242 ][ 220 ],
   alphaCSR[ 242 ][ 221 ],
   alphaCSR[ 242 ][ 222 ],
   alphaCSR[ 242 ][ 223 ],
   alphaCSR[ 242 ][ 224 ],
   alphaCSR[ 242 ][ 225 ],
   alphaCSR[ 242 ][ 226 ],
   alphaCSR[ 242 ][ 227 ],
   alphaCSR[ 242 ][ 228 ],
   alphaCSR[ 242 ][ 229 ],
   alphaCSR[ 242 ][ 230 ],
   alphaCSR[ 242 ][ 231 ],
   alphaCSR[ 242 ][ 232 ],
   alphaCSR[ 242 ][ 233 ],
   alphaCSR[ 242 ][ 234 ],
   alphaCSR[ 242 ][ 235 ],
   alphaCSR[ 242 ][ 236 ],
   alphaCSR[ 242 ][ 237 ],
   alphaCSR[ 242 ][ 238 ],
   alphaCSR[ 242 ][ 239 ],
   alphaCSR[ 242 ][ 240 ],
   alphaCSR[ 242 ][ 241 ],
   alphaCSR[ 242 ][ 242 ],
   alphaCSR[ 242 ][ 243 ],
   alphaCSR[ 242 ][ 244 ],
   alphaCSR[ 242 ][ 245 ],
   alphaCSR[ 242 ][ 246 ],
   alphaCSR[ 242 ][ 247 ],
   alphaCSR[ 242 ][ 248 ],
   alphaCSR[ 242 ][ 249 ],
   alphaCSR[ 242 ][ 250 ],
   alphaCSR[ 242 ][ 251 ],
   alphaCSR[ 242 ][ 252 ],
   alphaCSR[ 242 ][ 253 ],
   alphaCSR[ 242 ][ 254 ],
   alphaCSR[ 242 ][ 255 ],
   alphaCSR[ 242 ][ 256 ],
   alphaCSR[ 242 ][ 257 ],
   alphaCSR[ 242 ][ 258 ],
   alphaCSR[ 242 ][ 259 ],
   alphaCSR[ 242 ][ 260 ],
   alphaCSR[ 242 ][ 261 ],
   alphaCSR[ 242 ][ 262 ],
   alphaCSR[ 242 ][ 263 ],
   alphaCSR[ 242 ][ 264 ],
   alphaCSR[ 242 ][ 265 ],
   alphaCSR[ 242 ][ 266 ],
   alphaCSR[ 242 ][ 267 ],
   alphaCSR[ 242 ][ 268 ],
   alphaCSR[ 242 ][ 269 ],
   alphaCSR[ 242 ][ 270 ],
   alphaCSR[ 242 ][ 271 ],
   alphaCSR[ 242 ][ 272 ],
   alphaCSR[ 242 ][ 273 ],
   alphaCSR[ 242 ][ 274 ],
   alphaCSR[ 242 ][ 275 ],
   alphaCSR[ 242 ][ 276 ],
   alphaCSR[ 242 ][ 277 ],
   alphaCSR[ 242 ][ 278 ],
   alphaCSR[ 242 ][ 279 ],
   alphaCSR[ 242 ][ 280 ],
   alphaCSR[ 242 ][ 281 ],
   alphaCSR[ 242 ][ 282 ],
   alphaCSR[ 242 ][ 283 ],
   alphaCSR[ 242 ][ 284 ],
   alphaCSR[ 242 ][ 285 ],
   alphaCSR[ 242 ][ 286 ],
   alphaCSR[ 242 ][ 287 ],
   alphaCSR[ 242 ][ 288 ],
   alphaCSR[ 242 ][ 289 ],
   alphaCSR[ 242 ][ 290 ],
   alphaCSR[ 242 ][ 291 ],
   alphaCSR[ 242 ][ 292 ],
   alphaCSR[ 242 ][ 293 ],
   alphaCSR[ 242 ][ 294 ],
   alphaCSR[ 242 ][ 295 ],
   alphaCSR[ 242 ][ 296 ],
   alphaCSR[ 242 ][ 297 ],
   alphaCSR[ 242 ][ 298 ],
   alphaCSR[ 242 ][ 299 ],
   alphaCSR[ 242 ][ 300 ],
   alphaCSR[ 242 ][ 301 ],
   alphaCSR[ 242 ][ 302 ],
   alphaCSR[ 242 ][ 303 ],
   alphaCSR[ 242 ][ 304 ],
   alphaCSR[ 242 ][ 305 ],
   alphaCSR[ 242 ][ 306 ],
   alphaCSR[ 242 ][ 307 ],
   alphaCSR[ 242 ][ 308 ],
   alphaCSR[ 242 ][ 309 ],
   alphaCSR[ 242 ][ 310 ],
   alphaCSR[ 242 ][ 311 ],
   alphaCSR[ 242 ][ 312 ],
   alphaCSR[ 242 ][ 313 ],
   alphaCSR[ 242 ][ 314 ],
   alphaCSR[ 242 ][ 315 ],
   alphaCSR[ 242 ][ 316 ],
   alphaCSR[ 242 ][ 317 ],
   alphaCSR[ 242 ][ 318 ],
   alphaCSR[ 242 ][ 319 ],
   alphaCSR[ 242 ][ 320 ],
   alphaCSR[ 242 ][ 321 ],
   alphaCSR[ 242 ][ 322 ],
   alphaCSR[ 242 ][ 323 ],
   alphaCSR[ 242 ][ 324 ],
   alphaCSR[ 242 ][ 325 ],
   alphaCSR[ 242 ][ 326 ],
   alphaCSR[ 242 ][ 327 ],
   alphaCSR[ 242 ][ 328 ],
   alphaCSR[ 242 ][ 329 ],
   alphaCSR[ 242 ][ 330 ],
   alphaCSR[ 242 ][ 331 ],
   alphaCSR[ 242 ][ 332 ],
   alphaCSR[ 242 ][ 333 ],
   alphaCSR[ 242 ][ 334 ],
   alphaCSR[ 242 ][ 335 ],
   alphaCSR[ 242 ][ 336 ],
   alphaCSR[ 242 ][ 337 ],
   alphaCSR[ 242 ][ 338 ],
   alphaCSR[ 242 ][ 339 ],
   alphaCSR[ 242 ][ 340 ],
   alphaCSR[ 242 ][ 341 ],
   alphaCSR[ 242 ][ 342 ],
   alphaCSR[ 242 ][ 343 ],
   alphaCSR[ 242 ][ 344 ],
   alphaCSR[ 242 ][ 345 ],
   alphaCSR[ 242 ][ 346 ],
   alphaCSR[ 242 ][ 347 ],
   alphaCSR[ 242 ][ 348 ],
   alphaCSR[ 242 ][ 349 ],
   alphaCSR[ 242 ][ 350 ],
   alphaCSR[ 242 ][ 351 ],
   alphaCSR[ 242 ][ 352 ],
   alphaCSR[ 242 ][ 353 ],
   alphaCSR[ 242 ][ 354 ],
   alphaCSR[ 242 ][ 355 ],
   alphaCSR[ 242 ][ 356 ],
   alphaCSR[ 242 ][ 357 ],
   alphaCSR[ 242 ][ 358 ],
   alphaCSR[ 242 ][ 359 ],
   alphaCSR[ 242 ][ 360 ],
   alphaCSR[ 242 ][ 361 ],
   alphaCSR[ 242 ][ 362 ],
   alphaCSR[ 242 ][ 363 ],
   alphaCSR[ 242 ][ 364 ],
   alphaCSR[ 242 ][ 365 ],
   alphaCSR[ 242 ][ 366 ],
   alphaCSR[ 242 ][ 367 ],
   alphaCSR[ 242 ][ 368 ],
   alphaCSR[ 242 ][ 369 ],
   alphaCSR[ 242 ][ 370 ],
   alphaCSR[ 242 ][ 371 ],
   alphaCSR[ 242 ][ 372 ],
   alphaCSR[ 242 ][ 373 ],
   alphaCSR[ 242 ][ 374 ],
   alphaCSR[ 242 ][ 375 ],
   alphaCSR[ 242 ][ 376 ],
   alphaCSR[ 242 ][ 377 ],
   alphaCSR[ 242 ][ 378 ],
   alphaCSR[ 242 ][ 379 ],
   alphaCSR[ 242 ][ 380 ],
   alphaCSR[ 242 ][ 381 ],
   alphaCSR[ 242 ][ 382 ],
   alphaCSR[ 242 ][ 383 ],
   alphaCSR[ 243 ][ 0 ],
   alphaCSR[ 243 ][ 1 ],
   alphaCSR[ 243 ][ 2 ],
   alphaCSR[ 243 ][ 3 ],
   alphaCSR[ 243 ][ 4 ],
   alphaCSR[ 243 ][ 5 ],
   alphaCSR[ 243 ][ 6 ],
   alphaCSR[ 243 ][ 7 ],
   alphaCSR[ 243 ][ 8 ],
   alphaCSR[ 243 ][ 9 ],
   alphaCSR[ 243 ][ 10 ],
   alphaCSR[ 243 ][ 11 ],
   alphaCSR[ 243 ][ 12 ],
   alphaCSR[ 243 ][ 13 ],
   alphaCSR[ 243 ][ 14 ],
   alphaCSR[ 243 ][ 15 ],
   alphaCSR[ 243 ][ 16 ],
   alphaCSR[ 243 ][ 17 ],
   alphaCSR[ 243 ][ 18 ],
   alphaCSR[ 243 ][ 19 ],
   alphaCSR[ 243 ][ 20 ],
   alphaCSR[ 243 ][ 21 ],
   alphaCSR[ 243 ][ 22 ],
   alphaCSR[ 243 ][ 23 ],
   alphaCSR[ 243 ][ 24 ],
   alphaCSR[ 243 ][ 25 ],
   alphaCSR[ 243 ][ 26 ],
   alphaCSR[ 243 ][ 27 ],
   alphaCSR[ 243 ][ 28 ],
   alphaCSR[ 243 ][ 29 ],
   alphaCSR[ 243 ][ 30 ],
   alphaCSR[ 243 ][ 31 ],
   alphaCSR[ 243 ][ 32 ],
   alphaCSR[ 243 ][ 33 ],
   alphaCSR[ 243 ][ 34 ],
   alphaCSR[ 243 ][ 35 ],
   alphaCSR[ 243 ][ 36 ],
   alphaCSR[ 243 ][ 37 ],
   alphaCSR[ 243 ][ 38 ],
   alphaCSR[ 243 ][ 39 ],
   alphaCSR[ 243 ][ 40 ],
   alphaCSR[ 243 ][ 41 ],
   alphaCSR[ 243 ][ 42 ],
   alphaCSR[ 243 ][ 43 ],
   alphaCSR[ 243 ][ 44 ],
   alphaCSR[ 243 ][ 45 ],
   alphaCSR[ 243 ][ 46 ],
   alphaCSR[ 243 ][ 47 ],
   alphaCSR[ 243 ][ 48 ],
   alphaCSR[ 243 ][ 49 ],
   alphaCSR[ 243 ][ 50 ],
   alphaCSR[ 243 ][ 51 ],
   alphaCSR[ 243 ][ 52 ],
   alphaCSR[ 243 ][ 53 ],
   alphaCSR[ 243 ][ 54 ],
   alphaCSR[ 243 ][ 55 ],
   alphaCSR[ 243 ][ 56 ],
   alphaCSR[ 243 ][ 57 ],
   alphaCSR[ 243 ][ 58 ],
   alphaCSR[ 243 ][ 59 ],
   alphaCSR[ 243 ][ 60 ],
   alphaCSR[ 243 ][ 61 ],
   alphaCSR[ 243 ][ 62 ],
   alphaCSR[ 243 ][ 63 ],
   alphaCSR[ 243 ][ 64 ],
   alphaCSR[ 243 ][ 65 ],
   alphaCSR[ 243 ][ 66 ],
   alphaCSR[ 243 ][ 67 ],
   alphaCSR[ 243 ][ 68 ],
   alphaCSR[ 243 ][ 69 ],
   alphaCSR[ 243 ][ 70 ],
   alphaCSR[ 243 ][ 71 ],
   alphaCSR[ 243 ][ 72 ],
   alphaCSR[ 243 ][ 73 ],
   alphaCSR[ 243 ][ 74 ],
   alphaCSR[ 243 ][ 75 ],
   alphaCSR[ 243 ][ 76 ],
   alphaCSR[ 243 ][ 77 ],
   alphaCSR[ 243 ][ 78 ],
   alphaCSR[ 243 ][ 79 ],
   alphaCSR[ 243 ][ 80 ],
   alphaCSR[ 243 ][ 81 ],
   alphaCSR[ 243 ][ 82 ],
   alphaCSR[ 243 ][ 83 ],
   alphaCSR[ 243 ][ 84 ],
   alphaCSR[ 243 ][ 85 ],
   alphaCSR[ 243 ][ 86 ],
   alphaCSR[ 243 ][ 87 ],
   alphaCSR[ 243 ][ 88 ],
   alphaCSR[ 243 ][ 89 ],
   alphaCSR[ 243 ][ 90 ],
   alphaCSR[ 243 ][ 91 ],
   alphaCSR[ 243 ][ 92 ],
   alphaCSR[ 243 ][ 93 ],
   alphaCSR[ 243 ][ 94 ],
   alphaCSR[ 243 ][ 95 ],
   alphaCSR[ 243 ][ 96 ],
   alphaCSR[ 243 ][ 97 ],
   alphaCSR[ 243 ][ 98 ],
   alphaCSR[ 243 ][ 99 ],
   alphaCSR[ 243 ][ 100 ],
   alphaCSR[ 243 ][ 101 ],
   alphaCSR[ 243 ][ 102 ],
   alphaCSR[ 243 ][ 103 ],
   alphaCSR[ 243 ][ 104 ],
   alphaCSR[ 243 ][ 105 ],
   alphaCSR[ 243 ][ 106 ],
   alphaCSR[ 243 ][ 107 ],
   alphaCSR[ 243 ][ 108 ],
   alphaCSR[ 243 ][ 109 ],
   alphaCSR[ 243 ][ 110 ],
   alphaCSR[ 243 ][ 111 ],
   alphaCSR[ 243 ][ 112 ],
   alphaCSR[ 243 ][ 113 ],
   alphaCSR[ 243 ][ 114 ],
   alphaCSR[ 243 ][ 115 ],
   alphaCSR[ 243 ][ 116 ],
   alphaCSR[ 243 ][ 117 ],
   alphaCSR[ 243 ][ 118 ],
   alphaCSR[ 243 ][ 119 ],
   alphaCSR[ 243 ][ 120 ],
   alphaCSR[ 243 ][ 121 ],
   alphaCSR[ 243 ][ 122 ],
   alphaCSR[ 243 ][ 123 ],
   alphaCSR[ 243 ][ 124 ],
   alphaCSR[ 243 ][ 125 ],
   alphaCSR[ 243 ][ 126 ],
   alphaCSR[ 243 ][ 127 ],
   alphaCSR[ 243 ][ 128 ],
   alphaCSR[ 243 ][ 129 ],
   alphaCSR[ 243 ][ 130 ],
   alphaCSR[ 243 ][ 131 ],
   alphaCSR[ 243 ][ 132 ],
   alphaCSR[ 243 ][ 133 ],
   alphaCSR[ 243 ][ 134 ],
   alphaCSR[ 243 ][ 135 ],
   alphaCSR[ 243 ][ 136 ],
   alphaCSR[ 243 ][ 137 ],
   alphaCSR[ 243 ][ 138 ],
   alphaCSR[ 243 ][ 139 ],
   alphaCSR[ 243 ][ 140 ],
   alphaCSR[ 243 ][ 141 ],
   alphaCSR[ 243 ][ 142 ],
   alphaCSR[ 243 ][ 143 ],
   alphaCSR[ 243 ][ 144 ],
   alphaCSR[ 243 ][ 145 ],
   alphaCSR[ 243 ][ 146 ],
   alphaCSR[ 243 ][ 147 ],
   alphaCSR[ 243 ][ 148 ],
   alphaCSR[ 243 ][ 149 ],
   alphaCSR[ 243 ][ 150 ],
   alphaCSR[ 243 ][ 151 ],
   alphaCSR[ 243 ][ 152 ],
   alphaCSR[ 243 ][ 153 ],
   alphaCSR[ 243 ][ 154 ],
   alphaCSR[ 243 ][ 155 ],
   alphaCSR[ 243 ][ 156 ],
   alphaCSR[ 243 ][ 157 ],
   alphaCSR[ 243 ][ 158 ],
   alphaCSR[ 243 ][ 159 ],
   alphaCSR[ 243 ][ 160 ],
   alphaCSR[ 243 ][ 161 ],
   alphaCSR[ 243 ][ 162 ],
   alphaCSR[ 243 ][ 163 ],
   alphaCSR[ 243 ][ 164 ],
   alphaCSR[ 243 ][ 165 ],
   alphaCSR[ 243 ][ 166 ],
   alphaCSR[ 243 ][ 167 ],
   alphaCSR[ 243 ][ 168 ],
   alphaCSR[ 243 ][ 169 ],
   alphaCSR[ 243 ][ 170 ],
   alphaCSR[ 243 ][ 171 ],
   alphaCSR[ 243 ][ 172 ],
   alphaCSR[ 243 ][ 173 ],
   alphaCSR[ 243 ][ 174 ],
   alphaCSR[ 243 ][ 175 ],
   alphaCSR[ 243 ][ 176 ],
   alphaCSR[ 243 ][ 177 ],
   alphaCSR[ 243 ][ 178 ],
   alphaCSR[ 243 ][ 179 ],
   alphaCSR[ 243 ][ 180 ],
   alphaCSR[ 243 ][ 181 ],
   alphaCSR[ 243 ][ 182 ],
   alphaCSR[ 243 ][ 183 ],
   alphaCSR[ 243 ][ 184 ],
   alphaCSR[ 243 ][ 185 ],
   alphaCSR[ 243 ][ 186 ],
   alphaCSR[ 243 ][ 187 ],
   alphaCSR[ 243 ][ 188 ],
   alphaCSR[ 243 ][ 189 ],
   alphaCSR[ 243 ][ 190 ],
   alphaCSR[ 243 ][ 191 ],
   alphaCSR[ 243 ][ 192 ],
   alphaCSR[ 243 ][ 193 ],
   alphaCSR[ 243 ][ 194 ],
   alphaCSR[ 243 ][ 195 ],
   alphaCSR[ 243 ][ 196 ],
   alphaCSR[ 243 ][ 197 ],
   alphaCSR[ 243 ][ 198 ],
   alphaCSR[ 243 ][ 199 ],
   alphaCSR[ 243 ][ 200 ],
   alphaCSR[ 243 ][ 201 ],
   alphaCSR[ 243 ][ 202 ],
   alphaCSR[ 243 ][ 203 ],
   alphaCSR[ 243 ][ 204 ],
   alphaCSR[ 243 ][ 205 ],
   alphaCSR[ 243 ][ 206 ],
   alphaCSR[ 243 ][ 207 ],
   alphaCSR[ 243 ][ 208 ],
   alphaCSR[ 243 ][ 209 ],
   alphaCSR[ 243 ][ 210 ],
   alphaCSR[ 243 ][ 211 ],
   alphaCSR[ 243 ][ 212 ],
   alphaCSR[ 243 ][ 213 ],
   alphaCSR[ 243 ][ 214 ],
   alphaCSR[ 243 ][ 215 ],
   alphaCSR[ 243 ][ 216 ],
   alphaCSR[ 243 ][ 217 ],
   alphaCSR[ 243 ][ 218 ],
   alphaCSR[ 243 ][ 219 ],
   alphaCSR[ 243 ][ 220 ],
   alphaCSR[ 243 ][ 221 ],
   alphaCSR[ 243 ][ 222 ],
   alphaCSR[ 243 ][ 223 ],
   alphaCSR[ 243 ][ 224 ],
   alphaCSR[ 243 ][ 225 ],
   alphaCSR[ 243 ][ 226 ],
   alphaCSR[ 243 ][ 227 ],
   alphaCSR[ 243 ][ 228 ],
   alphaCSR[ 243 ][ 229 ],
   alphaCSR[ 243 ][ 230 ],
   alphaCSR[ 243 ][ 231 ],
   alphaCSR[ 243 ][ 232 ],
   alphaCSR[ 243 ][ 233 ],
   alphaCSR[ 243 ][ 234 ],
   alphaCSR[ 243 ][ 235 ],
   alphaCSR[ 243 ][ 236 ],
   alphaCSR[ 243 ][ 237 ],
   alphaCSR[ 243 ][ 238 ],
   alphaCSR[ 243 ][ 239 ],
   alphaCSR[ 243 ][ 240 ],
   alphaCSR[ 243 ][ 241 ],
   alphaCSR[ 243 ][ 242 ],
   alphaCSR[ 243 ][ 243 ],
   alphaCSR[ 243 ][ 244 ],
   alphaCSR[ 243 ][ 245 ],
   alphaCSR[ 243 ][ 246 ],
   alphaCSR[ 243 ][ 247 ],
   alphaCSR[ 243 ][ 248 ],
   alphaCSR[ 243 ][ 249 ],
   alphaCSR[ 243 ][ 250 ],
   alphaCSR[ 243 ][ 251 ],
   alphaCSR[ 243 ][ 252 ],
   alphaCSR[ 243 ][ 253 ],
   alphaCSR[ 243 ][ 254 ],
   alphaCSR[ 243 ][ 255 ],
   alphaCSR[ 243 ][ 256 ],
   alphaCSR[ 243 ][ 257 ],
   alphaCSR[ 243 ][ 258 ],
   alphaCSR[ 243 ][ 259 ],
   alphaCSR[ 243 ][ 260 ],
   alphaCSR[ 243 ][ 261 ],
   alphaCSR[ 243 ][ 262 ],
   alphaCSR[ 243 ][ 263 ],
   alphaCSR[ 243 ][ 264 ],
   alphaCSR[ 243 ][ 265 ],
   alphaCSR[ 243 ][ 266 ],
   alphaCSR[ 243 ][ 267 ],
   alphaCSR[ 243 ][ 268 ],
   alphaCSR[ 243 ][ 269 ],
   alphaCSR[ 243 ][ 270 ],
   alphaCSR[ 243 ][ 271 ],
   alphaCSR[ 243 ][ 272 ],
   alphaCSR[ 243 ][ 273 ],
   alphaCSR[ 243 ][ 274 ],
   alphaCSR[ 243 ][ 275 ],
   alphaCSR[ 243 ][ 276 ],
   alphaCSR[ 243 ][ 277 ],
   alphaCSR[ 243 ][ 278 ],
   alphaCSR[ 243 ][ 279 ],
   alphaCSR[ 243 ][ 280 ],
   alphaCSR[ 243 ][ 281 ],
   alphaCSR[ 243 ][ 282 ],
   alphaCSR[ 243 ][ 283 ],
   alphaCSR[ 243 ][ 284 ],
   alphaCSR[ 243 ][ 285 ],
   alphaCSR[ 243 ][ 286 ],
   alphaCSR[ 243 ][ 287 ],
   alphaCSR[ 243 ][ 288 ],
   alphaCSR[ 243 ][ 289 ],
   alphaCSR[ 243 ][ 290 ],
   alphaCSR[ 243 ][ 291 ],
   alphaCSR[ 243 ][ 292 ],
   alphaCSR[ 243 ][ 293 ],
   alphaCSR[ 243 ][ 294 ],
   alphaCSR[ 243 ][ 295 ],
   alphaCSR[ 243 ][ 296 ],
   alphaCSR[ 243 ][ 297 ],
   alphaCSR[ 243 ][ 298 ],
   alphaCSR[ 243 ][ 299 ],
   alphaCSR[ 243 ][ 300 ],
   alphaCSR[ 243 ][ 301 ],
   alphaCSR[ 243 ][ 302 ],
   alphaCSR[ 243 ][ 303 ],
   alphaCSR[ 243 ][ 304 ],
   alphaCSR[ 243 ][ 305 ],
   alphaCSR[ 243 ][ 306 ],
   alphaCSR[ 243 ][ 307 ],
   alphaCSR[ 243 ][ 308 ],
   alphaCSR[ 243 ][ 309 ],
   alphaCSR[ 243 ][ 310 ],
   alphaCSR[ 243 ][ 311 ],
   alphaCSR[ 243 ][ 312 ],
   alphaCSR[ 243 ][ 313 ],
   alphaCSR[ 243 ][ 314 ],
   alphaCSR[ 243 ][ 315 ],
   alphaCSR[ 243 ][ 316 ],
   alphaCSR[ 243 ][ 317 ],
   alphaCSR[ 243 ][ 318 ],
   alphaCSR[ 243 ][ 319 ],
   alphaCSR[ 243 ][ 320 ],
   alphaCSR[ 243 ][ 321 ],
   alphaCSR[ 243 ][ 322 ],
   alphaCSR[ 243 ][ 323 ],
   alphaCSR[ 243 ][ 324 ],
   alphaCSR[ 243 ][ 325 ],
   alphaCSR[ 243 ][ 326 ],
   alphaCSR[ 243 ][ 327 ],
   alphaCSR[ 243 ][ 328 ],
   alphaCSR[ 243 ][ 329 ],
   alphaCSR[ 243 ][ 330 ],
   alphaCSR[ 243 ][ 331 ],
   alphaCSR[ 243 ][ 332 ],
   alphaCSR[ 243 ][ 333 ],
   alphaCSR[ 243 ][ 334 ],
   alphaCSR[ 243 ][ 335 ],
   alphaCSR[ 243 ][ 336 ],
   alphaCSR[ 243 ][ 337 ],
   alphaCSR[ 243 ][ 338 ],
   alphaCSR[ 243 ][ 339 ],
   alphaCSR[ 243 ][ 340 ],
   alphaCSR[ 243 ][ 341 ],
   alphaCSR[ 243 ][ 342 ],
   alphaCSR[ 243 ][ 343 ],
   alphaCSR[ 243 ][ 344 ],
   alphaCSR[ 243 ][ 345 ],
   alphaCSR[ 243 ][ 346 ],
   alphaCSR[ 243 ][ 347 ],
   alphaCSR[ 243 ][ 348 ],
   alphaCSR[ 243 ][ 349 ],
   alphaCSR[ 243 ][ 350 ],
   alphaCSR[ 243 ][ 351 ],
   alphaCSR[ 243 ][ 352 ],
   alphaCSR[ 243 ][ 353 ],
   alphaCSR[ 243 ][ 354 ],
   alphaCSR[ 243 ][ 355 ],
   alphaCSR[ 243 ][ 356 ],
   alphaCSR[ 243 ][ 357 ],
   alphaCSR[ 243 ][ 358 ],
   alphaCSR[ 243 ][ 359 ],
   alphaCSR[ 243 ][ 360 ],
   alphaCSR[ 243 ][ 361 ],
   alphaCSR[ 243 ][ 362 ],
   alphaCSR[ 243 ][ 363 ],
   alphaCSR[ 243 ][ 364 ],
   alphaCSR[ 243 ][ 365 ],
   alphaCSR[ 243 ][ 366 ],
   alphaCSR[ 243 ][ 367 ],
   alphaCSR[ 243 ][ 368 ],
   alphaCSR[ 243 ][ 369 ],
   alphaCSR[ 243 ][ 370 ],
   alphaCSR[ 243 ][ 371 ],
   alphaCSR[ 243 ][ 372 ],
   alphaCSR[ 243 ][ 373 ],
   alphaCSR[ 243 ][ 374 ],
   alphaCSR[ 243 ][ 375 ],
   alphaCSR[ 243 ][ 376 ],
   alphaCSR[ 243 ][ 377 ],
   alphaCSR[ 243 ][ 378 ],
   alphaCSR[ 243 ][ 379 ],
   alphaCSR[ 243 ][ 380 ],
   alphaCSR[ 243 ][ 381 ],
   alphaCSR[ 243 ][ 382 ],
   alphaCSR[ 243 ][ 383 ],
   alphaCSR[ 244 ][ 0 ],
   alphaCSR[ 244 ][ 1 ],
   alphaCSR[ 244 ][ 2 ],
   alphaCSR[ 244 ][ 3 ],
   alphaCSR[ 244 ][ 4 ],
   alphaCSR[ 244 ][ 5 ],
   alphaCSR[ 244 ][ 6 ],
   alphaCSR[ 244 ][ 7 ],
   alphaCSR[ 244 ][ 8 ],
   alphaCSR[ 244 ][ 9 ],
   alphaCSR[ 244 ][ 10 ],
   alphaCSR[ 244 ][ 11 ],
   alphaCSR[ 244 ][ 12 ],
   alphaCSR[ 244 ][ 13 ],
   alphaCSR[ 244 ][ 14 ],
   alphaCSR[ 244 ][ 15 ],
   alphaCSR[ 244 ][ 16 ],
   alphaCSR[ 244 ][ 17 ],
   alphaCSR[ 244 ][ 18 ],
   alphaCSR[ 244 ][ 19 ],
   alphaCSR[ 244 ][ 20 ],
   alphaCSR[ 244 ][ 21 ],
   alphaCSR[ 244 ][ 22 ],
   alphaCSR[ 244 ][ 23 ],
   alphaCSR[ 244 ][ 24 ],
   alphaCSR[ 244 ][ 25 ],
   alphaCSR[ 244 ][ 26 ],
   alphaCSR[ 244 ][ 27 ],
   alphaCSR[ 244 ][ 28 ],
   alphaCSR[ 244 ][ 29 ],
   alphaCSR[ 244 ][ 30 ],
   alphaCSR[ 244 ][ 31 ],
   alphaCSR[ 244 ][ 32 ],
   alphaCSR[ 244 ][ 33 ],
   alphaCSR[ 244 ][ 34 ],
   alphaCSR[ 244 ][ 35 ],
   alphaCSR[ 244 ][ 36 ],
   alphaCSR[ 244 ][ 37 ],
   alphaCSR[ 244 ][ 38 ],
   alphaCSR[ 244 ][ 39 ],
   alphaCSR[ 244 ][ 40 ],
   alphaCSR[ 244 ][ 41 ],
   alphaCSR[ 244 ][ 42 ],
   alphaCSR[ 244 ][ 43 ],
   alphaCSR[ 244 ][ 44 ],
   alphaCSR[ 244 ][ 45 ],
   alphaCSR[ 244 ][ 46 ],
   alphaCSR[ 244 ][ 47 ],
   alphaCSR[ 244 ][ 48 ],
   alphaCSR[ 244 ][ 49 ],
   alphaCSR[ 244 ][ 50 ],
   alphaCSR[ 244 ][ 51 ],
   alphaCSR[ 244 ][ 52 ],
   alphaCSR[ 244 ][ 53 ],
   alphaCSR[ 244 ][ 54 ],
   alphaCSR[ 244 ][ 55 ],
   alphaCSR[ 244 ][ 56 ],
   alphaCSR[ 244 ][ 57 ],
   alphaCSR[ 244 ][ 58 ],
   alphaCSR[ 244 ][ 59 ],
   alphaCSR[ 244 ][ 60 ],
   alphaCSR[ 244 ][ 61 ],
   alphaCSR[ 244 ][ 62 ],
   alphaCSR[ 244 ][ 63 ],
   alphaCSR[ 244 ][ 64 ],
   alphaCSR[ 244 ][ 65 ],
   alphaCSR[ 244 ][ 66 ],
   alphaCSR[ 244 ][ 67 ],
   alphaCSR[ 244 ][ 68 ],
   alphaCSR[ 244 ][ 69 ],
   alphaCSR[ 244 ][ 70 ],
   alphaCSR[ 244 ][ 71 ],
   alphaCSR[ 244 ][ 72 ],
   alphaCSR[ 244 ][ 73 ],
   alphaCSR[ 244 ][ 74 ],
   alphaCSR[ 244 ][ 75 ],
   alphaCSR[ 244 ][ 76 ],
   alphaCSR[ 244 ][ 77 ],
   alphaCSR[ 244 ][ 78 ],
   alphaCSR[ 244 ][ 79 ],
   alphaCSR[ 244 ][ 80 ],
   alphaCSR[ 244 ][ 81 ],
   alphaCSR[ 244 ][ 82 ],
   alphaCSR[ 244 ][ 83 ],
   alphaCSR[ 244 ][ 84 ],
   alphaCSR[ 244 ][ 85 ],
   alphaCSR[ 244 ][ 86 ],
   alphaCSR[ 244 ][ 87 ],
   alphaCSR[ 244 ][ 88 ],
   alphaCSR[ 244 ][ 89 ],
   alphaCSR[ 244 ][ 90 ],
   alphaCSR[ 244 ][ 91 ],
   alphaCSR[ 244 ][ 92 ],
   alphaCSR[ 244 ][ 93 ],
   alphaCSR[ 244 ][ 94 ],
   alphaCSR[ 244 ][ 95 ],
   alphaCSR[ 244 ][ 96 ],
   alphaCSR[ 244 ][ 97 ],
   alphaCSR[ 244 ][ 98 ],
   alphaCSR[ 244 ][ 99 ],
   alphaCSR[ 244 ][ 100 ],
   alphaCSR[ 244 ][ 101 ],
   alphaCSR[ 244 ][ 102 ],
   alphaCSR[ 244 ][ 103 ],
   alphaCSR[ 244 ][ 104 ],
   alphaCSR[ 244 ][ 105 ],
   alphaCSR[ 244 ][ 106 ],
   alphaCSR[ 244 ][ 107 ],
   alphaCSR[ 244 ][ 108 ],
   alphaCSR[ 244 ][ 109 ],
   alphaCSR[ 244 ][ 110 ],
   alphaCSR[ 244 ][ 111 ],
   alphaCSR[ 244 ][ 112 ],
   alphaCSR[ 244 ][ 113 ],
   alphaCSR[ 244 ][ 114 ],
   alphaCSR[ 244 ][ 115 ],
   alphaCSR[ 244 ][ 116 ],
   alphaCSR[ 244 ][ 117 ],
   alphaCSR[ 244 ][ 118 ],
   alphaCSR[ 244 ][ 119 ],
   alphaCSR[ 244 ][ 120 ],
   alphaCSR[ 244 ][ 121 ],
   alphaCSR[ 244 ][ 122 ],
   alphaCSR[ 244 ][ 123 ],
   alphaCSR[ 244 ][ 124 ],
   alphaCSR[ 244 ][ 125 ],
   alphaCSR[ 244 ][ 126 ],
   alphaCSR[ 244 ][ 127 ],
   alphaCSR[ 244 ][ 128 ],
   alphaCSR[ 244 ][ 129 ],
   alphaCSR[ 244 ][ 130 ],
   alphaCSR[ 244 ][ 131 ],
   alphaCSR[ 244 ][ 132 ],
   alphaCSR[ 244 ][ 133 ],
   alphaCSR[ 244 ][ 134 ],
   alphaCSR[ 244 ][ 135 ],
   alphaCSR[ 244 ][ 136 ],
   alphaCSR[ 244 ][ 137 ],
   alphaCSR[ 244 ][ 138 ],
   alphaCSR[ 244 ][ 139 ],
   alphaCSR[ 244 ][ 140 ],
   alphaCSR[ 244 ][ 141 ],
   alphaCSR[ 244 ][ 142 ],
   alphaCSR[ 244 ][ 143 ],
   alphaCSR[ 244 ][ 144 ],
   alphaCSR[ 244 ][ 145 ],
   alphaCSR[ 244 ][ 146 ],
   alphaCSR[ 244 ][ 147 ],
   alphaCSR[ 244 ][ 148 ],
   alphaCSR[ 244 ][ 149 ],
   alphaCSR[ 244 ][ 150 ],
   alphaCSR[ 244 ][ 151 ],
   alphaCSR[ 244 ][ 152 ],
   alphaCSR[ 244 ][ 153 ],
   alphaCSR[ 244 ][ 154 ],
   alphaCSR[ 244 ][ 155 ],
   alphaCSR[ 244 ][ 156 ],
   alphaCSR[ 244 ][ 157 ],
   alphaCSR[ 244 ][ 158 ],
   alphaCSR[ 244 ][ 159 ],
   alphaCSR[ 244 ][ 160 ],
   alphaCSR[ 244 ][ 161 ],
   alphaCSR[ 244 ][ 162 ],
   alphaCSR[ 244 ][ 163 ],
   alphaCSR[ 244 ][ 164 ],
   alphaCSR[ 244 ][ 165 ],
   alphaCSR[ 244 ][ 166 ],
   alphaCSR[ 244 ][ 167 ],
   alphaCSR[ 244 ][ 168 ],
   alphaCSR[ 244 ][ 169 ],
   alphaCSR[ 244 ][ 170 ],
   alphaCSR[ 244 ][ 171 ],
   alphaCSR[ 244 ][ 172 ],
   alphaCSR[ 244 ][ 173 ],
   alphaCSR[ 244 ][ 174 ],
   alphaCSR[ 244 ][ 175 ],
   alphaCSR[ 244 ][ 176 ],
   alphaCSR[ 244 ][ 177 ],
   alphaCSR[ 244 ][ 178 ],
   alphaCSR[ 244 ][ 179 ],
   alphaCSR[ 244 ][ 180 ],
   alphaCSR[ 244 ][ 181 ],
   alphaCSR[ 244 ][ 182 ],
   alphaCSR[ 244 ][ 183 ],
   alphaCSR[ 244 ][ 184 ],
   alphaCSR[ 244 ][ 185 ],
   alphaCSR[ 244 ][ 186 ],
   alphaCSR[ 244 ][ 187 ],
   alphaCSR[ 244 ][ 188 ],
   alphaCSR[ 244 ][ 189 ],
   alphaCSR[ 244 ][ 190 ],
   alphaCSR[ 244 ][ 191 ],
   alphaCSR[ 244 ][ 192 ],
   alphaCSR[ 244 ][ 193 ],
   alphaCSR[ 244 ][ 194 ],
   alphaCSR[ 244 ][ 195 ],
   alphaCSR[ 244 ][ 196 ],
   alphaCSR[ 244 ][ 197 ],
   alphaCSR[ 244 ][ 198 ],
   alphaCSR[ 244 ][ 199 ],
   alphaCSR[ 244 ][ 200 ],
   alphaCSR[ 244 ][ 201 ],
   alphaCSR[ 244 ][ 202 ],
   alphaCSR[ 244 ][ 203 ],
   alphaCSR[ 244 ][ 204 ],
   alphaCSR[ 244 ][ 205 ],
   alphaCSR[ 244 ][ 206 ],
   alphaCSR[ 244 ][ 207 ],
   alphaCSR[ 244 ][ 208 ],
   alphaCSR[ 244 ][ 209 ],
   alphaCSR[ 244 ][ 210 ],
   alphaCSR[ 244 ][ 211 ],
   alphaCSR[ 244 ][ 212 ],
   alphaCSR[ 244 ][ 213 ],
   alphaCSR[ 244 ][ 214 ],
   alphaCSR[ 244 ][ 215 ],
   alphaCSR[ 244 ][ 216 ],
   alphaCSR[ 244 ][ 217 ],
   alphaCSR[ 244 ][ 218 ],
   alphaCSR[ 244 ][ 219 ],
   alphaCSR[ 244 ][ 220 ],
   alphaCSR[ 244 ][ 221 ],
   alphaCSR[ 244 ][ 222 ],
   alphaCSR[ 244 ][ 223 ],
   alphaCSR[ 244 ][ 224 ],
   alphaCSR[ 244 ][ 225 ],
   alphaCSR[ 244 ][ 226 ],
   alphaCSR[ 244 ][ 227 ],
   alphaCSR[ 244 ][ 228 ],
   alphaCSR[ 244 ][ 229 ],
   alphaCSR[ 244 ][ 230 ],
   alphaCSR[ 244 ][ 231 ],
   alphaCSR[ 244 ][ 232 ],
   alphaCSR[ 244 ][ 233 ],
   alphaCSR[ 244 ][ 234 ],
   alphaCSR[ 244 ][ 235 ],
   alphaCSR[ 244 ][ 236 ],
   alphaCSR[ 244 ][ 237 ],
   alphaCSR[ 244 ][ 238 ],
   alphaCSR[ 244 ][ 239 ],
   alphaCSR[ 244 ][ 240 ],
   alphaCSR[ 244 ][ 241 ],
   alphaCSR[ 244 ][ 242 ],
   alphaCSR[ 244 ][ 243 ],
   alphaCSR[ 244 ][ 244 ],
   alphaCSR[ 244 ][ 245 ],
   alphaCSR[ 244 ][ 246 ],
   alphaCSR[ 244 ][ 247 ],
   alphaCSR[ 244 ][ 248 ],
   alphaCSR[ 244 ][ 249 ],
   alphaCSR[ 244 ][ 250 ],
   alphaCSR[ 244 ][ 251 ],
   alphaCSR[ 244 ][ 252 ],
   alphaCSR[ 244 ][ 253 ],
   alphaCSR[ 244 ][ 254 ],
   alphaCSR[ 244 ][ 255 ],
   alphaCSR[ 244 ][ 256 ],
   alphaCSR[ 244 ][ 257 ],
   alphaCSR[ 244 ][ 258 ],
   alphaCSR[ 244 ][ 259 ],
   alphaCSR[ 244 ][ 260 ],
   alphaCSR[ 244 ][ 261 ],
   alphaCSR[ 244 ][ 262 ],
   alphaCSR[ 244 ][ 263 ],
   alphaCSR[ 244 ][ 264 ],
   alphaCSR[ 244 ][ 265 ],
   alphaCSR[ 244 ][ 266 ],
   alphaCSR[ 244 ][ 267 ],
   alphaCSR[ 244 ][ 268 ],
   alphaCSR[ 244 ][ 269 ],
   alphaCSR[ 244 ][ 270 ],
   alphaCSR[ 244 ][ 271 ],
   alphaCSR[ 244 ][ 272 ],
   alphaCSR[ 244 ][ 273 ],
   alphaCSR[ 244 ][ 274 ],
   alphaCSR[ 244 ][ 275 ],
   alphaCSR[ 244 ][ 276 ],
   alphaCSR[ 244 ][ 277 ],
   alphaCSR[ 244 ][ 278 ],
   alphaCSR[ 244 ][ 279 ],
   alphaCSR[ 244 ][ 280 ],
   alphaCSR[ 244 ][ 281 ],
   alphaCSR[ 244 ][ 282 ],
   alphaCSR[ 244 ][ 283 ],
   alphaCSR[ 244 ][ 284 ],
   alphaCSR[ 244 ][ 285 ],
   alphaCSR[ 244 ][ 286 ],
   alphaCSR[ 244 ][ 287 ],
   alphaCSR[ 244 ][ 288 ],
   alphaCSR[ 244 ][ 289 ],
   alphaCSR[ 244 ][ 290 ],
   alphaCSR[ 244 ][ 291 ],
   alphaCSR[ 244 ][ 292 ],
   alphaCSR[ 244 ][ 293 ],
   alphaCSR[ 244 ][ 294 ],
   alphaCSR[ 244 ][ 295 ],
   alphaCSR[ 244 ][ 296 ],
   alphaCSR[ 244 ][ 297 ],
   alphaCSR[ 244 ][ 298 ],
   alphaCSR[ 244 ][ 299 ],
   alphaCSR[ 244 ][ 300 ],
   alphaCSR[ 244 ][ 301 ],
   alphaCSR[ 244 ][ 302 ],
   alphaCSR[ 244 ][ 303 ],
   alphaCSR[ 244 ][ 304 ],
   alphaCSR[ 244 ][ 305 ],
   alphaCSR[ 244 ][ 306 ],
   alphaCSR[ 244 ][ 307 ],
   alphaCSR[ 244 ][ 308 ],
   alphaCSR[ 244 ][ 309 ],
   alphaCSR[ 244 ][ 310 ],
   alphaCSR[ 244 ][ 311 ],
   alphaCSR[ 244 ][ 312 ],
   alphaCSR[ 244 ][ 313 ],
   alphaCSR[ 244 ][ 314 ],
   alphaCSR[ 244 ][ 315 ],
   alphaCSR[ 244 ][ 316 ],
   alphaCSR[ 244 ][ 317 ],
   alphaCSR[ 244 ][ 318 ],
   alphaCSR[ 244 ][ 319 ],
   alphaCSR[ 244 ][ 320 ],
   alphaCSR[ 244 ][ 321 ],
   alphaCSR[ 244 ][ 322 ],
   alphaCSR[ 244 ][ 323 ],
   alphaCSR[ 244 ][ 324 ],
   alphaCSR[ 244 ][ 325 ],
   alphaCSR[ 244 ][ 326 ],
   alphaCSR[ 244 ][ 327 ],
   alphaCSR[ 244 ][ 328 ],
   alphaCSR[ 244 ][ 329 ],
   alphaCSR[ 244 ][ 330 ],
   alphaCSR[ 244 ][ 331 ],
   alphaCSR[ 244 ][ 332 ],
   alphaCSR[ 244 ][ 333 ],
   alphaCSR[ 244 ][ 334 ],
   alphaCSR[ 244 ][ 335 ],
   alphaCSR[ 244 ][ 336 ],
   alphaCSR[ 244 ][ 337 ],
   alphaCSR[ 244 ][ 338 ],
   alphaCSR[ 244 ][ 339 ],
   alphaCSR[ 244 ][ 340 ],
   alphaCSR[ 244 ][ 341 ],
   alphaCSR[ 244 ][ 342 ],
   alphaCSR[ 244 ][ 343 ],
   alphaCSR[ 244 ][ 344 ],
   alphaCSR[ 244 ][ 345 ],
   alphaCSR[ 244 ][ 346 ],
   alphaCSR[ 244 ][ 347 ],
   alphaCSR[ 244 ][ 348 ],
   alphaCSR[ 244 ][ 349 ],
   alphaCSR[ 244 ][ 350 ],
   alphaCSR[ 244 ][ 351 ],
   alphaCSR[ 244 ][ 352 ],
   alphaCSR[ 244 ][ 353 ],
   alphaCSR[ 244 ][ 354 ],
   alphaCSR[ 244 ][ 355 ],
   alphaCSR[ 244 ][ 356 ],
   alphaCSR[ 244 ][ 357 ],
   alphaCSR[ 244 ][ 358 ],
   alphaCSR[ 244 ][ 359 ],
   alphaCSR[ 244 ][ 360 ],
   alphaCSR[ 244 ][ 361 ],
   alphaCSR[ 244 ][ 362 ],
   alphaCSR[ 244 ][ 363 ],
   alphaCSR[ 244 ][ 364 ],
   alphaCSR[ 244 ][ 365 ],
   alphaCSR[ 244 ][ 366 ],
   alphaCSR[ 244 ][ 367 ],
   alphaCSR[ 244 ][ 368 ],
   alphaCSR[ 244 ][ 369 ],
   alphaCSR[ 244 ][ 370 ],
   alphaCSR[ 244 ][ 371 ],
   alphaCSR[ 244 ][ 372 ],
   alphaCSR[ 244 ][ 373 ],
   alphaCSR[ 244 ][ 374 ],
   alphaCSR[ 244 ][ 375 ],
   alphaCSR[ 244 ][ 376 ],
   alphaCSR[ 244 ][ 377 ],
   alphaCSR[ 244 ][ 378 ],
   alphaCSR[ 244 ][ 379 ],
   alphaCSR[ 244 ][ 380 ],
   alphaCSR[ 244 ][ 381 ],
   alphaCSR[ 244 ][ 382 ],
   alphaCSR[ 244 ][ 383 ],
   alphaCSR[ 245 ][ 0 ],
   alphaCSR[ 245 ][ 1 ],
   alphaCSR[ 245 ][ 2 ],
   alphaCSR[ 245 ][ 3 ],
   alphaCSR[ 245 ][ 4 ],
   alphaCSR[ 245 ][ 5 ],
   alphaCSR[ 245 ][ 6 ],
   alphaCSR[ 245 ][ 7 ],
   alphaCSR[ 245 ][ 8 ],
   alphaCSR[ 245 ][ 9 ],
   alphaCSR[ 245 ][ 10 ],
   alphaCSR[ 245 ][ 11 ],
   alphaCSR[ 245 ][ 12 ],
   alphaCSR[ 245 ][ 13 ],
   alphaCSR[ 245 ][ 14 ],
   alphaCSR[ 245 ][ 15 ],
   alphaCSR[ 245 ][ 16 ],
   alphaCSR[ 245 ][ 17 ],
   alphaCSR[ 245 ][ 18 ],
   alphaCSR[ 245 ][ 19 ],
   alphaCSR[ 245 ][ 20 ],
   alphaCSR[ 245 ][ 21 ],
   alphaCSR[ 245 ][ 22 ],
   alphaCSR[ 245 ][ 23 ],
   alphaCSR[ 245 ][ 24 ],
   alphaCSR[ 245 ][ 25 ],
   alphaCSR[ 245 ][ 26 ],
   alphaCSR[ 245 ][ 27 ],
   alphaCSR[ 245 ][ 28 ],
   alphaCSR[ 245 ][ 29 ],
   alphaCSR[ 245 ][ 30 ],
   alphaCSR[ 245 ][ 31 ],
   alphaCSR[ 245 ][ 32 ],
   alphaCSR[ 245 ][ 33 ],
   alphaCSR[ 245 ][ 34 ],
   alphaCSR[ 245 ][ 35 ],
   alphaCSR[ 245 ][ 36 ],
   alphaCSR[ 245 ][ 37 ],
   alphaCSR[ 245 ][ 38 ],
   alphaCSR[ 245 ][ 39 ],
   alphaCSR[ 245 ][ 40 ],
   alphaCSR[ 245 ][ 41 ],
   alphaCSR[ 245 ][ 42 ],
   alphaCSR[ 245 ][ 43 ],
   alphaCSR[ 245 ][ 44 ],
   alphaCSR[ 245 ][ 45 ],
   alphaCSR[ 245 ][ 46 ],
   alphaCSR[ 245 ][ 47 ],
   alphaCSR[ 245 ][ 48 ],
   alphaCSR[ 245 ][ 49 ],
   alphaCSR[ 245 ][ 50 ],
   alphaCSR[ 245 ][ 51 ],
   alphaCSR[ 245 ][ 52 ],
   alphaCSR[ 245 ][ 53 ],
   alphaCSR[ 245 ][ 54 ],
   alphaCSR[ 245 ][ 55 ],
   alphaCSR[ 245 ][ 56 ],
   alphaCSR[ 245 ][ 57 ],
   alphaCSR[ 245 ][ 58 ],
   alphaCSR[ 245 ][ 59 ],
   alphaCSR[ 245 ][ 60 ],
   alphaCSR[ 245 ][ 61 ],
   alphaCSR[ 245 ][ 62 ],
   alphaCSR[ 245 ][ 63 ],
   alphaCSR[ 245 ][ 64 ],
   alphaCSR[ 245 ][ 65 ],
   alphaCSR[ 245 ][ 66 ],
   alphaCSR[ 245 ][ 67 ],
   alphaCSR[ 245 ][ 68 ],
   alphaCSR[ 245 ][ 69 ],
   alphaCSR[ 245 ][ 70 ],
   alphaCSR[ 245 ][ 71 ],
   alphaCSR[ 245 ][ 72 ],
   alphaCSR[ 245 ][ 73 ],
   alphaCSR[ 245 ][ 74 ],
   alphaCSR[ 245 ][ 75 ],
   alphaCSR[ 245 ][ 76 ],
   alphaCSR[ 245 ][ 77 ],
   alphaCSR[ 245 ][ 78 ],
   alphaCSR[ 245 ][ 79 ],
   alphaCSR[ 245 ][ 80 ],
   alphaCSR[ 245 ][ 81 ],
   alphaCSR[ 245 ][ 82 ],
   alphaCSR[ 245 ][ 83 ],
   alphaCSR[ 245 ][ 84 ],
   alphaCSR[ 245 ][ 85 ],
   alphaCSR[ 245 ][ 86 ],
   alphaCSR[ 245 ][ 87 ],
   alphaCSR[ 245 ][ 88 ],
   alphaCSR[ 245 ][ 89 ],
   alphaCSR[ 245 ][ 90 ],
   alphaCSR[ 245 ][ 91 ],
   alphaCSR[ 245 ][ 92 ],
   alphaCSR[ 245 ][ 93 ],
   alphaCSR[ 245 ][ 94 ],
   alphaCSR[ 245 ][ 95 ],
   alphaCSR[ 245 ][ 96 ],
   alphaCSR[ 245 ][ 97 ],
   alphaCSR[ 245 ][ 98 ],
   alphaCSR[ 245 ][ 99 ],
   alphaCSR[ 245 ][ 100 ],
   alphaCSR[ 245 ][ 101 ],
   alphaCSR[ 245 ][ 102 ],
   alphaCSR[ 245 ][ 103 ],
   alphaCSR[ 245 ][ 104 ],
   alphaCSR[ 245 ][ 105 ],
   alphaCSR[ 245 ][ 106 ],
   alphaCSR[ 245 ][ 107 ],
   alphaCSR[ 245 ][ 108 ],
   alphaCSR[ 245 ][ 109 ],
   alphaCSR[ 245 ][ 110 ],
   alphaCSR[ 245 ][ 111 ],
   alphaCSR[ 245 ][ 112 ],
   alphaCSR[ 245 ][ 113 ],
   alphaCSR[ 245 ][ 114 ],
   alphaCSR[ 245 ][ 115 ],
   alphaCSR[ 245 ][ 116 ],
   alphaCSR[ 245 ][ 117 ],
   alphaCSR[ 245 ][ 118 ],
   alphaCSR[ 245 ][ 119 ],
   alphaCSR[ 245 ][ 120 ],
   alphaCSR[ 245 ][ 121 ],
   alphaCSR[ 245 ][ 122 ],
   alphaCSR[ 245 ][ 123 ],
   alphaCSR[ 245 ][ 124 ],
   alphaCSR[ 245 ][ 125 ],
   alphaCSR[ 245 ][ 126 ],
   alphaCSR[ 245 ][ 127 ],
   alphaCSR[ 245 ][ 128 ],
   alphaCSR[ 245 ][ 129 ],
   alphaCSR[ 245 ][ 130 ],
   alphaCSR[ 245 ][ 131 ],
   alphaCSR[ 245 ][ 132 ],
   alphaCSR[ 245 ][ 133 ],
   alphaCSR[ 245 ][ 134 ],
   alphaCSR[ 245 ][ 135 ],
   alphaCSR[ 245 ][ 136 ],
   alphaCSR[ 245 ][ 137 ],
   alphaCSR[ 245 ][ 138 ],
   alphaCSR[ 245 ][ 139 ],
   alphaCSR[ 245 ][ 140 ],
   alphaCSR[ 245 ][ 141 ],
   alphaCSR[ 245 ][ 142 ],
   alphaCSR[ 245 ][ 143 ],
   alphaCSR[ 245 ][ 144 ],
   alphaCSR[ 245 ][ 145 ],
   alphaCSR[ 245 ][ 146 ],
   alphaCSR[ 245 ][ 147 ],
   alphaCSR[ 245 ][ 148 ],
   alphaCSR[ 245 ][ 149 ],
   alphaCSR[ 245 ][ 150 ],
   alphaCSR[ 245 ][ 151 ],
   alphaCSR[ 245 ][ 152 ],
   alphaCSR[ 245 ][ 153 ],
   alphaCSR[ 245 ][ 154 ],
   alphaCSR[ 245 ][ 155 ],
   alphaCSR[ 245 ][ 156 ],
   alphaCSR[ 245 ][ 157 ],
   alphaCSR[ 245 ][ 158 ],
   alphaCSR[ 245 ][ 159 ],
   alphaCSR[ 245 ][ 160 ],
   alphaCSR[ 245 ][ 161 ],
   alphaCSR[ 245 ][ 162 ],
   alphaCSR[ 245 ][ 163 ],
   alphaCSR[ 245 ][ 164 ],
   alphaCSR[ 245 ][ 165 ],
   alphaCSR[ 245 ][ 166 ],
   alphaCSR[ 245 ][ 167 ],
   alphaCSR[ 245 ][ 168 ],
   alphaCSR[ 245 ][ 169 ],
   alphaCSR[ 245 ][ 170 ],
   alphaCSR[ 245 ][ 171 ],
   alphaCSR[ 245 ][ 172 ],
   alphaCSR[ 245 ][ 173 ],
   alphaCSR[ 245 ][ 174 ],
   alphaCSR[ 245 ][ 175 ],
   alphaCSR[ 245 ][ 176 ],
   alphaCSR[ 245 ][ 177 ],
   alphaCSR[ 245 ][ 178 ],
   alphaCSR[ 245 ][ 179 ],
   alphaCSR[ 245 ][ 180 ],
   alphaCSR[ 245 ][ 181 ],
   alphaCSR[ 245 ][ 182 ],
   alphaCSR[ 245 ][ 183 ],
   alphaCSR[ 245 ][ 184 ],
   alphaCSR[ 245 ][ 185 ],
   alphaCSR[ 245 ][ 186 ],
   alphaCSR[ 245 ][ 187 ],
   alphaCSR[ 245 ][ 188 ],
   alphaCSR[ 245 ][ 189 ],
   alphaCSR[ 245 ][ 190 ],
   alphaCSR[ 245 ][ 191 ],
   alphaCSR[ 245 ][ 192 ],
   alphaCSR[ 245 ][ 193 ],
   alphaCSR[ 245 ][ 194 ],
   alphaCSR[ 245 ][ 195 ],
   alphaCSR[ 245 ][ 196 ],
   alphaCSR[ 245 ][ 197 ],
   alphaCSR[ 245 ][ 198 ],
   alphaCSR[ 245 ][ 199 ],
   alphaCSR[ 245 ][ 200 ],
   alphaCSR[ 245 ][ 201 ],
   alphaCSR[ 245 ][ 202 ],
   alphaCSR[ 245 ][ 203 ],
   alphaCSR[ 245 ][ 204 ],
   alphaCSR[ 245 ][ 205 ],
   alphaCSR[ 245 ][ 206 ],
   alphaCSR[ 245 ][ 207 ],
   alphaCSR[ 245 ][ 208 ],
   alphaCSR[ 245 ][ 209 ],
   alphaCSR[ 245 ][ 210 ],
   alphaCSR[ 245 ][ 211 ],
   alphaCSR[ 245 ][ 212 ],
   alphaCSR[ 245 ][ 213 ],
   alphaCSR[ 245 ][ 214 ],
   alphaCSR[ 245 ][ 215 ],
   alphaCSR[ 245 ][ 216 ],
   alphaCSR[ 245 ][ 217 ],
   alphaCSR[ 245 ][ 218 ],
   alphaCSR[ 245 ][ 219 ],
   alphaCSR[ 245 ][ 220 ],
   alphaCSR[ 245 ][ 221 ],
   alphaCSR[ 245 ][ 222 ],
   alphaCSR[ 245 ][ 223 ],
   alphaCSR[ 245 ][ 224 ],
   alphaCSR[ 245 ][ 225 ],
   alphaCSR[ 245 ][ 226 ],
   alphaCSR[ 245 ][ 227 ],
   alphaCSR[ 245 ][ 228 ],
   alphaCSR[ 245 ][ 229 ],
   alphaCSR[ 245 ][ 230 ],
   alphaCSR[ 245 ][ 231 ],
   alphaCSR[ 245 ][ 232 ],
   alphaCSR[ 245 ][ 233 ],
   alphaCSR[ 245 ][ 234 ],
   alphaCSR[ 245 ][ 235 ],
   alphaCSR[ 245 ][ 236 ],
   alphaCSR[ 245 ][ 237 ],
   alphaCSR[ 245 ][ 238 ],
   alphaCSR[ 245 ][ 239 ],
   alphaCSR[ 245 ][ 240 ],
   alphaCSR[ 245 ][ 241 ],
   alphaCSR[ 245 ][ 242 ],
   alphaCSR[ 245 ][ 243 ],
   alphaCSR[ 245 ][ 244 ],
   alphaCSR[ 245 ][ 245 ],
   alphaCSR[ 245 ][ 246 ],
   alphaCSR[ 245 ][ 247 ],
   alphaCSR[ 245 ][ 248 ],
   alphaCSR[ 245 ][ 249 ],
   alphaCSR[ 245 ][ 250 ],
   alphaCSR[ 245 ][ 251 ],
   alphaCSR[ 245 ][ 252 ],
   alphaCSR[ 245 ][ 253 ],
   alphaCSR[ 245 ][ 254 ],
   alphaCSR[ 245 ][ 255 ],
   alphaCSR[ 245 ][ 256 ],
   alphaCSR[ 245 ][ 257 ],
   alphaCSR[ 245 ][ 258 ],
   alphaCSR[ 245 ][ 259 ],
   alphaCSR[ 245 ][ 260 ],
   alphaCSR[ 245 ][ 261 ],
   alphaCSR[ 245 ][ 262 ],
   alphaCSR[ 245 ][ 263 ],
   alphaCSR[ 245 ][ 264 ],
   alphaCSR[ 245 ][ 265 ],
   alphaCSR[ 245 ][ 266 ],
   alphaCSR[ 245 ][ 267 ],
   alphaCSR[ 245 ][ 268 ],
   alphaCSR[ 245 ][ 269 ],
   alphaCSR[ 245 ][ 270 ],
   alphaCSR[ 245 ][ 271 ],
   alphaCSR[ 245 ][ 272 ],
   alphaCSR[ 245 ][ 273 ],
   alphaCSR[ 245 ][ 274 ],
   alphaCSR[ 245 ][ 275 ],
   alphaCSR[ 245 ][ 276 ],
   alphaCSR[ 245 ][ 277 ],
   alphaCSR[ 245 ][ 278 ],
   alphaCSR[ 245 ][ 279 ],
   alphaCSR[ 245 ][ 280 ],
   alphaCSR[ 245 ][ 281 ],
   alphaCSR[ 245 ][ 282 ],
   alphaCSR[ 245 ][ 283 ],
   alphaCSR[ 245 ][ 284 ],
   alphaCSR[ 245 ][ 285 ],
   alphaCSR[ 245 ][ 286 ],
   alphaCSR[ 245 ][ 287 ],
   alphaCSR[ 245 ][ 288 ],
   alphaCSR[ 245 ][ 289 ],
   alphaCSR[ 245 ][ 290 ],
   alphaCSR[ 245 ][ 291 ],
   alphaCSR[ 245 ][ 292 ],
   alphaCSR[ 245 ][ 293 ],
   alphaCSR[ 245 ][ 294 ],
   alphaCSR[ 245 ][ 295 ],
   alphaCSR[ 245 ][ 296 ],
   alphaCSR[ 245 ][ 297 ],
   alphaCSR[ 245 ][ 298 ],
   alphaCSR[ 245 ][ 299 ],
   alphaCSR[ 245 ][ 300 ],
   alphaCSR[ 245 ][ 301 ],
   alphaCSR[ 245 ][ 302 ],
   alphaCSR[ 245 ][ 303 ],
   alphaCSR[ 245 ][ 304 ],
   alphaCSR[ 245 ][ 305 ],
   alphaCSR[ 245 ][ 306 ],
   alphaCSR[ 245 ][ 307 ],
   alphaCSR[ 245 ][ 308 ],
   alphaCSR[ 245 ][ 309 ],
   alphaCSR[ 245 ][ 310 ],
   alphaCSR[ 245 ][ 311 ],
   alphaCSR[ 245 ][ 312 ],
   alphaCSR[ 245 ][ 313 ],
   alphaCSR[ 245 ][ 314 ],
   alphaCSR[ 245 ][ 315 ],
   alphaCSR[ 245 ][ 316 ],
   alphaCSR[ 245 ][ 317 ],
   alphaCSR[ 245 ][ 318 ],
   alphaCSR[ 245 ][ 319 ],
   alphaCSR[ 245 ][ 320 ],
   alphaCSR[ 245 ][ 321 ],
   alphaCSR[ 245 ][ 322 ],
   alphaCSR[ 245 ][ 323 ],
   alphaCSR[ 245 ][ 324 ],
   alphaCSR[ 245 ][ 325 ],
   alphaCSR[ 245 ][ 326 ],
   alphaCSR[ 245 ][ 327 ],
   alphaCSR[ 245 ][ 328 ],
   alphaCSR[ 245 ][ 329 ],
   alphaCSR[ 245 ][ 330 ],
   alphaCSR[ 245 ][ 331 ],
   alphaCSR[ 245 ][ 332 ],
   alphaCSR[ 245 ][ 333 ],
   alphaCSR[ 245 ][ 334 ],
   alphaCSR[ 245 ][ 335 ],
   alphaCSR[ 245 ][ 336 ],
   alphaCSR[ 245 ][ 337 ],
   alphaCSR[ 245 ][ 338 ],
   alphaCSR[ 245 ][ 339 ],
   alphaCSR[ 245 ][ 340 ],
   alphaCSR[ 245 ][ 341 ],
   alphaCSR[ 245 ][ 342 ],
   alphaCSR[ 245 ][ 343 ],
   alphaCSR[ 245 ][ 344 ],
   alphaCSR[ 245 ][ 345 ],
   alphaCSR[ 245 ][ 346 ],
   alphaCSR[ 245 ][ 347 ],
   alphaCSR[ 245 ][ 348 ],
   alphaCSR[ 245 ][ 349 ],
   alphaCSR[ 245 ][ 350 ],
   alphaCSR[ 245 ][ 351 ],
   alphaCSR[ 245 ][ 352 ],
   alphaCSR[ 245 ][ 353 ],
   alphaCSR[ 245 ][ 354 ],
   alphaCSR[ 245 ][ 355 ],
   alphaCSR[ 245 ][ 356 ],
   alphaCSR[ 245 ][ 357 ],
   alphaCSR[ 245 ][ 358 ],
   alphaCSR[ 245 ][ 359 ],
   alphaCSR[ 245 ][ 360 ],
   alphaCSR[ 245 ][ 361 ],
   alphaCSR[ 245 ][ 362 ],
   alphaCSR[ 245 ][ 363 ],
   alphaCSR[ 245 ][ 364 ],
   alphaCSR[ 245 ][ 365 ],
   alphaCSR[ 245 ][ 366 ],
   alphaCSR[ 245 ][ 367 ],
   alphaCSR[ 245 ][ 368 ],
   alphaCSR[ 245 ][ 369 ],
   alphaCSR[ 245 ][ 370 ],
   alphaCSR[ 245 ][ 371 ],
   alphaCSR[ 245 ][ 372 ],
   alphaCSR[ 245 ][ 373 ],
   alphaCSR[ 245 ][ 374 ],
   alphaCSR[ 245 ][ 375 ],
   alphaCSR[ 245 ][ 376 ],
   alphaCSR[ 245 ][ 377 ],
   alphaCSR[ 245 ][ 378 ],
   alphaCSR[ 245 ][ 379 ],
   alphaCSR[ 245 ][ 380 ],
   alphaCSR[ 245 ][ 381 ],
   alphaCSR[ 245 ][ 382 ],
   alphaCSR[ 245 ][ 383 ],
   alphaCSR[ 246 ][ 0 ],
   alphaCSR[ 246 ][ 1 ],
   alphaCSR[ 246 ][ 2 ],
   alphaCSR[ 246 ][ 3 ],
   alphaCSR[ 246 ][ 4 ],
   alphaCSR[ 246 ][ 5 ],
   alphaCSR[ 246 ][ 6 ],
   alphaCSR[ 246 ][ 7 ],
   alphaCSR[ 246 ][ 8 ],
   alphaCSR[ 246 ][ 9 ],
   alphaCSR[ 246 ][ 10 ],
   alphaCSR[ 246 ][ 11 ],
   alphaCSR[ 246 ][ 12 ],
   alphaCSR[ 246 ][ 13 ],
   alphaCSR[ 246 ][ 14 ],
   alphaCSR[ 246 ][ 15 ],
   alphaCSR[ 246 ][ 16 ],
   alphaCSR[ 246 ][ 17 ],
   alphaCSR[ 246 ][ 18 ],
   alphaCSR[ 246 ][ 19 ],
   alphaCSR[ 246 ][ 20 ],
   alphaCSR[ 246 ][ 21 ],
   alphaCSR[ 246 ][ 22 ],
   alphaCSR[ 246 ][ 23 ],
   alphaCSR[ 246 ][ 24 ],
   alphaCSR[ 246 ][ 25 ],
   alphaCSR[ 246 ][ 26 ],
   alphaCSR[ 246 ][ 27 ],
   alphaCSR[ 246 ][ 28 ],
   alphaCSR[ 246 ][ 29 ],
   alphaCSR[ 246 ][ 30 ],
   alphaCSR[ 246 ][ 31 ],
   alphaCSR[ 246 ][ 32 ],
   alphaCSR[ 246 ][ 33 ],
   alphaCSR[ 246 ][ 34 ],
   alphaCSR[ 246 ][ 35 ],
   alphaCSR[ 246 ][ 36 ],
   alphaCSR[ 246 ][ 37 ],
   alphaCSR[ 246 ][ 38 ],
   alphaCSR[ 246 ][ 39 ],
   alphaCSR[ 246 ][ 40 ],
   alphaCSR[ 246 ][ 41 ],
   alphaCSR[ 246 ][ 42 ],
   alphaCSR[ 246 ][ 43 ],
   alphaCSR[ 246 ][ 44 ],
   alphaCSR[ 246 ][ 45 ],
   alphaCSR[ 246 ][ 46 ],
   alphaCSR[ 246 ][ 47 ],
   alphaCSR[ 246 ][ 48 ],
   alphaCSR[ 246 ][ 49 ],
   alphaCSR[ 246 ][ 50 ],
   alphaCSR[ 246 ][ 51 ],
   alphaCSR[ 246 ][ 52 ],
   alphaCSR[ 246 ][ 53 ],
   alphaCSR[ 246 ][ 54 ],
   alphaCSR[ 246 ][ 55 ],
   alphaCSR[ 246 ][ 56 ],
   alphaCSR[ 246 ][ 57 ],
   alphaCSR[ 246 ][ 58 ],
   alphaCSR[ 246 ][ 59 ],
   alphaCSR[ 246 ][ 60 ],
   alphaCSR[ 246 ][ 61 ],
   alphaCSR[ 246 ][ 62 ],
   alphaCSR[ 246 ][ 63 ],
   alphaCSR[ 246 ][ 64 ],
   alphaCSR[ 246 ][ 65 ],
   alphaCSR[ 246 ][ 66 ],
   alphaCSR[ 246 ][ 67 ],
   alphaCSR[ 246 ][ 68 ],
   alphaCSR[ 246 ][ 69 ],
   alphaCSR[ 246 ][ 70 ],
   alphaCSR[ 246 ][ 71 ],
   alphaCSR[ 246 ][ 72 ],
   alphaCSR[ 246 ][ 73 ],
   alphaCSR[ 246 ][ 74 ],
   alphaCSR[ 246 ][ 75 ],
   alphaCSR[ 246 ][ 76 ],
   alphaCSR[ 246 ][ 77 ],
   alphaCSR[ 246 ][ 78 ],
   alphaCSR[ 246 ][ 79 ],
   alphaCSR[ 246 ][ 80 ],
   alphaCSR[ 246 ][ 81 ],
   alphaCSR[ 246 ][ 82 ],
   alphaCSR[ 246 ][ 83 ],
   alphaCSR[ 246 ][ 84 ],
   alphaCSR[ 246 ][ 85 ],
   alphaCSR[ 246 ][ 86 ],
   alphaCSR[ 246 ][ 87 ],
   alphaCSR[ 246 ][ 88 ],
   alphaCSR[ 246 ][ 89 ],
   alphaCSR[ 246 ][ 90 ],
   alphaCSR[ 246 ][ 91 ],
   alphaCSR[ 246 ][ 92 ],
   alphaCSR[ 246 ][ 93 ],
   alphaCSR[ 246 ][ 94 ],
   alphaCSR[ 246 ][ 95 ],
   alphaCSR[ 246 ][ 96 ],
   alphaCSR[ 246 ][ 97 ],
   alphaCSR[ 246 ][ 98 ],
   alphaCSR[ 246 ][ 99 ],
   alphaCSR[ 246 ][ 100 ],
   alphaCSR[ 246 ][ 101 ],
   alphaCSR[ 246 ][ 102 ],
   alphaCSR[ 246 ][ 103 ],
   alphaCSR[ 246 ][ 104 ],
   alphaCSR[ 246 ][ 105 ],
   alphaCSR[ 246 ][ 106 ],
   alphaCSR[ 246 ][ 107 ],
   alphaCSR[ 246 ][ 108 ],
   alphaCSR[ 246 ][ 109 ],
   alphaCSR[ 246 ][ 110 ],
   alphaCSR[ 246 ][ 111 ],
   alphaCSR[ 246 ][ 112 ],
   alphaCSR[ 246 ][ 113 ],
   alphaCSR[ 246 ][ 114 ],
   alphaCSR[ 246 ][ 115 ],
   alphaCSR[ 246 ][ 116 ],
   alphaCSR[ 246 ][ 117 ],
   alphaCSR[ 246 ][ 118 ],
   alphaCSR[ 246 ][ 119 ],
   alphaCSR[ 246 ][ 120 ],
   alphaCSR[ 246 ][ 121 ],
   alphaCSR[ 246 ][ 122 ],
   alphaCSR[ 246 ][ 123 ],
   alphaCSR[ 246 ][ 124 ],
   alphaCSR[ 246 ][ 125 ],
   alphaCSR[ 246 ][ 126 ],
   alphaCSR[ 246 ][ 127 ],
   alphaCSR[ 246 ][ 128 ],
   alphaCSR[ 246 ][ 129 ],
   alphaCSR[ 246 ][ 130 ],
   alphaCSR[ 246 ][ 131 ],
   alphaCSR[ 246 ][ 132 ],
   alphaCSR[ 246 ][ 133 ],
   alphaCSR[ 246 ][ 134 ],
   alphaCSR[ 246 ][ 135 ],
   alphaCSR[ 246 ][ 136 ],
   alphaCSR[ 246 ][ 137 ],
   alphaCSR[ 246 ][ 138 ],
   alphaCSR[ 246 ][ 139 ],
   alphaCSR[ 246 ][ 140 ],
   alphaCSR[ 246 ][ 141 ],
   alphaCSR[ 246 ][ 142 ],
   alphaCSR[ 246 ][ 143 ],
   alphaCSR[ 246 ][ 144 ],
   alphaCSR[ 246 ][ 145 ],
   alphaCSR[ 246 ][ 146 ],
   alphaCSR[ 246 ][ 147 ],
   alphaCSR[ 246 ][ 148 ],
   alphaCSR[ 246 ][ 149 ],
   alphaCSR[ 246 ][ 150 ],
   alphaCSR[ 246 ][ 151 ],
   alphaCSR[ 246 ][ 152 ],
   alphaCSR[ 246 ][ 153 ],
   alphaCSR[ 246 ][ 154 ],
   alphaCSR[ 246 ][ 155 ],
   alphaCSR[ 246 ][ 156 ],
   alphaCSR[ 246 ][ 157 ],
   alphaCSR[ 246 ][ 158 ],
   alphaCSR[ 246 ][ 159 ],
   alphaCSR[ 246 ][ 160 ],
   alphaCSR[ 246 ][ 161 ],
   alphaCSR[ 246 ][ 162 ],
   alphaCSR[ 246 ][ 163 ],
   alphaCSR[ 246 ][ 164 ],
   alphaCSR[ 246 ][ 165 ],
   alphaCSR[ 246 ][ 166 ],
   alphaCSR[ 246 ][ 167 ],
   alphaCSR[ 246 ][ 168 ],
   alphaCSR[ 246 ][ 169 ],
   alphaCSR[ 246 ][ 170 ],
   alphaCSR[ 246 ][ 171 ],
   alphaCSR[ 246 ][ 172 ],
   alphaCSR[ 246 ][ 173 ],
   alphaCSR[ 246 ][ 174 ],
   alphaCSR[ 246 ][ 175 ],
   alphaCSR[ 246 ][ 176 ],
   alphaCSR[ 246 ][ 177 ],
   alphaCSR[ 246 ][ 178 ],
   alphaCSR[ 246 ][ 179 ],
   alphaCSR[ 246 ][ 180 ],
   alphaCSR[ 246 ][ 181 ],
   alphaCSR[ 246 ][ 182 ],
   alphaCSR[ 246 ][ 183 ],
   alphaCSR[ 246 ][ 184 ],
   alphaCSR[ 246 ][ 185 ],
   alphaCSR[ 246 ][ 186 ],
   alphaCSR[ 246 ][ 187 ],
   alphaCSR[ 246 ][ 188 ],
   alphaCSR[ 246 ][ 189 ],
   alphaCSR[ 246 ][ 190 ],
   alphaCSR[ 246 ][ 191 ],
   alphaCSR[ 246 ][ 192 ],
   alphaCSR[ 246 ][ 193 ],
   alphaCSR[ 246 ][ 194 ],
   alphaCSR[ 246 ][ 195 ],
   alphaCSR[ 246 ][ 196 ],
   alphaCSR[ 246 ][ 197 ],
   alphaCSR[ 246 ][ 198 ],
   alphaCSR[ 246 ][ 199 ],
   alphaCSR[ 246 ][ 200 ],
   alphaCSR[ 246 ][ 201 ],
   alphaCSR[ 246 ][ 202 ],
   alphaCSR[ 246 ][ 203 ],
   alphaCSR[ 246 ][ 204 ],
   alphaCSR[ 246 ][ 205 ],
   alphaCSR[ 246 ][ 206 ],
   alphaCSR[ 246 ][ 207 ],
   alphaCSR[ 246 ][ 208 ],
   alphaCSR[ 246 ][ 209 ],
   alphaCSR[ 246 ][ 210 ],
   alphaCSR[ 246 ][ 211 ],
   alphaCSR[ 246 ][ 212 ],
   alphaCSR[ 246 ][ 213 ],
   alphaCSR[ 246 ][ 214 ],
   alphaCSR[ 246 ][ 215 ],
   alphaCSR[ 246 ][ 216 ],
   alphaCSR[ 246 ][ 217 ],
   alphaCSR[ 246 ][ 218 ],
   alphaCSR[ 246 ][ 219 ],
   alphaCSR[ 246 ][ 220 ],
   alphaCSR[ 246 ][ 221 ],
   alphaCSR[ 246 ][ 222 ],
   alphaCSR[ 246 ][ 223 ],
   alphaCSR[ 246 ][ 224 ],
   alphaCSR[ 246 ][ 225 ],
   alphaCSR[ 246 ][ 226 ],
   alphaCSR[ 246 ][ 227 ],
   alphaCSR[ 246 ][ 228 ],
   alphaCSR[ 246 ][ 229 ],
   alphaCSR[ 246 ][ 230 ],
   alphaCSR[ 246 ][ 231 ],
   alphaCSR[ 246 ][ 232 ],
   alphaCSR[ 246 ][ 233 ],
   alphaCSR[ 246 ][ 234 ],
   alphaCSR[ 246 ][ 235 ],
   alphaCSR[ 246 ][ 236 ],
   alphaCSR[ 246 ][ 237 ],
   alphaCSR[ 246 ][ 238 ],
   alphaCSR[ 246 ][ 239 ],
   alphaCSR[ 246 ][ 240 ],
   alphaCSR[ 246 ][ 241 ],
   alphaCSR[ 246 ][ 242 ],
   alphaCSR[ 246 ][ 243 ],
   alphaCSR[ 246 ][ 244 ],
   alphaCSR[ 246 ][ 245 ],
   alphaCSR[ 246 ][ 246 ],
   alphaCSR[ 246 ][ 247 ],
   alphaCSR[ 246 ][ 248 ],
   alphaCSR[ 246 ][ 249 ],
   alphaCSR[ 246 ][ 250 ],
   alphaCSR[ 246 ][ 251 ],
   alphaCSR[ 246 ][ 252 ],
   alphaCSR[ 246 ][ 253 ],
   alphaCSR[ 246 ][ 254 ],
   alphaCSR[ 246 ][ 255 ],
   alphaCSR[ 246 ][ 256 ],
   alphaCSR[ 246 ][ 257 ],
   alphaCSR[ 246 ][ 258 ],
   alphaCSR[ 246 ][ 259 ],
   alphaCSR[ 246 ][ 260 ],
   alphaCSR[ 246 ][ 261 ],
   alphaCSR[ 246 ][ 262 ],
   alphaCSR[ 246 ][ 263 ],
   alphaCSR[ 246 ][ 264 ],
   alphaCSR[ 246 ][ 265 ],
   alphaCSR[ 246 ][ 266 ],
   alphaCSR[ 246 ][ 267 ],
   alphaCSR[ 246 ][ 268 ],
   alphaCSR[ 246 ][ 269 ],
   alphaCSR[ 246 ][ 270 ],
   alphaCSR[ 246 ][ 271 ],
   alphaCSR[ 246 ][ 272 ],
   alphaCSR[ 246 ][ 273 ],
   alphaCSR[ 246 ][ 274 ],
   alphaCSR[ 246 ][ 275 ],
   alphaCSR[ 246 ][ 276 ],
   alphaCSR[ 246 ][ 277 ],
   alphaCSR[ 246 ][ 278 ],
   alphaCSR[ 246 ][ 279 ],
   alphaCSR[ 246 ][ 280 ],
   alphaCSR[ 246 ][ 281 ],
   alphaCSR[ 246 ][ 282 ],
   alphaCSR[ 246 ][ 283 ],
   alphaCSR[ 246 ][ 284 ],
   alphaCSR[ 246 ][ 285 ],
   alphaCSR[ 246 ][ 286 ],
   alphaCSR[ 246 ][ 287 ],
   alphaCSR[ 246 ][ 288 ],
   alphaCSR[ 246 ][ 289 ],
   alphaCSR[ 246 ][ 290 ],
   alphaCSR[ 246 ][ 291 ],
   alphaCSR[ 246 ][ 292 ],
   alphaCSR[ 246 ][ 293 ],
   alphaCSR[ 246 ][ 294 ],
   alphaCSR[ 246 ][ 295 ],
   alphaCSR[ 246 ][ 296 ],
   alphaCSR[ 246 ][ 297 ],
   alphaCSR[ 246 ][ 298 ],
   alphaCSR[ 246 ][ 299 ],
   alphaCSR[ 246 ][ 300 ],
   alphaCSR[ 246 ][ 301 ],
   alphaCSR[ 246 ][ 302 ],
   alphaCSR[ 246 ][ 303 ],
   alphaCSR[ 246 ][ 304 ],
   alphaCSR[ 246 ][ 305 ],
   alphaCSR[ 246 ][ 306 ],
   alphaCSR[ 246 ][ 307 ],
   alphaCSR[ 246 ][ 308 ],
   alphaCSR[ 246 ][ 309 ],
   alphaCSR[ 246 ][ 310 ],
   alphaCSR[ 246 ][ 311 ],
   alphaCSR[ 246 ][ 312 ],
   alphaCSR[ 246 ][ 313 ],
   alphaCSR[ 246 ][ 314 ],
   alphaCSR[ 246 ][ 315 ],
   alphaCSR[ 246 ][ 316 ],
   alphaCSR[ 246 ][ 317 ],
   alphaCSR[ 246 ][ 318 ],
   alphaCSR[ 246 ][ 319 ],
   alphaCSR[ 246 ][ 320 ],
   alphaCSR[ 246 ][ 321 ],
   alphaCSR[ 246 ][ 322 ],
   alphaCSR[ 246 ][ 323 ],
   alphaCSR[ 246 ][ 324 ],
   alphaCSR[ 246 ][ 325 ],
   alphaCSR[ 246 ][ 326 ],
   alphaCSR[ 246 ][ 327 ],
   alphaCSR[ 246 ][ 328 ],
   alphaCSR[ 246 ][ 329 ],
   alphaCSR[ 246 ][ 330 ],
   alphaCSR[ 246 ][ 331 ],
   alphaCSR[ 246 ][ 332 ],
   alphaCSR[ 246 ][ 333 ],
   alphaCSR[ 246 ][ 334 ],
   alphaCSR[ 246 ][ 335 ],
   alphaCSR[ 246 ][ 336 ],
   alphaCSR[ 246 ][ 337 ],
   alphaCSR[ 246 ][ 338 ],
   alphaCSR[ 246 ][ 339 ],
   alphaCSR[ 246 ][ 340 ],
   alphaCSR[ 246 ][ 341 ],
   alphaCSR[ 246 ][ 342 ],
   alphaCSR[ 246 ][ 343 ],
   alphaCSR[ 246 ][ 344 ],
   alphaCSR[ 246 ][ 345 ],
   alphaCSR[ 246 ][ 346 ],
   alphaCSR[ 246 ][ 347 ],
   alphaCSR[ 246 ][ 348 ],
   alphaCSR[ 246 ][ 349 ],
   alphaCSR[ 246 ][ 350 ],
   alphaCSR[ 246 ][ 351 ],
   alphaCSR[ 246 ][ 352 ],
   alphaCSR[ 246 ][ 353 ],
   alphaCSR[ 246 ][ 354 ],
   alphaCSR[ 246 ][ 355 ],
   alphaCSR[ 246 ][ 356 ],
   alphaCSR[ 246 ][ 357 ],
   alphaCSR[ 246 ][ 358 ],
   alphaCSR[ 246 ][ 359 ],
   alphaCSR[ 246 ][ 360 ],
   alphaCSR[ 246 ][ 361 ],
   alphaCSR[ 246 ][ 362 ],
   alphaCSR[ 246 ][ 363 ],
   alphaCSR[ 246 ][ 364 ],
   alphaCSR[ 246 ][ 365 ],
   alphaCSR[ 246 ][ 366 ],
   alphaCSR[ 246 ][ 367 ],
   alphaCSR[ 246 ][ 368 ],
   alphaCSR[ 246 ][ 369 ],
   alphaCSR[ 246 ][ 370 ],
   alphaCSR[ 246 ][ 371 ],
   alphaCSR[ 246 ][ 372 ],
   alphaCSR[ 246 ][ 373 ],
   alphaCSR[ 246 ][ 374 ],
   alphaCSR[ 246 ][ 375 ],
   alphaCSR[ 246 ][ 376 ],
   alphaCSR[ 246 ][ 377 ],
   alphaCSR[ 246 ][ 378 ],
   alphaCSR[ 246 ][ 379 ],
   alphaCSR[ 246 ][ 380 ],
   alphaCSR[ 246 ][ 381 ],
   alphaCSR[ 246 ][ 382 ],
   alphaCSR[ 246 ][ 383 ],
   alphaCSR[ 247 ][ 0 ],
   alphaCSR[ 247 ][ 1 ],
   alphaCSR[ 247 ][ 2 ],
   alphaCSR[ 247 ][ 3 ],
   alphaCSR[ 247 ][ 4 ],
   alphaCSR[ 247 ][ 5 ],
   alphaCSR[ 247 ][ 6 ],
   alphaCSR[ 247 ][ 7 ],
   alphaCSR[ 247 ][ 8 ],
   alphaCSR[ 247 ][ 9 ],
   alphaCSR[ 247 ][ 10 ],
   alphaCSR[ 247 ][ 11 ],
   alphaCSR[ 247 ][ 12 ],
   alphaCSR[ 247 ][ 13 ],
   alphaCSR[ 247 ][ 14 ],
   alphaCSR[ 247 ][ 15 ],
   alphaCSR[ 247 ][ 16 ],
   alphaCSR[ 247 ][ 17 ],
   alphaCSR[ 247 ][ 18 ],
   alphaCSR[ 247 ][ 19 ],
   alphaCSR[ 247 ][ 20 ],
   alphaCSR[ 247 ][ 21 ],
   alphaCSR[ 247 ][ 22 ],
   alphaCSR[ 247 ][ 23 ],
   alphaCSR[ 247 ][ 24 ],
   alphaCSR[ 247 ][ 25 ],
   alphaCSR[ 247 ][ 26 ],
   alphaCSR[ 247 ][ 27 ],
   alphaCSR[ 247 ][ 28 ],
   alphaCSR[ 247 ][ 29 ],
   alphaCSR[ 247 ][ 30 ],
   alphaCSR[ 247 ][ 31 ],
   alphaCSR[ 247 ][ 32 ],
   alphaCSR[ 247 ][ 33 ],
   alphaCSR[ 247 ][ 34 ],
   alphaCSR[ 247 ][ 35 ],
   alphaCSR[ 247 ][ 36 ],
   alphaCSR[ 247 ][ 37 ],
   alphaCSR[ 247 ][ 38 ],
   alphaCSR[ 247 ][ 39 ],
   alphaCSR[ 247 ][ 40 ],
   alphaCSR[ 247 ][ 41 ],
   alphaCSR[ 247 ][ 42 ],
   alphaCSR[ 247 ][ 43 ],
   alphaCSR[ 247 ][ 44 ],
   alphaCSR[ 247 ][ 45 ],
   alphaCSR[ 247 ][ 46 ],
   alphaCSR[ 247 ][ 47 ],
   alphaCSR[ 247 ][ 48 ],
   alphaCSR[ 247 ][ 49 ],
   alphaCSR[ 247 ][ 50 ],
   alphaCSR[ 247 ][ 51 ],
   alphaCSR[ 247 ][ 52 ],
   alphaCSR[ 247 ][ 53 ],
   alphaCSR[ 247 ][ 54 ],
   alphaCSR[ 247 ][ 55 ],
   alphaCSR[ 247 ][ 56 ],
   alphaCSR[ 247 ][ 57 ],
   alphaCSR[ 247 ][ 58 ],
   alphaCSR[ 247 ][ 59 ],
   alphaCSR[ 247 ][ 60 ],
   alphaCSR[ 247 ][ 61 ],
   alphaCSR[ 247 ][ 62 ],
   alphaCSR[ 247 ][ 63 ],
   alphaCSR[ 247 ][ 64 ],
   alphaCSR[ 247 ][ 65 ],
   alphaCSR[ 247 ][ 66 ],
   alphaCSR[ 247 ][ 67 ],
   alphaCSR[ 247 ][ 68 ],
   alphaCSR[ 247 ][ 69 ],
   alphaCSR[ 247 ][ 70 ],
   alphaCSR[ 247 ][ 71 ],
   alphaCSR[ 247 ][ 72 ],
   alphaCSR[ 247 ][ 73 ],
   alphaCSR[ 247 ][ 74 ],
   alphaCSR[ 247 ][ 75 ],
   alphaCSR[ 247 ][ 76 ],
   alphaCSR[ 247 ][ 77 ],
   alphaCSR[ 247 ][ 78 ],
   alphaCSR[ 247 ][ 79 ],
   alphaCSR[ 247 ][ 80 ],
   alphaCSR[ 247 ][ 81 ],
   alphaCSR[ 247 ][ 82 ],
   alphaCSR[ 247 ][ 83 ],
   alphaCSR[ 247 ][ 84 ],
   alphaCSR[ 247 ][ 85 ],
   alphaCSR[ 247 ][ 86 ],
   alphaCSR[ 247 ][ 87 ],
   alphaCSR[ 247 ][ 88 ],
   alphaCSR[ 247 ][ 89 ],
   alphaCSR[ 247 ][ 90 ],
   alphaCSR[ 247 ][ 91 ],
   alphaCSR[ 247 ][ 92 ],
   alphaCSR[ 247 ][ 93 ],
   alphaCSR[ 247 ][ 94 ],
   alphaCSR[ 247 ][ 95 ],
   alphaCSR[ 247 ][ 96 ],
   alphaCSR[ 247 ][ 97 ],
   alphaCSR[ 247 ][ 98 ],
   alphaCSR[ 247 ][ 99 ],
   alphaCSR[ 247 ][ 100 ],
   alphaCSR[ 247 ][ 101 ],
   alphaCSR[ 247 ][ 102 ],
   alphaCSR[ 247 ][ 103 ],
   alphaCSR[ 247 ][ 104 ],
   alphaCSR[ 247 ][ 105 ],
   alphaCSR[ 247 ][ 106 ],
   alphaCSR[ 247 ][ 107 ],
   alphaCSR[ 247 ][ 108 ],
   alphaCSR[ 247 ][ 109 ],
   alphaCSR[ 247 ][ 110 ],
   alphaCSR[ 247 ][ 111 ],
   alphaCSR[ 247 ][ 112 ],
   alphaCSR[ 247 ][ 113 ],
   alphaCSR[ 247 ][ 114 ],
   alphaCSR[ 247 ][ 115 ],
   alphaCSR[ 247 ][ 116 ],
   alphaCSR[ 247 ][ 117 ],
   alphaCSR[ 247 ][ 118 ],
   alphaCSR[ 247 ][ 119 ],
   alphaCSR[ 247 ][ 120 ],
   alphaCSR[ 247 ][ 121 ],
   alphaCSR[ 247 ][ 122 ],
   alphaCSR[ 247 ][ 123 ],
   alphaCSR[ 247 ][ 124 ],
   alphaCSR[ 247 ][ 125 ],
   alphaCSR[ 247 ][ 126 ],
   alphaCSR[ 247 ][ 127 ],
   alphaCSR[ 247 ][ 128 ],
   alphaCSR[ 247 ][ 129 ],
   alphaCSR[ 247 ][ 130 ],
   alphaCSR[ 247 ][ 131 ],
   alphaCSR[ 247 ][ 132 ],
   alphaCSR[ 247 ][ 133 ],
   alphaCSR[ 247 ][ 134 ],
   alphaCSR[ 247 ][ 135 ],
   alphaCSR[ 247 ][ 136 ],
   alphaCSR[ 247 ][ 137 ],
   alphaCSR[ 247 ][ 138 ],
   alphaCSR[ 247 ][ 139 ],
   alphaCSR[ 247 ][ 140 ],
   alphaCSR[ 247 ][ 141 ],
   alphaCSR[ 247 ][ 142 ],
   alphaCSR[ 247 ][ 143 ],
   alphaCSR[ 247 ][ 144 ],
   alphaCSR[ 247 ][ 145 ],
   alphaCSR[ 247 ][ 146 ],
   alphaCSR[ 247 ][ 147 ],
   alphaCSR[ 247 ][ 148 ],
   alphaCSR[ 247 ][ 149 ],
   alphaCSR[ 247 ][ 150 ],
   alphaCSR[ 247 ][ 151 ],
   alphaCSR[ 247 ][ 152 ],
   alphaCSR[ 247 ][ 153 ],
   alphaCSR[ 247 ][ 154 ],
   alphaCSR[ 247 ][ 155 ],
   alphaCSR[ 247 ][ 156 ],
   alphaCSR[ 247 ][ 157 ],
   alphaCSR[ 247 ][ 158 ],
   alphaCSR[ 247 ][ 159 ],
   alphaCSR[ 247 ][ 160 ],
   alphaCSR[ 247 ][ 161 ],
   alphaCSR[ 247 ][ 162 ],
   alphaCSR[ 247 ][ 163 ],
   alphaCSR[ 247 ][ 164 ],
   alphaCSR[ 247 ][ 165 ],
   alphaCSR[ 247 ][ 166 ],
   alphaCSR[ 247 ][ 167 ],
   alphaCSR[ 247 ][ 168 ],
   alphaCSR[ 247 ][ 169 ],
   alphaCSR[ 247 ][ 170 ],
   alphaCSR[ 247 ][ 171 ],
   alphaCSR[ 247 ][ 172 ],
   alphaCSR[ 247 ][ 173 ],
   alphaCSR[ 247 ][ 174 ],
   alphaCSR[ 247 ][ 175 ],
   alphaCSR[ 247 ][ 176 ],
   alphaCSR[ 247 ][ 177 ],
   alphaCSR[ 247 ][ 178 ],
   alphaCSR[ 247 ][ 179 ],
   alphaCSR[ 247 ][ 180 ],
   alphaCSR[ 247 ][ 181 ],
   alphaCSR[ 247 ][ 182 ],
   alphaCSR[ 247 ][ 183 ],
   alphaCSR[ 247 ][ 184 ],
   alphaCSR[ 247 ][ 185 ],
   alphaCSR[ 247 ][ 186 ],
   alphaCSR[ 247 ][ 187 ],
   alphaCSR[ 247 ][ 188 ],
   alphaCSR[ 247 ][ 189 ],
   alphaCSR[ 247 ][ 190 ],
   alphaCSR[ 247 ][ 191 ],
   alphaCSR[ 247 ][ 192 ],
   alphaCSR[ 247 ][ 193 ],
   alphaCSR[ 247 ][ 194 ],
   alphaCSR[ 247 ][ 195 ],
   alphaCSR[ 247 ][ 196 ],
   alphaCSR[ 247 ][ 197 ],
   alphaCSR[ 247 ][ 198 ],
   alphaCSR[ 247 ][ 199 ],
   alphaCSR[ 247 ][ 200 ],
   alphaCSR[ 247 ][ 201 ],
   alphaCSR[ 247 ][ 202 ],
   alphaCSR[ 247 ][ 203 ],
   alphaCSR[ 247 ][ 204 ],
   alphaCSR[ 247 ][ 205 ],
   alphaCSR[ 247 ][ 206 ],
   alphaCSR[ 247 ][ 207 ],
   alphaCSR[ 247 ][ 208 ],
   alphaCSR[ 247 ][ 209 ],
   alphaCSR[ 247 ][ 210 ],
   alphaCSR[ 247 ][ 211 ],
   alphaCSR[ 247 ][ 212 ],
   alphaCSR[ 247 ][ 213 ],
   alphaCSR[ 247 ][ 214 ],
   alphaCSR[ 247 ][ 215 ],
   alphaCSR[ 247 ][ 216 ],
   alphaCSR[ 247 ][ 217 ],
   alphaCSR[ 247 ][ 218 ],
   alphaCSR[ 247 ][ 219 ],
   alphaCSR[ 247 ][ 220 ],
   alphaCSR[ 247 ][ 221 ],
   alphaCSR[ 247 ][ 222 ],
   alphaCSR[ 247 ][ 223 ],
   alphaCSR[ 247 ][ 224 ],
   alphaCSR[ 247 ][ 225 ],
   alphaCSR[ 247 ][ 226 ],
   alphaCSR[ 247 ][ 227 ],
   alphaCSR[ 247 ][ 228 ],
   alphaCSR[ 247 ][ 229 ],
   alphaCSR[ 247 ][ 230 ],
   alphaCSR[ 247 ][ 231 ],
   alphaCSR[ 247 ][ 232 ],
   alphaCSR[ 247 ][ 233 ],
   alphaCSR[ 247 ][ 234 ],
   alphaCSR[ 247 ][ 235 ],
   alphaCSR[ 247 ][ 236 ],
   alphaCSR[ 247 ][ 237 ],
   alphaCSR[ 247 ][ 238 ],
   alphaCSR[ 247 ][ 239 ],
   alphaCSR[ 247 ][ 240 ],
   alphaCSR[ 247 ][ 241 ],
   alphaCSR[ 247 ][ 242 ],
   alphaCSR[ 247 ][ 243 ],
   alphaCSR[ 247 ][ 244 ],
   alphaCSR[ 247 ][ 245 ],
   alphaCSR[ 247 ][ 246 ],
   alphaCSR[ 247 ][ 247 ],
   alphaCSR[ 247 ][ 248 ],
   alphaCSR[ 247 ][ 249 ],
   alphaCSR[ 247 ][ 250 ],
   alphaCSR[ 247 ][ 251 ],
   alphaCSR[ 247 ][ 252 ],
   alphaCSR[ 247 ][ 253 ],
   alphaCSR[ 247 ][ 254 ],
   alphaCSR[ 247 ][ 255 ],
   alphaCSR[ 247 ][ 256 ],
   alphaCSR[ 247 ][ 257 ],
   alphaCSR[ 247 ][ 258 ],
   alphaCSR[ 247 ][ 259 ],
   alphaCSR[ 247 ][ 260 ],
   alphaCSR[ 247 ][ 261 ],
   alphaCSR[ 247 ][ 262 ],
   alphaCSR[ 247 ][ 263 ],
   alphaCSR[ 247 ][ 264 ],
   alphaCSR[ 247 ][ 265 ],
   alphaCSR[ 247 ][ 266 ],
   alphaCSR[ 247 ][ 267 ],
   alphaCSR[ 247 ][ 268 ],
   alphaCSR[ 247 ][ 269 ],
   alphaCSR[ 247 ][ 270 ],
   alphaCSR[ 247 ][ 271 ],
   alphaCSR[ 247 ][ 272 ],
   alphaCSR[ 247 ][ 273 ],
   alphaCSR[ 247 ][ 274 ],
   alphaCSR[ 247 ][ 275 ],
   alphaCSR[ 247 ][ 276 ],
   alphaCSR[ 247 ][ 277 ],
   alphaCSR[ 247 ][ 278 ],
   alphaCSR[ 247 ][ 279 ],
   alphaCSR[ 247 ][ 280 ],
   alphaCSR[ 247 ][ 281 ],
   alphaCSR[ 247 ][ 282 ],
   alphaCSR[ 247 ][ 283 ],
   alphaCSR[ 247 ][ 284 ],
   alphaCSR[ 247 ][ 285 ],
   alphaCSR[ 247 ][ 286 ],
   alphaCSR[ 247 ][ 287 ],
   alphaCSR[ 247 ][ 288 ],
   alphaCSR[ 247 ][ 289 ],
   alphaCSR[ 247 ][ 290 ],
   alphaCSR[ 247 ][ 291 ],
   alphaCSR[ 247 ][ 292 ],
   alphaCSR[ 247 ][ 293 ],
   alphaCSR[ 247 ][ 294 ],
   alphaCSR[ 247 ][ 295 ],
   alphaCSR[ 247 ][ 296 ],
   alphaCSR[ 247 ][ 297 ],
   alphaCSR[ 247 ][ 298 ],
   alphaCSR[ 247 ][ 299 ],
   alphaCSR[ 247 ][ 300 ],
   alphaCSR[ 247 ][ 301 ],
   alphaCSR[ 247 ][ 302 ],
   alphaCSR[ 247 ][ 303 ],
   alphaCSR[ 247 ][ 304 ],
   alphaCSR[ 247 ][ 305 ],
   alphaCSR[ 247 ][ 306 ],
   alphaCSR[ 247 ][ 307 ],
   alphaCSR[ 247 ][ 308 ],
   alphaCSR[ 247 ][ 309 ],
   alphaCSR[ 247 ][ 310 ],
   alphaCSR[ 247 ][ 311 ],
   alphaCSR[ 247 ][ 312 ],
   alphaCSR[ 247 ][ 313 ],
   alphaCSR[ 247 ][ 314 ],
   alphaCSR[ 247 ][ 315 ],
   alphaCSR[ 247 ][ 316 ],
   alphaCSR[ 247 ][ 317 ],
   alphaCSR[ 247 ][ 318 ],
   alphaCSR[ 247 ][ 319 ],
   alphaCSR[ 247 ][ 320 ],
   alphaCSR[ 247 ][ 321 ],
   alphaCSR[ 247 ][ 322 ],
   alphaCSR[ 247 ][ 323 ],
   alphaCSR[ 247 ][ 324 ],
   alphaCSR[ 247 ][ 325 ],
   alphaCSR[ 247 ][ 326 ],
   alphaCSR[ 247 ][ 327 ],
   alphaCSR[ 247 ][ 328 ],
   alphaCSR[ 247 ][ 329 ],
   alphaCSR[ 247 ][ 330 ],
   alphaCSR[ 247 ][ 331 ],
   alphaCSR[ 247 ][ 332 ],
   alphaCSR[ 247 ][ 333 ],
   alphaCSR[ 247 ][ 334 ],
   alphaCSR[ 247 ][ 335 ],
   alphaCSR[ 247 ][ 336 ],
   alphaCSR[ 247 ][ 337 ],
   alphaCSR[ 247 ][ 338 ],
   alphaCSR[ 247 ][ 339 ],
   alphaCSR[ 247 ][ 340 ],
   alphaCSR[ 247 ][ 341 ],
   alphaCSR[ 247 ][ 342 ],
   alphaCSR[ 247 ][ 343 ],
   alphaCSR[ 247 ][ 344 ],
   alphaCSR[ 247 ][ 345 ],
   alphaCSR[ 247 ][ 346 ],
   alphaCSR[ 247 ][ 347 ],
   alphaCSR[ 247 ][ 348 ],
   alphaCSR[ 247 ][ 349 ],
   alphaCSR[ 247 ][ 350 ],
   alphaCSR[ 247 ][ 351 ],
   alphaCSR[ 247 ][ 352 ],
   alphaCSR[ 247 ][ 353 ],
   alphaCSR[ 247 ][ 354 ],
   alphaCSR[ 247 ][ 355 ],
   alphaCSR[ 247 ][ 356 ],
   alphaCSR[ 247 ][ 357 ],
   alphaCSR[ 247 ][ 358 ],
   alphaCSR[ 247 ][ 359 ],
   alphaCSR[ 247 ][ 360 ],
   alphaCSR[ 247 ][ 361 ],
   alphaCSR[ 247 ][ 362 ],
   alphaCSR[ 247 ][ 363 ],
   alphaCSR[ 247 ][ 364 ],
   alphaCSR[ 247 ][ 365 ],
   alphaCSR[ 247 ][ 366 ],
   alphaCSR[ 247 ][ 367 ],
   alphaCSR[ 247 ][ 368 ],
   alphaCSR[ 247 ][ 369 ],
   alphaCSR[ 247 ][ 370 ],
   alphaCSR[ 247 ][ 371 ],
   alphaCSR[ 247 ][ 372 ],
   alphaCSR[ 247 ][ 373 ],
   alphaCSR[ 247 ][ 374 ],
   alphaCSR[ 247 ][ 375 ],
   alphaCSR[ 247 ][ 376 ],
   alphaCSR[ 247 ][ 377 ],
   alphaCSR[ 247 ][ 378 ],
   alphaCSR[ 247 ][ 379 ],
   alphaCSR[ 247 ][ 380 ],
   alphaCSR[ 247 ][ 381 ],
   alphaCSR[ 247 ][ 382 ],
   alphaCSR[ 247 ][ 383 ],
   alphaCSR[ 248 ][ 0 ],
   alphaCSR[ 248 ][ 1 ],
   alphaCSR[ 248 ][ 2 ],
   alphaCSR[ 248 ][ 3 ],
   alphaCSR[ 248 ][ 4 ],
   alphaCSR[ 248 ][ 5 ],
   alphaCSR[ 248 ][ 6 ],
   alphaCSR[ 248 ][ 7 ],
   alphaCSR[ 248 ][ 8 ],
   alphaCSR[ 248 ][ 9 ],
   alphaCSR[ 248 ][ 10 ],
   alphaCSR[ 248 ][ 11 ],
   alphaCSR[ 248 ][ 12 ],
   alphaCSR[ 248 ][ 13 ],
   alphaCSR[ 248 ][ 14 ],
   alphaCSR[ 248 ][ 15 ],
   alphaCSR[ 248 ][ 16 ],
   alphaCSR[ 248 ][ 17 ],
   alphaCSR[ 248 ][ 18 ],
   alphaCSR[ 248 ][ 19 ],
   alphaCSR[ 248 ][ 20 ],
   alphaCSR[ 248 ][ 21 ],
   alphaCSR[ 248 ][ 22 ],
   alphaCSR[ 248 ][ 23 ],
   alphaCSR[ 248 ][ 24 ],
   alphaCSR[ 248 ][ 25 ],
   alphaCSR[ 248 ][ 26 ],
   alphaCSR[ 248 ][ 27 ],
   alphaCSR[ 248 ][ 28 ],
   alphaCSR[ 248 ][ 29 ],
   alphaCSR[ 248 ][ 30 ],
   alphaCSR[ 248 ][ 31 ],
   alphaCSR[ 248 ][ 32 ],
   alphaCSR[ 248 ][ 33 ],
   alphaCSR[ 248 ][ 34 ],
   alphaCSR[ 248 ][ 35 ],
   alphaCSR[ 248 ][ 36 ],
   alphaCSR[ 248 ][ 37 ],
   alphaCSR[ 248 ][ 38 ],
   alphaCSR[ 248 ][ 39 ],
   alphaCSR[ 248 ][ 40 ],
   alphaCSR[ 248 ][ 41 ],
   alphaCSR[ 248 ][ 42 ],
   alphaCSR[ 248 ][ 43 ],
   alphaCSR[ 248 ][ 44 ],
   alphaCSR[ 248 ][ 45 ],
   alphaCSR[ 248 ][ 46 ],
   alphaCSR[ 248 ][ 47 ],
   alphaCSR[ 248 ][ 48 ],
   alphaCSR[ 248 ][ 49 ],
   alphaCSR[ 248 ][ 50 ],
   alphaCSR[ 248 ][ 51 ],
   alphaCSR[ 248 ][ 52 ],
   alphaCSR[ 248 ][ 53 ],
   alphaCSR[ 248 ][ 54 ],
   alphaCSR[ 248 ][ 55 ],
   alphaCSR[ 248 ][ 56 ],
   alphaCSR[ 248 ][ 57 ],
   alphaCSR[ 248 ][ 58 ],
   alphaCSR[ 248 ][ 59 ],
   alphaCSR[ 248 ][ 60 ],
   alphaCSR[ 248 ][ 61 ],
   alphaCSR[ 248 ][ 62 ],
   alphaCSR[ 248 ][ 63 ],
   alphaCSR[ 248 ][ 64 ],
   alphaCSR[ 248 ][ 65 ],
   alphaCSR[ 248 ][ 66 ],
   alphaCSR[ 248 ][ 67 ],
   alphaCSR[ 248 ][ 68 ],
   alphaCSR[ 248 ][ 69 ],
   alphaCSR[ 248 ][ 70 ],
   alphaCSR[ 248 ][ 71 ],
   alphaCSR[ 248 ][ 72 ],
   alphaCSR[ 248 ][ 73 ],
   alphaCSR[ 248 ][ 74 ],
   alphaCSR[ 248 ][ 75 ],
   alphaCSR[ 248 ][ 76 ],
   alphaCSR[ 248 ][ 77 ],
   alphaCSR[ 248 ][ 78 ],
   alphaCSR[ 248 ][ 79 ],
   alphaCSR[ 248 ][ 80 ],
   alphaCSR[ 248 ][ 81 ],
   alphaCSR[ 248 ][ 82 ],
   alphaCSR[ 248 ][ 83 ],
   alphaCSR[ 248 ][ 84 ],
   alphaCSR[ 248 ][ 85 ],
   alphaCSR[ 248 ][ 86 ],
   alphaCSR[ 248 ][ 87 ],
   alphaCSR[ 248 ][ 88 ],
   alphaCSR[ 248 ][ 89 ],
   alphaCSR[ 248 ][ 90 ],
   alphaCSR[ 248 ][ 91 ],
   alphaCSR[ 248 ][ 92 ],
   alphaCSR[ 248 ][ 93 ],
   alphaCSR[ 248 ][ 94 ],
   alphaCSR[ 248 ][ 95 ],
   alphaCSR[ 248 ][ 96 ],
   alphaCSR[ 248 ][ 97 ],
   alphaCSR[ 248 ][ 98 ],
   alphaCSR[ 248 ][ 99 ],
   alphaCSR[ 248 ][ 100 ],
   alphaCSR[ 248 ][ 101 ],
   alphaCSR[ 248 ][ 102 ],
   alphaCSR[ 248 ][ 103 ],
   alphaCSR[ 248 ][ 104 ],
   alphaCSR[ 248 ][ 105 ],
   alphaCSR[ 248 ][ 106 ],
   alphaCSR[ 248 ][ 107 ],
   alphaCSR[ 248 ][ 108 ],
   alphaCSR[ 248 ][ 109 ],
   alphaCSR[ 248 ][ 110 ],
   alphaCSR[ 248 ][ 111 ],
   alphaCSR[ 248 ][ 112 ],
   alphaCSR[ 248 ][ 113 ],
   alphaCSR[ 248 ][ 114 ],
   alphaCSR[ 248 ][ 115 ],
   alphaCSR[ 248 ][ 116 ],
   alphaCSR[ 248 ][ 117 ],
   alphaCSR[ 248 ][ 118 ],
   alphaCSR[ 248 ][ 119 ],
   alphaCSR[ 248 ][ 120 ],
   alphaCSR[ 248 ][ 121 ],
   alphaCSR[ 248 ][ 122 ],
   alphaCSR[ 248 ][ 123 ],
   alphaCSR[ 248 ][ 124 ],
   alphaCSR[ 248 ][ 125 ],
   alphaCSR[ 248 ][ 126 ],
   alphaCSR[ 248 ][ 127 ],
   alphaCSR[ 248 ][ 128 ],
   alphaCSR[ 248 ][ 129 ],
   alphaCSR[ 248 ][ 130 ],
   alphaCSR[ 248 ][ 131 ],
   alphaCSR[ 248 ][ 132 ],
   alphaCSR[ 248 ][ 133 ],
   alphaCSR[ 248 ][ 134 ],
   alphaCSR[ 248 ][ 135 ],
   alphaCSR[ 248 ][ 136 ],
   alphaCSR[ 248 ][ 137 ],
   alphaCSR[ 248 ][ 138 ],
   alphaCSR[ 248 ][ 139 ],
   alphaCSR[ 248 ][ 140 ],
   alphaCSR[ 248 ][ 141 ],
   alphaCSR[ 248 ][ 142 ],
   alphaCSR[ 248 ][ 143 ],
   alphaCSR[ 248 ][ 144 ],
   alphaCSR[ 248 ][ 145 ],
   alphaCSR[ 248 ][ 146 ],
   alphaCSR[ 248 ][ 147 ],
   alphaCSR[ 248 ][ 148 ],
   alphaCSR[ 248 ][ 149 ],
   alphaCSR[ 248 ][ 150 ],
   alphaCSR[ 248 ][ 151 ],
   alphaCSR[ 248 ][ 152 ],
   alphaCSR[ 248 ][ 153 ],
   alphaCSR[ 248 ][ 154 ],
   alphaCSR[ 248 ][ 155 ],
   alphaCSR[ 248 ][ 156 ],
   alphaCSR[ 248 ][ 157 ],
   alphaCSR[ 248 ][ 158 ],
   alphaCSR[ 248 ][ 159 ],
   alphaCSR[ 248 ][ 160 ],
   alphaCSR[ 248 ][ 161 ],
   alphaCSR[ 248 ][ 162 ],
   alphaCSR[ 248 ][ 163 ],
   alphaCSR[ 248 ][ 164 ],
   alphaCSR[ 248 ][ 165 ],
   alphaCSR[ 248 ][ 166 ],
   alphaCSR[ 248 ][ 167 ],
   alphaCSR[ 248 ][ 168 ],
   alphaCSR[ 248 ][ 169 ],
   alphaCSR[ 248 ][ 170 ],
   alphaCSR[ 248 ][ 171 ],
   alphaCSR[ 248 ][ 172 ],
   alphaCSR[ 248 ][ 173 ],
   alphaCSR[ 248 ][ 174 ],
   alphaCSR[ 248 ][ 175 ],
   alphaCSR[ 248 ][ 176 ],
   alphaCSR[ 248 ][ 177 ],
   alphaCSR[ 248 ][ 178 ],
   alphaCSR[ 248 ][ 179 ],
   alphaCSR[ 248 ][ 180 ],
   alphaCSR[ 248 ][ 181 ],
   alphaCSR[ 248 ][ 182 ],
   alphaCSR[ 248 ][ 183 ],
   alphaCSR[ 248 ][ 184 ],
   alphaCSR[ 248 ][ 185 ],
   alphaCSR[ 248 ][ 186 ],
   alphaCSR[ 248 ][ 187 ],
   alphaCSR[ 248 ][ 188 ],
   alphaCSR[ 248 ][ 189 ],
   alphaCSR[ 248 ][ 190 ],
   alphaCSR[ 248 ][ 191 ],
   alphaCSR[ 248 ][ 192 ],
   alphaCSR[ 248 ][ 193 ],
   alphaCSR[ 248 ][ 194 ],
   alphaCSR[ 248 ][ 195 ],
   alphaCSR[ 248 ][ 196 ],
   alphaCSR[ 248 ][ 197 ],
   alphaCSR[ 248 ][ 198 ],
   alphaCSR[ 248 ][ 199 ],
   alphaCSR[ 248 ][ 200 ],
   alphaCSR[ 248 ][ 201 ],
   alphaCSR[ 248 ][ 202 ],
   alphaCSR[ 248 ][ 203 ],
   alphaCSR[ 248 ][ 204 ],
   alphaCSR[ 248 ][ 205 ],
   alphaCSR[ 248 ][ 206 ],
   alphaCSR[ 248 ][ 207 ],
   alphaCSR[ 248 ][ 208 ],
   alphaCSR[ 248 ][ 209 ],
   alphaCSR[ 248 ][ 210 ],
   alphaCSR[ 248 ][ 211 ],
   alphaCSR[ 248 ][ 212 ],
   alphaCSR[ 248 ][ 213 ],
   alphaCSR[ 248 ][ 214 ],
   alphaCSR[ 248 ][ 215 ],
   alphaCSR[ 248 ][ 216 ],
   alphaCSR[ 248 ][ 217 ],
   alphaCSR[ 248 ][ 218 ],
   alphaCSR[ 248 ][ 219 ],
   alphaCSR[ 248 ][ 220 ],
   alphaCSR[ 248 ][ 221 ],
   alphaCSR[ 248 ][ 222 ],
   alphaCSR[ 248 ][ 223 ],
   alphaCSR[ 248 ][ 224 ],
   alphaCSR[ 248 ][ 225 ],
   alphaCSR[ 248 ][ 226 ],
   alphaCSR[ 248 ][ 227 ],
   alphaCSR[ 248 ][ 228 ],
   alphaCSR[ 248 ][ 229 ],
   alphaCSR[ 248 ][ 230 ],
   alphaCSR[ 248 ][ 231 ],
   alphaCSR[ 248 ][ 232 ],
   alphaCSR[ 248 ][ 233 ],
   alphaCSR[ 248 ][ 234 ],
   alphaCSR[ 248 ][ 235 ],
   alphaCSR[ 248 ][ 236 ],
   alphaCSR[ 248 ][ 237 ],
   alphaCSR[ 248 ][ 238 ],
   alphaCSR[ 248 ][ 239 ],
   alphaCSR[ 248 ][ 240 ],
   alphaCSR[ 248 ][ 241 ],
   alphaCSR[ 248 ][ 242 ],
   alphaCSR[ 248 ][ 243 ],
   alphaCSR[ 248 ][ 244 ],
   alphaCSR[ 248 ][ 245 ],
   alphaCSR[ 248 ][ 246 ],
   alphaCSR[ 248 ][ 247 ],
   alphaCSR[ 248 ][ 248 ],
   alphaCSR[ 248 ][ 249 ],
   alphaCSR[ 248 ][ 250 ],
   alphaCSR[ 248 ][ 251 ],
   alphaCSR[ 248 ][ 252 ],
   alphaCSR[ 248 ][ 253 ],
   alphaCSR[ 248 ][ 254 ],
   alphaCSR[ 248 ][ 255 ],
   alphaCSR[ 248 ][ 256 ],
   alphaCSR[ 248 ][ 257 ],
   alphaCSR[ 248 ][ 258 ],
   alphaCSR[ 248 ][ 259 ],
   alphaCSR[ 248 ][ 260 ],
   alphaCSR[ 248 ][ 261 ],
   alphaCSR[ 248 ][ 262 ],
   alphaCSR[ 248 ][ 263 ],
   alphaCSR[ 248 ][ 264 ],
   alphaCSR[ 248 ][ 265 ],
   alphaCSR[ 248 ][ 266 ],
   alphaCSR[ 248 ][ 267 ],
   alphaCSR[ 248 ][ 268 ],
   alphaCSR[ 248 ][ 269 ],
   alphaCSR[ 248 ][ 270 ],
   alphaCSR[ 248 ][ 271 ],
   alphaCSR[ 248 ][ 272 ],
   alphaCSR[ 248 ][ 273 ],
   alphaCSR[ 248 ][ 274 ],
   alphaCSR[ 248 ][ 275 ],
   alphaCSR[ 248 ][ 276 ],
   alphaCSR[ 248 ][ 277 ],
   alphaCSR[ 248 ][ 278 ],
   alphaCSR[ 248 ][ 279 ],
   alphaCSR[ 248 ][ 280 ],
   alphaCSR[ 248 ][ 281 ],
   alphaCSR[ 248 ][ 282 ],
   alphaCSR[ 248 ][ 283 ],
   alphaCSR[ 248 ][ 284 ],
   alphaCSR[ 248 ][ 285 ],
   alphaCSR[ 248 ][ 286 ],
   alphaCSR[ 248 ][ 287 ],
   alphaCSR[ 248 ][ 288 ],
   alphaCSR[ 248 ][ 289 ],
   alphaCSR[ 248 ][ 290 ],
   alphaCSR[ 248 ][ 291 ],
   alphaCSR[ 248 ][ 292 ],
   alphaCSR[ 248 ][ 293 ],
   alphaCSR[ 248 ][ 294 ],
   alphaCSR[ 248 ][ 295 ],
   alphaCSR[ 248 ][ 296 ],
   alphaCSR[ 248 ][ 297 ],
   alphaCSR[ 248 ][ 298 ],
   alphaCSR[ 248 ][ 299 ],
   alphaCSR[ 248 ][ 300 ],
   alphaCSR[ 248 ][ 301 ],
   alphaCSR[ 248 ][ 302 ],
   alphaCSR[ 248 ][ 303 ],
   alphaCSR[ 248 ][ 304 ],
   alphaCSR[ 248 ][ 305 ],
   alphaCSR[ 248 ][ 306 ],
   alphaCSR[ 248 ][ 307 ],
   alphaCSR[ 248 ][ 308 ],
   alphaCSR[ 248 ][ 309 ],
   alphaCSR[ 248 ][ 310 ],
   alphaCSR[ 248 ][ 311 ],
   alphaCSR[ 248 ][ 312 ],
   alphaCSR[ 248 ][ 313 ],
   alphaCSR[ 248 ][ 314 ],
   alphaCSR[ 248 ][ 315 ],
   alphaCSR[ 248 ][ 316 ],
   alphaCSR[ 248 ][ 317 ],
   alphaCSR[ 248 ][ 318 ],
   alphaCSR[ 248 ][ 319 ],
   alphaCSR[ 248 ][ 320 ],
   alphaCSR[ 248 ][ 321 ],
   alphaCSR[ 248 ][ 322 ],
   alphaCSR[ 248 ][ 323 ],
   alphaCSR[ 248 ][ 324 ],
   alphaCSR[ 248 ][ 325 ],
   alphaCSR[ 248 ][ 326 ],
   alphaCSR[ 248 ][ 327 ],
   alphaCSR[ 248 ][ 328 ],
   alphaCSR[ 248 ][ 329 ],
   alphaCSR[ 248 ][ 330 ],
   alphaCSR[ 248 ][ 331 ],
   alphaCSR[ 248 ][ 332 ],
   alphaCSR[ 248 ][ 333 ],
   alphaCSR[ 248 ][ 334 ],
   alphaCSR[ 248 ][ 335 ],
   alphaCSR[ 248 ][ 336 ],
   alphaCSR[ 248 ][ 337 ],
   alphaCSR[ 248 ][ 338 ],
   alphaCSR[ 248 ][ 339 ],
   alphaCSR[ 248 ][ 340 ],
   alphaCSR[ 248 ][ 341 ],
   alphaCSR[ 248 ][ 342 ],
   alphaCSR[ 248 ][ 343 ],
   alphaCSR[ 248 ][ 344 ],
   alphaCSR[ 248 ][ 345 ],
   alphaCSR[ 248 ][ 346 ],
   alphaCSR[ 248 ][ 347 ],
   alphaCSR[ 248 ][ 348 ],
   alphaCSR[ 248 ][ 349 ],
   alphaCSR[ 248 ][ 350 ],
   alphaCSR[ 248 ][ 351 ],
   alphaCSR[ 248 ][ 352 ],
   alphaCSR[ 248 ][ 353 ],
   alphaCSR[ 248 ][ 354 ],
   alphaCSR[ 248 ][ 355 ],
   alphaCSR[ 248 ][ 356 ],
   alphaCSR[ 248 ][ 357 ],
   alphaCSR[ 248 ][ 358 ],
   alphaCSR[ 248 ][ 359 ],
   alphaCSR[ 248 ][ 360 ],
   alphaCSR[ 248 ][ 361 ],
   alphaCSR[ 248 ][ 362 ],
   alphaCSR[ 248 ][ 363 ],
   alphaCSR[ 248 ][ 364 ],
   alphaCSR[ 248 ][ 365 ],
   alphaCSR[ 248 ][ 366 ],
   alphaCSR[ 248 ][ 367 ],
   alphaCSR[ 248 ][ 368 ],
   alphaCSR[ 248 ][ 369 ],
   alphaCSR[ 248 ][ 370 ],
   alphaCSR[ 248 ][ 371 ],
   alphaCSR[ 248 ][ 372 ],
   alphaCSR[ 248 ][ 373 ],
   alphaCSR[ 248 ][ 374 ],
   alphaCSR[ 248 ][ 375 ],
   alphaCSR[ 248 ][ 376 ],
   alphaCSR[ 248 ][ 377 ],
   alphaCSR[ 248 ][ 378 ],
   alphaCSR[ 248 ][ 379 ],
   alphaCSR[ 248 ][ 380 ],
   alphaCSR[ 248 ][ 381 ],
   alphaCSR[ 248 ][ 382 ],
   alphaCSR[ 248 ][ 383 ],
   alphaCSR[ 249 ][ 0 ],
   alphaCSR[ 249 ][ 1 ],
   alphaCSR[ 249 ][ 2 ],
   alphaCSR[ 249 ][ 3 ],
   alphaCSR[ 249 ][ 4 ],
   alphaCSR[ 249 ][ 5 ],
   alphaCSR[ 249 ][ 6 ],
   alphaCSR[ 249 ][ 7 ],
   alphaCSR[ 249 ][ 8 ],
   alphaCSR[ 249 ][ 9 ],
   alphaCSR[ 249 ][ 10 ],
   alphaCSR[ 249 ][ 11 ],
   alphaCSR[ 249 ][ 12 ],
   alphaCSR[ 249 ][ 13 ],
   alphaCSR[ 249 ][ 14 ],
   alphaCSR[ 249 ][ 15 ],
   alphaCSR[ 249 ][ 16 ],
   alphaCSR[ 249 ][ 17 ],
   alphaCSR[ 249 ][ 18 ],
   alphaCSR[ 249 ][ 19 ],
   alphaCSR[ 249 ][ 20 ],
   alphaCSR[ 249 ][ 21 ],
   alphaCSR[ 249 ][ 22 ],
   alphaCSR[ 249 ][ 23 ],
   alphaCSR[ 249 ][ 24 ],
   alphaCSR[ 249 ][ 25 ],
   alphaCSR[ 249 ][ 26 ],
   alphaCSR[ 249 ][ 27 ],
   alphaCSR[ 249 ][ 28 ],
   alphaCSR[ 249 ][ 29 ],
   alphaCSR[ 249 ][ 30 ],
   alphaCSR[ 249 ][ 31 ],
   alphaCSR[ 249 ][ 32 ],
   alphaCSR[ 249 ][ 33 ],
   alphaCSR[ 249 ][ 34 ],
   alphaCSR[ 249 ][ 35 ],
   alphaCSR[ 249 ][ 36 ],
   alphaCSR[ 249 ][ 37 ],
   alphaCSR[ 249 ][ 38 ],
   alphaCSR[ 249 ][ 39 ],
   alphaCSR[ 249 ][ 40 ],
   alphaCSR[ 249 ][ 41 ],
   alphaCSR[ 249 ][ 42 ],
   alphaCSR[ 249 ][ 43 ],
   alphaCSR[ 249 ][ 44 ],
   alphaCSR[ 249 ][ 45 ],
   alphaCSR[ 249 ][ 46 ],
   alphaCSR[ 249 ][ 47 ],
   alphaCSR[ 249 ][ 48 ],
   alphaCSR[ 249 ][ 49 ],
   alphaCSR[ 249 ][ 50 ],
   alphaCSR[ 249 ][ 51 ],
   alphaCSR[ 249 ][ 52 ],
   alphaCSR[ 249 ][ 53 ],
   alphaCSR[ 249 ][ 54 ],
   alphaCSR[ 249 ][ 55 ],
   alphaCSR[ 249 ][ 56 ],
   alphaCSR[ 249 ][ 57 ],
   alphaCSR[ 249 ][ 58 ],
   alphaCSR[ 249 ][ 59 ],
   alphaCSR[ 249 ][ 60 ],
   alphaCSR[ 249 ][ 61 ],
   alphaCSR[ 249 ][ 62 ],
   alphaCSR[ 249 ][ 63 ],
   alphaCSR[ 249 ][ 64 ],
   alphaCSR[ 249 ][ 65 ],
   alphaCSR[ 249 ][ 66 ],
   alphaCSR[ 249 ][ 67 ],
   alphaCSR[ 249 ][ 68 ],
   alphaCSR[ 249 ][ 69 ],
   alphaCSR[ 249 ][ 70 ],
   alphaCSR[ 249 ][ 71 ],
   alphaCSR[ 249 ][ 72 ],
   alphaCSR[ 249 ][ 73 ],
   alphaCSR[ 249 ][ 74 ],
   alphaCSR[ 249 ][ 75 ],
   alphaCSR[ 249 ][ 76 ],
   alphaCSR[ 249 ][ 77 ],
   alphaCSR[ 249 ][ 78 ],
   alphaCSR[ 249 ][ 79 ],
   alphaCSR[ 249 ][ 80 ],
   alphaCSR[ 249 ][ 81 ],
   alphaCSR[ 249 ][ 82 ],
   alphaCSR[ 249 ][ 83 ],
   alphaCSR[ 249 ][ 84 ],
   alphaCSR[ 249 ][ 85 ],
   alphaCSR[ 249 ][ 86 ],
   alphaCSR[ 249 ][ 87 ],
   alphaCSR[ 249 ][ 88 ],
   alphaCSR[ 249 ][ 89 ],
   alphaCSR[ 249 ][ 90 ],
   alphaCSR[ 249 ][ 91 ],
   alphaCSR[ 249 ][ 92 ],
   alphaCSR[ 249 ][ 93 ],
   alphaCSR[ 249 ][ 94 ],
   alphaCSR[ 249 ][ 95 ],
   alphaCSR[ 249 ][ 96 ],
   alphaCSR[ 249 ][ 97 ],
   alphaCSR[ 249 ][ 98 ],
   alphaCSR[ 249 ][ 99 ],
   alphaCSR[ 249 ][ 100 ],
   alphaCSR[ 249 ][ 101 ],
   alphaCSR[ 249 ][ 102 ],
   alphaCSR[ 249 ][ 103 ],
   alphaCSR[ 249 ][ 104 ],
   alphaCSR[ 249 ][ 105 ],
   alphaCSR[ 249 ][ 106 ],
   alphaCSR[ 249 ][ 107 ],
   alphaCSR[ 249 ][ 108 ],
   alphaCSR[ 249 ][ 109 ],
   alphaCSR[ 249 ][ 110 ],
   alphaCSR[ 249 ][ 111 ],
   alphaCSR[ 249 ][ 112 ],
   alphaCSR[ 249 ][ 113 ],
   alphaCSR[ 249 ][ 114 ],
   alphaCSR[ 249 ][ 115 ],
   alphaCSR[ 249 ][ 116 ],
   alphaCSR[ 249 ][ 117 ],
   alphaCSR[ 249 ][ 118 ],
   alphaCSR[ 249 ][ 119 ],
   alphaCSR[ 249 ][ 120 ],
   alphaCSR[ 249 ][ 121 ],
   alphaCSR[ 249 ][ 122 ],
   alphaCSR[ 249 ][ 123 ],
   alphaCSR[ 249 ][ 124 ],
   alphaCSR[ 249 ][ 125 ],
   alphaCSR[ 249 ][ 126 ],
   alphaCSR[ 249 ][ 127 ],
   alphaCSR[ 249 ][ 128 ],
   alphaCSR[ 249 ][ 129 ],
   alphaCSR[ 249 ][ 130 ],
   alphaCSR[ 249 ][ 131 ],
   alphaCSR[ 249 ][ 132 ],
   alphaCSR[ 249 ][ 133 ],
   alphaCSR[ 249 ][ 134 ],
   alphaCSR[ 249 ][ 135 ],
   alphaCSR[ 249 ][ 136 ],
   alphaCSR[ 249 ][ 137 ],
   alphaCSR[ 249 ][ 138 ],
   alphaCSR[ 249 ][ 139 ],
   alphaCSR[ 249 ][ 140 ],
   alphaCSR[ 249 ][ 141 ],
   alphaCSR[ 249 ][ 142 ],
   alphaCSR[ 249 ][ 143 ],
   alphaCSR[ 249 ][ 144 ],
   alphaCSR[ 249 ][ 145 ],
   alphaCSR[ 249 ][ 146 ],
   alphaCSR[ 249 ][ 147 ],
   alphaCSR[ 249 ][ 148 ],
   alphaCSR[ 249 ][ 149 ],
   alphaCSR[ 249 ][ 150 ],
   alphaCSR[ 249 ][ 151 ],
   alphaCSR[ 249 ][ 152 ],
   alphaCSR[ 249 ][ 153 ],
   alphaCSR[ 249 ][ 154 ],
   alphaCSR[ 249 ][ 155 ],
   alphaCSR[ 249 ][ 156 ],
   alphaCSR[ 249 ][ 157 ],
   alphaCSR[ 249 ][ 158 ],
   alphaCSR[ 249 ][ 159 ],
   alphaCSR[ 249 ][ 160 ],
   alphaCSR[ 249 ][ 161 ],
   alphaCSR[ 249 ][ 162 ],
   alphaCSR[ 249 ][ 163 ],
   alphaCSR[ 249 ][ 164 ],
   alphaCSR[ 249 ][ 165 ],
   alphaCSR[ 249 ][ 166 ],
   alphaCSR[ 249 ][ 167 ],
   alphaCSR[ 249 ][ 168 ],
   alphaCSR[ 249 ][ 169 ],
   alphaCSR[ 249 ][ 170 ],
   alphaCSR[ 249 ][ 171 ],
   alphaCSR[ 249 ][ 172 ],
   alphaCSR[ 249 ][ 173 ],
   alphaCSR[ 249 ][ 174 ],
   alphaCSR[ 249 ][ 175 ],
   alphaCSR[ 249 ][ 176 ],
   alphaCSR[ 249 ][ 177 ],
   alphaCSR[ 249 ][ 178 ],
   alphaCSR[ 249 ][ 179 ],
   alphaCSR[ 249 ][ 180 ],
   alphaCSR[ 249 ][ 181 ],
   alphaCSR[ 249 ][ 182 ],
   alphaCSR[ 249 ][ 183 ],
   alphaCSR[ 249 ][ 184 ],
   alphaCSR[ 249 ][ 185 ],
   alphaCSR[ 249 ][ 186 ],
   alphaCSR[ 249 ][ 187 ],
   alphaCSR[ 249 ][ 188 ],
   alphaCSR[ 249 ][ 189 ],
   alphaCSR[ 249 ][ 190 ],
   alphaCSR[ 249 ][ 191 ],
   alphaCSR[ 249 ][ 192 ],
   alphaCSR[ 249 ][ 193 ],
   alphaCSR[ 249 ][ 194 ],
   alphaCSR[ 249 ][ 195 ],
   alphaCSR[ 249 ][ 196 ],
   alphaCSR[ 249 ][ 197 ],
   alphaCSR[ 249 ][ 198 ],
   alphaCSR[ 249 ][ 199 ],
   alphaCSR[ 249 ][ 200 ],
   alphaCSR[ 249 ][ 201 ],
   alphaCSR[ 249 ][ 202 ],
   alphaCSR[ 249 ][ 203 ],
   alphaCSR[ 249 ][ 204 ],
   alphaCSR[ 249 ][ 205 ],
   alphaCSR[ 249 ][ 206 ],
   alphaCSR[ 249 ][ 207 ],
   alphaCSR[ 249 ][ 208 ],
   alphaCSR[ 249 ][ 209 ],
   alphaCSR[ 249 ][ 210 ],
   alphaCSR[ 249 ][ 211 ],
   alphaCSR[ 249 ][ 212 ],
   alphaCSR[ 249 ][ 213 ],
   alphaCSR[ 249 ][ 214 ],
   alphaCSR[ 249 ][ 215 ],
   alphaCSR[ 249 ][ 216 ],
   alphaCSR[ 249 ][ 217 ],
   alphaCSR[ 249 ][ 218 ],
   alphaCSR[ 249 ][ 219 ],
   alphaCSR[ 249 ][ 220 ],
   alphaCSR[ 249 ][ 221 ],
   alphaCSR[ 249 ][ 222 ],
   alphaCSR[ 249 ][ 223 ],
   alphaCSR[ 249 ][ 224 ],
   alphaCSR[ 249 ][ 225 ],
   alphaCSR[ 249 ][ 226 ],
   alphaCSR[ 249 ][ 227 ],
   alphaCSR[ 249 ][ 228 ],
   alphaCSR[ 249 ][ 229 ],
   alphaCSR[ 249 ][ 230 ],
   alphaCSR[ 249 ][ 231 ],
   alphaCSR[ 249 ][ 232 ],
   alphaCSR[ 249 ][ 233 ],
   alphaCSR[ 249 ][ 234 ],
   alphaCSR[ 249 ][ 235 ],
   alphaCSR[ 249 ][ 236 ],
   alphaCSR[ 249 ][ 237 ],
   alphaCSR[ 249 ][ 238 ],
   alphaCSR[ 249 ][ 239 ],
   alphaCSR[ 249 ][ 240 ],
   alphaCSR[ 249 ][ 241 ],
   alphaCSR[ 249 ][ 242 ],
   alphaCSR[ 249 ][ 243 ],
   alphaCSR[ 249 ][ 244 ],
   alphaCSR[ 249 ][ 245 ],
   alphaCSR[ 249 ][ 246 ],
   alphaCSR[ 249 ][ 247 ],
   alphaCSR[ 249 ][ 248 ],
   alphaCSR[ 249 ][ 249 ],
   alphaCSR[ 249 ][ 250 ],
   alphaCSR[ 249 ][ 251 ],
   alphaCSR[ 249 ][ 252 ],
   alphaCSR[ 249 ][ 253 ],
   alphaCSR[ 249 ][ 254 ],
   alphaCSR[ 249 ][ 255 ],
   alphaCSR[ 249 ][ 256 ],
   alphaCSR[ 249 ][ 257 ],
   alphaCSR[ 249 ][ 258 ],
   alphaCSR[ 249 ][ 259 ],
   alphaCSR[ 249 ][ 260 ],
   alphaCSR[ 249 ][ 261 ],
   alphaCSR[ 249 ][ 262 ],
   alphaCSR[ 249 ][ 263 ],
   alphaCSR[ 249 ][ 264 ],
   alphaCSR[ 249 ][ 265 ],
   alphaCSR[ 249 ][ 266 ],
   alphaCSR[ 249 ][ 267 ],
   alphaCSR[ 249 ][ 268 ],
   alphaCSR[ 249 ][ 269 ],
   alphaCSR[ 249 ][ 270 ],
   alphaCSR[ 249 ][ 271 ],
   alphaCSR[ 249 ][ 272 ],
   alphaCSR[ 249 ][ 273 ],
   alphaCSR[ 249 ][ 274 ],
   alphaCSR[ 249 ][ 275 ],
   alphaCSR[ 249 ][ 276 ],
   alphaCSR[ 249 ][ 277 ],
   alphaCSR[ 249 ][ 278 ],
   alphaCSR[ 249 ][ 279 ],
   alphaCSR[ 249 ][ 280 ],
   alphaCSR[ 249 ][ 281 ],
   alphaCSR[ 249 ][ 282 ],
   alphaCSR[ 249 ][ 283 ],
   alphaCSR[ 249 ][ 284 ],
   alphaCSR[ 249 ][ 285 ],
   alphaCSR[ 249 ][ 286 ],
   alphaCSR[ 249 ][ 287 ],
   alphaCSR[ 249 ][ 288 ],
   alphaCSR[ 249 ][ 289 ],
   alphaCSR[ 249 ][ 290 ],
   alphaCSR[ 249 ][ 291 ],
   alphaCSR[ 249 ][ 292 ],
   alphaCSR[ 249 ][ 293 ],
   alphaCSR[ 249 ][ 294 ],
   alphaCSR[ 249 ][ 295 ],
   alphaCSR[ 249 ][ 296 ],
   alphaCSR[ 249 ][ 297 ],
   alphaCSR[ 249 ][ 298 ],
   alphaCSR[ 249 ][ 299 ],
   alphaCSR[ 249 ][ 300 ],
   alphaCSR[ 249 ][ 301 ],
   alphaCSR[ 249 ][ 302 ],
   alphaCSR[ 249 ][ 303 ],
   alphaCSR[ 249 ][ 304 ],
   alphaCSR[ 249 ][ 305 ],
   alphaCSR[ 249 ][ 306 ],
   alphaCSR[ 249 ][ 307 ],
   alphaCSR[ 249 ][ 308 ],
   alphaCSR[ 249 ][ 309 ],
   alphaCSR[ 249 ][ 310 ],
   alphaCSR[ 249 ][ 311 ],
   alphaCSR[ 249 ][ 312 ],
   alphaCSR[ 249 ][ 313 ],
   alphaCSR[ 249 ][ 314 ],
   alphaCSR[ 249 ][ 315 ],
   alphaCSR[ 249 ][ 316 ],
   alphaCSR[ 249 ][ 317 ],
   alphaCSR[ 249 ][ 318 ],
   alphaCSR[ 249 ][ 319 ],
   alphaCSR[ 249 ][ 320 ],
   alphaCSR[ 249 ][ 321 ],
   alphaCSR[ 249 ][ 322 ],
   alphaCSR[ 249 ][ 323 ],
   alphaCSR[ 249 ][ 324 ],
   alphaCSR[ 249 ][ 325 ],
   alphaCSR[ 249 ][ 326 ],
   alphaCSR[ 249 ][ 327 ],
   alphaCSR[ 249 ][ 328 ],
   alphaCSR[ 249 ][ 329 ],
   alphaCSR[ 249 ][ 330 ],
   alphaCSR[ 249 ][ 331 ],
   alphaCSR[ 249 ][ 332 ],
   alphaCSR[ 249 ][ 333 ],
   alphaCSR[ 249 ][ 334 ],
   alphaCSR[ 249 ][ 335 ],
   alphaCSR[ 249 ][ 336 ],
   alphaCSR[ 249 ][ 337 ],
   alphaCSR[ 249 ][ 338 ],
   alphaCSR[ 249 ][ 339 ],
   alphaCSR[ 249 ][ 340 ],
   alphaCSR[ 249 ][ 341 ],
   alphaCSR[ 249 ][ 342 ],
   alphaCSR[ 249 ][ 343 ],
   alphaCSR[ 249 ][ 344 ],
   alphaCSR[ 249 ][ 345 ],
   alphaCSR[ 249 ][ 346 ],
   alphaCSR[ 249 ][ 347 ],
   alphaCSR[ 249 ][ 348 ],
   alphaCSR[ 249 ][ 349 ],
   alphaCSR[ 249 ][ 350 ],
   alphaCSR[ 249 ][ 351 ],
   alphaCSR[ 249 ][ 352 ],
   alphaCSR[ 249 ][ 353 ],
   alphaCSR[ 249 ][ 354 ],
   alphaCSR[ 249 ][ 355 ],
   alphaCSR[ 249 ][ 356 ],
   alphaCSR[ 249 ][ 357 ],
   alphaCSR[ 249 ][ 358 ],
   alphaCSR[ 249 ][ 359 ],
   alphaCSR[ 249 ][ 360 ],
   alphaCSR[ 249 ][ 361 ],
   alphaCSR[ 249 ][ 362 ],
   alphaCSR[ 249 ][ 363 ],
   alphaCSR[ 249 ][ 364 ],
   alphaCSR[ 249 ][ 365 ],
   alphaCSR[ 249 ][ 366 ],
   alphaCSR[ 249 ][ 367 ],
   alphaCSR[ 249 ][ 368 ],
   alphaCSR[ 249 ][ 369 ],
   alphaCSR[ 249 ][ 370 ],
   alphaCSR[ 249 ][ 371 ],
   alphaCSR[ 249 ][ 372 ],
   alphaCSR[ 249 ][ 373 ],
   alphaCSR[ 249 ][ 374 ],
   alphaCSR[ 249 ][ 375 ],
   alphaCSR[ 249 ][ 376 ],
   alphaCSR[ 249 ][ 377 ],
   alphaCSR[ 249 ][ 378 ],
   alphaCSR[ 249 ][ 379 ],
   alphaCSR[ 249 ][ 380 ],
   alphaCSR[ 249 ][ 381 ],
   alphaCSR[ 249 ][ 382 ],
   alphaCSR[ 249 ][ 383 ],
   alphaCSR[ 250 ][ 0 ],
   alphaCSR[ 250 ][ 1 ],
   alphaCSR[ 250 ][ 2 ],
   alphaCSR[ 250 ][ 3 ],
   alphaCSR[ 250 ][ 4 ],
   alphaCSR[ 250 ][ 5 ],
   alphaCSR[ 250 ][ 6 ],
   alphaCSR[ 250 ][ 7 ],
   alphaCSR[ 250 ][ 8 ],
   alphaCSR[ 250 ][ 9 ],
   alphaCSR[ 250 ][ 10 ],
   alphaCSR[ 250 ][ 11 ],
   alphaCSR[ 250 ][ 12 ],
   alphaCSR[ 250 ][ 13 ],
   alphaCSR[ 250 ][ 14 ],
   alphaCSR[ 250 ][ 15 ],
   alphaCSR[ 250 ][ 16 ],
   alphaCSR[ 250 ][ 17 ],
   alphaCSR[ 250 ][ 18 ],
   alphaCSR[ 250 ][ 19 ],
   alphaCSR[ 250 ][ 20 ],
   alphaCSR[ 250 ][ 21 ],
   alphaCSR[ 250 ][ 22 ],
   alphaCSR[ 250 ][ 23 ],
   alphaCSR[ 250 ][ 24 ],
   alphaCSR[ 250 ][ 25 ],
   alphaCSR[ 250 ][ 26 ],
   alphaCSR[ 250 ][ 27 ],
   alphaCSR[ 250 ][ 28 ],
   alphaCSR[ 250 ][ 29 ],
   alphaCSR[ 250 ][ 30 ],
   alphaCSR[ 250 ][ 31 ],
   alphaCSR[ 250 ][ 32 ],
   alphaCSR[ 250 ][ 33 ],
   alphaCSR[ 250 ][ 34 ],
   alphaCSR[ 250 ][ 35 ],
   alphaCSR[ 250 ][ 36 ],
   alphaCSR[ 250 ][ 37 ],
   alphaCSR[ 250 ][ 38 ],
   alphaCSR[ 250 ][ 39 ],
   alphaCSR[ 250 ][ 40 ],
   alphaCSR[ 250 ][ 41 ],
   alphaCSR[ 250 ][ 42 ],
   alphaCSR[ 250 ][ 43 ],
   alphaCSR[ 250 ][ 44 ],
   alphaCSR[ 250 ][ 45 ],
   alphaCSR[ 250 ][ 46 ],
   alphaCSR[ 250 ][ 47 ],
   alphaCSR[ 250 ][ 48 ],
   alphaCSR[ 250 ][ 49 ],
   alphaCSR[ 250 ][ 50 ],
   alphaCSR[ 250 ][ 51 ],
   alphaCSR[ 250 ][ 52 ],
   alphaCSR[ 250 ][ 53 ],
   alphaCSR[ 250 ][ 54 ],
   alphaCSR[ 250 ][ 55 ],
   alphaCSR[ 250 ][ 56 ],
   alphaCSR[ 250 ][ 57 ],
   alphaCSR[ 250 ][ 58 ],
   alphaCSR[ 250 ][ 59 ],
   alphaCSR[ 250 ][ 60 ],
   alphaCSR[ 250 ][ 61 ],
   alphaCSR[ 250 ][ 62 ],
   alphaCSR[ 250 ][ 63 ],
   alphaCSR[ 250 ][ 64 ],
   alphaCSR[ 250 ][ 65 ],
   alphaCSR[ 250 ][ 66 ],
   alphaCSR[ 250 ][ 67 ],
   alphaCSR[ 250 ][ 68 ],
   alphaCSR[ 250 ][ 69 ],
   alphaCSR[ 250 ][ 70 ],
   alphaCSR[ 250 ][ 71 ],
   alphaCSR[ 250 ][ 72 ],
   alphaCSR[ 250 ][ 73 ],
   alphaCSR[ 250 ][ 74 ],
   alphaCSR[ 250 ][ 75 ],
   alphaCSR[ 250 ][ 76 ],
   alphaCSR[ 250 ][ 77 ],
   alphaCSR[ 250 ][ 78 ],
   alphaCSR[ 250 ][ 79 ],
   alphaCSR[ 250 ][ 80 ],
   alphaCSR[ 250 ][ 81 ],
   alphaCSR[ 250 ][ 82 ],
   alphaCSR[ 250 ][ 83 ],
   alphaCSR[ 250 ][ 84 ],
   alphaCSR[ 250 ][ 85 ],
   alphaCSR[ 250 ][ 86 ],
   alphaCSR[ 250 ][ 87 ],
   alphaCSR[ 250 ][ 88 ],
   alphaCSR[ 250 ][ 89 ],
   alphaCSR[ 250 ][ 90 ],
   alphaCSR[ 250 ][ 91 ],
   alphaCSR[ 250 ][ 92 ],
   alphaCSR[ 250 ][ 93 ],
   alphaCSR[ 250 ][ 94 ],
   alphaCSR[ 250 ][ 95 ],
   alphaCSR[ 250 ][ 96 ],
   alphaCSR[ 250 ][ 97 ],
   alphaCSR[ 250 ][ 98 ],
   alphaCSR[ 250 ][ 99 ],
   alphaCSR[ 250 ][ 100 ],
   alphaCSR[ 250 ][ 101 ],
   alphaCSR[ 250 ][ 102 ],
   alphaCSR[ 250 ][ 103 ],
   alphaCSR[ 250 ][ 104 ],
   alphaCSR[ 250 ][ 105 ],
   alphaCSR[ 250 ][ 106 ],
   alphaCSR[ 250 ][ 107 ],
   alphaCSR[ 250 ][ 108 ],
   alphaCSR[ 250 ][ 109 ],
   alphaCSR[ 250 ][ 110 ],
   alphaCSR[ 250 ][ 111 ],
   alphaCSR[ 250 ][ 112 ],
   alphaCSR[ 250 ][ 113 ],
   alphaCSR[ 250 ][ 114 ],
   alphaCSR[ 250 ][ 115 ],
   alphaCSR[ 250 ][ 116 ],
   alphaCSR[ 250 ][ 117 ],
   alphaCSR[ 250 ][ 118 ],
   alphaCSR[ 250 ][ 119 ],
   alphaCSR[ 250 ][ 120 ],
   alphaCSR[ 250 ][ 121 ],
   alphaCSR[ 250 ][ 122 ],
   alphaCSR[ 250 ][ 123 ],
   alphaCSR[ 250 ][ 124 ],
   alphaCSR[ 250 ][ 125 ],
   alphaCSR[ 250 ][ 126 ],
   alphaCSR[ 250 ][ 127 ],
   alphaCSR[ 250 ][ 128 ],
   alphaCSR[ 250 ][ 129 ],
   alphaCSR[ 250 ][ 130 ],
   alphaCSR[ 250 ][ 131 ],
   alphaCSR[ 250 ][ 132 ],
   alphaCSR[ 250 ][ 133 ],
   alphaCSR[ 250 ][ 134 ],
   alphaCSR[ 250 ][ 135 ],
   alphaCSR[ 250 ][ 136 ],
   alphaCSR[ 250 ][ 137 ],
   alphaCSR[ 250 ][ 138 ],
   alphaCSR[ 250 ][ 139 ],
   alphaCSR[ 250 ][ 140 ],
   alphaCSR[ 250 ][ 141 ],
   alphaCSR[ 250 ][ 142 ],
   alphaCSR[ 250 ][ 143 ],
   alphaCSR[ 250 ][ 144 ],
   alphaCSR[ 250 ][ 145 ],
   alphaCSR[ 250 ][ 146 ],
   alphaCSR[ 250 ][ 147 ],
   alphaCSR[ 250 ][ 148 ],
   alphaCSR[ 250 ][ 149 ],
   alphaCSR[ 250 ][ 150 ],
   alphaCSR[ 250 ][ 151 ],
   alphaCSR[ 250 ][ 152 ],
   alphaCSR[ 250 ][ 153 ],
   alphaCSR[ 250 ][ 154 ],
   alphaCSR[ 250 ][ 155 ],
   alphaCSR[ 250 ][ 156 ],
   alphaCSR[ 250 ][ 157 ],
   alphaCSR[ 250 ][ 158 ],
   alphaCSR[ 250 ][ 159 ],
   alphaCSR[ 250 ][ 160 ],
   alphaCSR[ 250 ][ 161 ],
   alphaCSR[ 250 ][ 162 ],
   alphaCSR[ 250 ][ 163 ],
   alphaCSR[ 250 ][ 164 ],
   alphaCSR[ 250 ][ 165 ],
   alphaCSR[ 250 ][ 166 ],
   alphaCSR[ 250 ][ 167 ],
   alphaCSR[ 250 ][ 168 ],
   alphaCSR[ 250 ][ 169 ],
   alphaCSR[ 250 ][ 170 ],
   alphaCSR[ 250 ][ 171 ],
   alphaCSR[ 250 ][ 172 ],
   alphaCSR[ 250 ][ 173 ],
   alphaCSR[ 250 ][ 174 ],
   alphaCSR[ 250 ][ 175 ],
   alphaCSR[ 250 ][ 176 ],
   alphaCSR[ 250 ][ 177 ],
   alphaCSR[ 250 ][ 178 ],
   alphaCSR[ 250 ][ 179 ],
   alphaCSR[ 250 ][ 180 ],
   alphaCSR[ 250 ][ 181 ],
   alphaCSR[ 250 ][ 182 ],
   alphaCSR[ 250 ][ 183 ],
   alphaCSR[ 250 ][ 184 ],
   alphaCSR[ 250 ][ 185 ],
   alphaCSR[ 250 ][ 186 ],
   alphaCSR[ 250 ][ 187 ],
   alphaCSR[ 250 ][ 188 ],
   alphaCSR[ 250 ][ 189 ],
   alphaCSR[ 250 ][ 190 ],
   alphaCSR[ 250 ][ 191 ],
   alphaCSR[ 250 ][ 192 ],
   alphaCSR[ 250 ][ 193 ],
   alphaCSR[ 250 ][ 194 ],
   alphaCSR[ 250 ][ 195 ],
   alphaCSR[ 250 ][ 196 ],
   alphaCSR[ 250 ][ 197 ],
   alphaCSR[ 250 ][ 198 ],
   alphaCSR[ 250 ][ 199 ],
   alphaCSR[ 250 ][ 200 ],
   alphaCSR[ 250 ][ 201 ],
   alphaCSR[ 250 ][ 202 ],
   alphaCSR[ 250 ][ 203 ],
   alphaCSR[ 250 ][ 204 ],
   alphaCSR[ 250 ][ 205 ],
   alphaCSR[ 250 ][ 206 ],
   alphaCSR[ 250 ][ 207 ],
   alphaCSR[ 250 ][ 208 ],
   alphaCSR[ 250 ][ 209 ],
   alphaCSR[ 250 ][ 210 ],
   alphaCSR[ 250 ][ 211 ],
   alphaCSR[ 250 ][ 212 ],
   alphaCSR[ 250 ][ 213 ],
   alphaCSR[ 250 ][ 214 ],
   alphaCSR[ 250 ][ 215 ],
   alphaCSR[ 250 ][ 216 ],
   alphaCSR[ 250 ][ 217 ],
   alphaCSR[ 250 ][ 218 ],
   alphaCSR[ 250 ][ 219 ],
   alphaCSR[ 250 ][ 220 ],
   alphaCSR[ 250 ][ 221 ],
   alphaCSR[ 250 ][ 222 ],
   alphaCSR[ 250 ][ 223 ],
   alphaCSR[ 250 ][ 224 ],
   alphaCSR[ 250 ][ 225 ],
   alphaCSR[ 250 ][ 226 ],
   alphaCSR[ 250 ][ 227 ],
   alphaCSR[ 250 ][ 228 ],
   alphaCSR[ 250 ][ 229 ],
   alphaCSR[ 250 ][ 230 ],
   alphaCSR[ 250 ][ 231 ],
   alphaCSR[ 250 ][ 232 ],
   alphaCSR[ 250 ][ 233 ],
   alphaCSR[ 250 ][ 234 ],
   alphaCSR[ 250 ][ 235 ],
   alphaCSR[ 250 ][ 236 ],
   alphaCSR[ 250 ][ 237 ],
   alphaCSR[ 250 ][ 238 ],
   alphaCSR[ 250 ][ 239 ],
   alphaCSR[ 250 ][ 240 ],
   alphaCSR[ 250 ][ 241 ],
   alphaCSR[ 250 ][ 242 ],
   alphaCSR[ 250 ][ 243 ],
   alphaCSR[ 250 ][ 244 ],
   alphaCSR[ 250 ][ 245 ],
   alphaCSR[ 250 ][ 246 ],
   alphaCSR[ 250 ][ 247 ],
   alphaCSR[ 250 ][ 248 ],
   alphaCSR[ 250 ][ 249 ],
   alphaCSR[ 250 ][ 250 ],
   alphaCSR[ 250 ][ 251 ],
   alphaCSR[ 250 ][ 252 ],
   alphaCSR[ 250 ][ 253 ],
   alphaCSR[ 250 ][ 254 ],
   alphaCSR[ 250 ][ 255 ],
   alphaCSR[ 250 ][ 256 ],
   alphaCSR[ 250 ][ 257 ],
   alphaCSR[ 250 ][ 258 ],
   alphaCSR[ 250 ][ 259 ],
   alphaCSR[ 250 ][ 260 ],
   alphaCSR[ 250 ][ 261 ],
   alphaCSR[ 250 ][ 262 ],
   alphaCSR[ 250 ][ 263 ],
   alphaCSR[ 250 ][ 264 ],
   alphaCSR[ 250 ][ 265 ],
   alphaCSR[ 250 ][ 266 ],
   alphaCSR[ 250 ][ 267 ],
   alphaCSR[ 250 ][ 268 ],
   alphaCSR[ 250 ][ 269 ],
   alphaCSR[ 250 ][ 270 ],
   alphaCSR[ 250 ][ 271 ],
   alphaCSR[ 250 ][ 272 ],
   alphaCSR[ 250 ][ 273 ],
   alphaCSR[ 250 ][ 274 ],
   alphaCSR[ 250 ][ 275 ],
   alphaCSR[ 250 ][ 276 ],
   alphaCSR[ 250 ][ 277 ],
   alphaCSR[ 250 ][ 278 ],
   alphaCSR[ 250 ][ 279 ],
   alphaCSR[ 250 ][ 280 ],
   alphaCSR[ 250 ][ 281 ],
   alphaCSR[ 250 ][ 282 ],
   alphaCSR[ 250 ][ 283 ],
   alphaCSR[ 250 ][ 284 ],
   alphaCSR[ 250 ][ 285 ],
   alphaCSR[ 250 ][ 286 ],
   alphaCSR[ 250 ][ 287 ],
   alphaCSR[ 250 ][ 288 ],
   alphaCSR[ 250 ][ 289 ],
   alphaCSR[ 250 ][ 290 ],
   alphaCSR[ 250 ][ 291 ],
   alphaCSR[ 250 ][ 292 ],
   alphaCSR[ 250 ][ 293 ],
   alphaCSR[ 250 ][ 294 ],
   alphaCSR[ 250 ][ 295 ],
   alphaCSR[ 250 ][ 296 ],
   alphaCSR[ 250 ][ 297 ],
   alphaCSR[ 250 ][ 298 ],
   alphaCSR[ 250 ][ 299 ],
   alphaCSR[ 250 ][ 300 ],
   alphaCSR[ 250 ][ 301 ],
   alphaCSR[ 250 ][ 302 ],
   alphaCSR[ 250 ][ 303 ],
   alphaCSR[ 250 ][ 304 ],
   alphaCSR[ 250 ][ 305 ],
   alphaCSR[ 250 ][ 306 ],
   alphaCSR[ 250 ][ 307 ],
   alphaCSR[ 250 ][ 308 ],
   alphaCSR[ 250 ][ 309 ],
   alphaCSR[ 250 ][ 310 ],
   alphaCSR[ 250 ][ 311 ],
   alphaCSR[ 250 ][ 312 ],
   alphaCSR[ 250 ][ 313 ],
   alphaCSR[ 250 ][ 314 ],
   alphaCSR[ 250 ][ 315 ],
   alphaCSR[ 250 ][ 316 ],
   alphaCSR[ 250 ][ 317 ],
   alphaCSR[ 250 ][ 318 ],
   alphaCSR[ 250 ][ 319 ],
   alphaCSR[ 250 ][ 320 ],
   alphaCSR[ 250 ][ 321 ],
   alphaCSR[ 250 ][ 322 ],
   alphaCSR[ 250 ][ 323 ],
   alphaCSR[ 250 ][ 324 ],
   alphaCSR[ 250 ][ 325 ],
   alphaCSR[ 250 ][ 326 ],
   alphaCSR[ 250 ][ 327 ],
   alphaCSR[ 250 ][ 328 ],
   alphaCSR[ 250 ][ 329 ],
   alphaCSR[ 250 ][ 330 ],
   alphaCSR[ 250 ][ 331 ],
   alphaCSR[ 250 ][ 332 ],
   alphaCSR[ 250 ][ 333 ],
   alphaCSR[ 250 ][ 334 ],
   alphaCSR[ 250 ][ 335 ],
   alphaCSR[ 250 ][ 336 ],
   alphaCSR[ 250 ][ 337 ],
   alphaCSR[ 250 ][ 338 ],
   alphaCSR[ 250 ][ 339 ],
   alphaCSR[ 250 ][ 340 ],
   alphaCSR[ 250 ][ 341 ],
   alphaCSR[ 250 ][ 342 ],
   alphaCSR[ 250 ][ 343 ],
   alphaCSR[ 250 ][ 344 ],
   alphaCSR[ 250 ][ 345 ],
   alphaCSR[ 250 ][ 346 ],
   alphaCSR[ 250 ][ 347 ],
   alphaCSR[ 250 ][ 348 ],
   alphaCSR[ 250 ][ 349 ],
   alphaCSR[ 250 ][ 350 ],
   alphaCSR[ 250 ][ 351 ],
   alphaCSR[ 250 ][ 352 ],
   alphaCSR[ 250 ][ 353 ],
   alphaCSR[ 250 ][ 354 ],
   alphaCSR[ 250 ][ 355 ],
   alphaCSR[ 250 ][ 356 ],
   alphaCSR[ 250 ][ 357 ],
   alphaCSR[ 250 ][ 358 ],
   alphaCSR[ 250 ][ 359 ],
   alphaCSR[ 250 ][ 360 ],
   alphaCSR[ 250 ][ 361 ],
   alphaCSR[ 250 ][ 362 ],
   alphaCSR[ 250 ][ 363 ],
   alphaCSR[ 250 ][ 364 ],
   alphaCSR[ 250 ][ 365 ],
   alphaCSR[ 250 ][ 366 ],
   alphaCSR[ 250 ][ 367 ],
   alphaCSR[ 250 ][ 368 ],
   alphaCSR[ 250 ][ 369 ],
   alphaCSR[ 250 ][ 370 ],
   alphaCSR[ 250 ][ 371 ],
   alphaCSR[ 250 ][ 372 ],
   alphaCSR[ 250 ][ 373 ],
   alphaCSR[ 250 ][ 374 ],
   alphaCSR[ 250 ][ 375 ],
   alphaCSR[ 250 ][ 376 ],
   alphaCSR[ 250 ][ 377 ],
   alphaCSR[ 250 ][ 378 ],
   alphaCSR[ 250 ][ 379 ],
   alphaCSR[ 250 ][ 380 ],
   alphaCSR[ 250 ][ 381 ],
   alphaCSR[ 250 ][ 382 ],
   alphaCSR[ 250 ][ 383 ],
   alphaCSR[ 251 ][ 0 ],
   alphaCSR[ 251 ][ 1 ],
   alphaCSR[ 251 ][ 2 ],
   alphaCSR[ 251 ][ 3 ],
   alphaCSR[ 251 ][ 4 ],
   alphaCSR[ 251 ][ 5 ],
   alphaCSR[ 251 ][ 6 ],
   alphaCSR[ 251 ][ 7 ],
   alphaCSR[ 251 ][ 8 ],
   alphaCSR[ 251 ][ 9 ],
   alphaCSR[ 251 ][ 10 ],
   alphaCSR[ 251 ][ 11 ],
   alphaCSR[ 251 ][ 12 ],
   alphaCSR[ 251 ][ 13 ],
   alphaCSR[ 251 ][ 14 ],
   alphaCSR[ 251 ][ 15 ],
   alphaCSR[ 251 ][ 16 ],
   alphaCSR[ 251 ][ 17 ],
   alphaCSR[ 251 ][ 18 ],
   alphaCSR[ 251 ][ 19 ],
   alphaCSR[ 251 ][ 20 ],
   alphaCSR[ 251 ][ 21 ],
   alphaCSR[ 251 ][ 22 ],
   alphaCSR[ 251 ][ 23 ],
   alphaCSR[ 251 ][ 24 ],
   alphaCSR[ 251 ][ 25 ],
   alphaCSR[ 251 ][ 26 ],
   alphaCSR[ 251 ][ 27 ],
   alphaCSR[ 251 ][ 28 ],
   alphaCSR[ 251 ][ 29 ],
   alphaCSR[ 251 ][ 30 ],
   alphaCSR[ 251 ][ 31 ],
   alphaCSR[ 251 ][ 32 ],
   alphaCSR[ 251 ][ 33 ],
   alphaCSR[ 251 ][ 34 ],
   alphaCSR[ 251 ][ 35 ],
   alphaCSR[ 251 ][ 36 ],
   alphaCSR[ 251 ][ 37 ],
   alphaCSR[ 251 ][ 38 ],
   alphaCSR[ 251 ][ 39 ],
   alphaCSR[ 251 ][ 40 ],
   alphaCSR[ 251 ][ 41 ],
   alphaCSR[ 251 ][ 42 ],
   alphaCSR[ 251 ][ 43 ],
   alphaCSR[ 251 ][ 44 ],
   alphaCSR[ 251 ][ 45 ],
   alphaCSR[ 251 ][ 46 ],
   alphaCSR[ 251 ][ 47 ],
   alphaCSR[ 251 ][ 48 ],
   alphaCSR[ 251 ][ 49 ],
   alphaCSR[ 251 ][ 50 ],
   alphaCSR[ 251 ][ 51 ],
   alphaCSR[ 251 ][ 52 ],
   alphaCSR[ 251 ][ 53 ],
   alphaCSR[ 251 ][ 54 ],
   alphaCSR[ 251 ][ 55 ],
   alphaCSR[ 251 ][ 56 ],
   alphaCSR[ 251 ][ 57 ],
   alphaCSR[ 251 ][ 58 ],
   alphaCSR[ 251 ][ 59 ],
   alphaCSR[ 251 ][ 60 ],
   alphaCSR[ 251 ][ 61 ],
   alphaCSR[ 251 ][ 62 ],
   alphaCSR[ 251 ][ 63 ],
   alphaCSR[ 251 ][ 64 ],
   alphaCSR[ 251 ][ 65 ],
   alphaCSR[ 251 ][ 66 ],
   alphaCSR[ 251 ][ 67 ],
   alphaCSR[ 251 ][ 68 ],
   alphaCSR[ 251 ][ 69 ],
   alphaCSR[ 251 ][ 70 ],
   alphaCSR[ 251 ][ 71 ],
   alphaCSR[ 251 ][ 72 ],
   alphaCSR[ 251 ][ 73 ],
   alphaCSR[ 251 ][ 74 ],
   alphaCSR[ 251 ][ 75 ],
   alphaCSR[ 251 ][ 76 ],
   alphaCSR[ 251 ][ 77 ],
   alphaCSR[ 251 ][ 78 ],
   alphaCSR[ 251 ][ 79 ],
   alphaCSR[ 251 ][ 80 ],
   alphaCSR[ 251 ][ 81 ],
   alphaCSR[ 251 ][ 82 ],
   alphaCSR[ 251 ][ 83 ],
   alphaCSR[ 251 ][ 84 ],
   alphaCSR[ 251 ][ 85 ],
   alphaCSR[ 251 ][ 86 ],
   alphaCSR[ 251 ][ 87 ],
   alphaCSR[ 251 ][ 88 ],
   alphaCSR[ 251 ][ 89 ],
   alphaCSR[ 251 ][ 90 ],
   alphaCSR[ 251 ][ 91 ],
   alphaCSR[ 251 ][ 92 ],
   alphaCSR[ 251 ][ 93 ],
   alphaCSR[ 251 ][ 94 ],
   alphaCSR[ 251 ][ 95 ],
   alphaCSR[ 251 ][ 96 ],
   alphaCSR[ 251 ][ 97 ],
   alphaCSR[ 251 ][ 98 ],
   alphaCSR[ 251 ][ 99 ],
   alphaCSR[ 251 ][ 100 ],
   alphaCSR[ 251 ][ 101 ],
   alphaCSR[ 251 ][ 102 ],
   alphaCSR[ 251 ][ 103 ],
   alphaCSR[ 251 ][ 104 ],
   alphaCSR[ 251 ][ 105 ],
   alphaCSR[ 251 ][ 106 ],
   alphaCSR[ 251 ][ 107 ],
   alphaCSR[ 251 ][ 108 ],
   alphaCSR[ 251 ][ 109 ],
   alphaCSR[ 251 ][ 110 ],
   alphaCSR[ 251 ][ 111 ],
   alphaCSR[ 251 ][ 112 ],
   alphaCSR[ 251 ][ 113 ],
   alphaCSR[ 251 ][ 114 ],
   alphaCSR[ 251 ][ 115 ],
   alphaCSR[ 251 ][ 116 ],
   alphaCSR[ 251 ][ 117 ],
   alphaCSR[ 251 ][ 118 ],
   alphaCSR[ 251 ][ 119 ],
   alphaCSR[ 251 ][ 120 ],
   alphaCSR[ 251 ][ 121 ],
   alphaCSR[ 251 ][ 122 ],
   alphaCSR[ 251 ][ 123 ],
   alphaCSR[ 251 ][ 124 ],
   alphaCSR[ 251 ][ 125 ],
   alphaCSR[ 251 ][ 126 ],
   alphaCSR[ 251 ][ 127 ],
   alphaCSR[ 251 ][ 128 ],
   alphaCSR[ 251 ][ 129 ],
   alphaCSR[ 251 ][ 130 ],
   alphaCSR[ 251 ][ 131 ],
   alphaCSR[ 251 ][ 132 ],
   alphaCSR[ 251 ][ 133 ],
   alphaCSR[ 251 ][ 134 ],
   alphaCSR[ 251 ][ 135 ],
   alphaCSR[ 251 ][ 136 ],
   alphaCSR[ 251 ][ 137 ],
   alphaCSR[ 251 ][ 138 ],
   alphaCSR[ 251 ][ 139 ],
   alphaCSR[ 251 ][ 140 ],
   alphaCSR[ 251 ][ 141 ],
   alphaCSR[ 251 ][ 142 ],
   alphaCSR[ 251 ][ 143 ],
   alphaCSR[ 251 ][ 144 ],
   alphaCSR[ 251 ][ 145 ],
   alphaCSR[ 251 ][ 146 ],
   alphaCSR[ 251 ][ 147 ],
   alphaCSR[ 251 ][ 148 ],
   alphaCSR[ 251 ][ 149 ],
   alphaCSR[ 251 ][ 150 ],
   alphaCSR[ 251 ][ 151 ],
   alphaCSR[ 251 ][ 152 ],
   alphaCSR[ 251 ][ 153 ],
   alphaCSR[ 251 ][ 154 ],
   alphaCSR[ 251 ][ 155 ],
   alphaCSR[ 251 ][ 156 ],
   alphaCSR[ 251 ][ 157 ],
   alphaCSR[ 251 ][ 158 ],
   alphaCSR[ 251 ][ 159 ],
   alphaCSR[ 251 ][ 160 ],
   alphaCSR[ 251 ][ 161 ],
   alphaCSR[ 251 ][ 162 ],
   alphaCSR[ 251 ][ 163 ],
   alphaCSR[ 251 ][ 164 ],
   alphaCSR[ 251 ][ 165 ],
   alphaCSR[ 251 ][ 166 ],
   alphaCSR[ 251 ][ 167 ],
   alphaCSR[ 251 ][ 168 ],
   alphaCSR[ 251 ][ 169 ],
   alphaCSR[ 251 ][ 170 ],
   alphaCSR[ 251 ][ 171 ],
   alphaCSR[ 251 ][ 172 ],
   alphaCSR[ 251 ][ 173 ],
   alphaCSR[ 251 ][ 174 ],
   alphaCSR[ 251 ][ 175 ],
   alphaCSR[ 251 ][ 176 ],
   alphaCSR[ 251 ][ 177 ],
   alphaCSR[ 251 ][ 178 ],
   alphaCSR[ 251 ][ 179 ],
   alphaCSR[ 251 ][ 180 ],
   alphaCSR[ 251 ][ 181 ],
   alphaCSR[ 251 ][ 182 ],
   alphaCSR[ 251 ][ 183 ],
   alphaCSR[ 251 ][ 184 ],
   alphaCSR[ 251 ][ 185 ],
   alphaCSR[ 251 ][ 186 ],
   alphaCSR[ 251 ][ 187 ],
   alphaCSR[ 251 ][ 188 ],
   alphaCSR[ 251 ][ 189 ],
   alphaCSR[ 251 ][ 190 ],
   alphaCSR[ 251 ][ 191 ],
   alphaCSR[ 251 ][ 192 ],
   alphaCSR[ 251 ][ 193 ],
   alphaCSR[ 251 ][ 194 ],
   alphaCSR[ 251 ][ 195 ],
   alphaCSR[ 251 ][ 196 ],
   alphaCSR[ 251 ][ 197 ],
   alphaCSR[ 251 ][ 198 ],
   alphaCSR[ 251 ][ 199 ],
   alphaCSR[ 251 ][ 200 ],
   alphaCSR[ 251 ][ 201 ],
   alphaCSR[ 251 ][ 202 ],
   alphaCSR[ 251 ][ 203 ],
   alphaCSR[ 251 ][ 204 ],
   alphaCSR[ 251 ][ 205 ],
   alphaCSR[ 251 ][ 206 ],
   alphaCSR[ 251 ][ 207 ],
   alphaCSR[ 251 ][ 208 ],
   alphaCSR[ 251 ][ 209 ],
   alphaCSR[ 251 ][ 210 ],
   alphaCSR[ 251 ][ 211 ],
   alphaCSR[ 251 ][ 212 ],
   alphaCSR[ 251 ][ 213 ],
   alphaCSR[ 251 ][ 214 ],
   alphaCSR[ 251 ][ 215 ],
   alphaCSR[ 251 ][ 216 ],
   alphaCSR[ 251 ][ 217 ],
   alphaCSR[ 251 ][ 218 ],
   alphaCSR[ 251 ][ 219 ],
   alphaCSR[ 251 ][ 220 ],
   alphaCSR[ 251 ][ 221 ],
   alphaCSR[ 251 ][ 222 ],
   alphaCSR[ 251 ][ 223 ],
   alphaCSR[ 251 ][ 224 ],
   alphaCSR[ 251 ][ 225 ],
   alphaCSR[ 251 ][ 226 ],
   alphaCSR[ 251 ][ 227 ],
   alphaCSR[ 251 ][ 228 ],
   alphaCSR[ 251 ][ 229 ],
   alphaCSR[ 251 ][ 230 ],
   alphaCSR[ 251 ][ 231 ],
   alphaCSR[ 251 ][ 232 ],
   alphaCSR[ 251 ][ 233 ],
   alphaCSR[ 251 ][ 234 ],
   alphaCSR[ 251 ][ 235 ],
   alphaCSR[ 251 ][ 236 ],
   alphaCSR[ 251 ][ 237 ],
   alphaCSR[ 251 ][ 238 ],
   alphaCSR[ 251 ][ 239 ],
   alphaCSR[ 251 ][ 240 ],
   alphaCSR[ 251 ][ 241 ],
   alphaCSR[ 251 ][ 242 ],
   alphaCSR[ 251 ][ 243 ],
   alphaCSR[ 251 ][ 244 ],
   alphaCSR[ 251 ][ 245 ],
   alphaCSR[ 251 ][ 246 ],
   alphaCSR[ 251 ][ 247 ],
   alphaCSR[ 251 ][ 248 ],
   alphaCSR[ 251 ][ 249 ],
   alphaCSR[ 251 ][ 250 ],
   alphaCSR[ 251 ][ 251 ],
   alphaCSR[ 251 ][ 252 ],
   alphaCSR[ 251 ][ 253 ],
   alphaCSR[ 251 ][ 254 ],
   alphaCSR[ 251 ][ 255 ],
   alphaCSR[ 251 ][ 256 ],
   alphaCSR[ 251 ][ 257 ],
   alphaCSR[ 251 ][ 258 ],
   alphaCSR[ 251 ][ 259 ],
   alphaCSR[ 251 ][ 260 ],
   alphaCSR[ 251 ][ 261 ],
   alphaCSR[ 251 ][ 262 ],
   alphaCSR[ 251 ][ 263 ],
   alphaCSR[ 251 ][ 264 ],
   alphaCSR[ 251 ][ 265 ],
   alphaCSR[ 251 ][ 266 ],
   alphaCSR[ 251 ][ 267 ],
   alphaCSR[ 251 ][ 268 ],
   alphaCSR[ 251 ][ 269 ],
   alphaCSR[ 251 ][ 270 ],
   alphaCSR[ 251 ][ 271 ],
   alphaCSR[ 251 ][ 272 ],
   alphaCSR[ 251 ][ 273 ],
   alphaCSR[ 251 ][ 274 ],
   alphaCSR[ 251 ][ 275 ],
   alphaCSR[ 251 ][ 276 ],
   alphaCSR[ 251 ][ 277 ],
   alphaCSR[ 251 ][ 278 ],
   alphaCSR[ 251 ][ 279 ],
   alphaCSR[ 251 ][ 280 ],
   alphaCSR[ 251 ][ 281 ],
   alphaCSR[ 251 ][ 282 ],
   alphaCSR[ 251 ][ 283 ],
   alphaCSR[ 251 ][ 284 ],
   alphaCSR[ 251 ][ 285 ],
   alphaCSR[ 251 ][ 286 ],
   alphaCSR[ 251 ][ 287 ],
   alphaCSR[ 251 ][ 288 ],
   alphaCSR[ 251 ][ 289 ],
   alphaCSR[ 251 ][ 290 ],
   alphaCSR[ 251 ][ 291 ],
   alphaCSR[ 251 ][ 292 ],
   alphaCSR[ 251 ][ 293 ],
   alphaCSR[ 251 ][ 294 ],
   alphaCSR[ 251 ][ 295 ],
   alphaCSR[ 251 ][ 296 ],
   alphaCSR[ 251 ][ 297 ],
   alphaCSR[ 251 ][ 298 ],
   alphaCSR[ 251 ][ 299 ],
   alphaCSR[ 251 ][ 300 ],
   alphaCSR[ 251 ][ 301 ],
   alphaCSR[ 251 ][ 302 ],
   alphaCSR[ 251 ][ 303 ],
   alphaCSR[ 251 ][ 304 ],
   alphaCSR[ 251 ][ 305 ],
   alphaCSR[ 251 ][ 306 ],
   alphaCSR[ 251 ][ 307 ],
   alphaCSR[ 251 ][ 308 ],
   alphaCSR[ 251 ][ 309 ],
   alphaCSR[ 251 ][ 310 ],
   alphaCSR[ 251 ][ 311 ],
   alphaCSR[ 251 ][ 312 ],
   alphaCSR[ 251 ][ 313 ],
   alphaCSR[ 251 ][ 314 ],
   alphaCSR[ 251 ][ 315 ],
   alphaCSR[ 251 ][ 316 ],
   alphaCSR[ 251 ][ 317 ],
   alphaCSR[ 251 ][ 318 ],
   alphaCSR[ 251 ][ 319 ],
   alphaCSR[ 251 ][ 320 ],
   alphaCSR[ 251 ][ 321 ],
   alphaCSR[ 251 ][ 322 ],
   alphaCSR[ 251 ][ 323 ],
   alphaCSR[ 251 ][ 324 ],
   alphaCSR[ 251 ][ 325 ],
   alphaCSR[ 251 ][ 326 ],
   alphaCSR[ 251 ][ 327 ],
   alphaCSR[ 251 ][ 328 ],
   alphaCSR[ 251 ][ 329 ],
   alphaCSR[ 251 ][ 330 ],
   alphaCSR[ 251 ][ 331 ],
   alphaCSR[ 251 ][ 332 ],
   alphaCSR[ 251 ][ 333 ],
   alphaCSR[ 251 ][ 334 ],
   alphaCSR[ 251 ][ 335 ],
   alphaCSR[ 251 ][ 336 ],
   alphaCSR[ 251 ][ 337 ],
   alphaCSR[ 251 ][ 338 ],
   alphaCSR[ 251 ][ 339 ],
   alphaCSR[ 251 ][ 340 ],
   alphaCSR[ 251 ][ 341 ],
   alphaCSR[ 251 ][ 342 ],
   alphaCSR[ 251 ][ 343 ],
   alphaCSR[ 251 ][ 344 ],
   alphaCSR[ 251 ][ 345 ],
   alphaCSR[ 251 ][ 346 ],
   alphaCSR[ 251 ][ 347 ],
   alphaCSR[ 251 ][ 348 ],
   alphaCSR[ 251 ][ 349 ],
   alphaCSR[ 251 ][ 350 ],
   alphaCSR[ 251 ][ 351 ],
   alphaCSR[ 251 ][ 352 ],
   alphaCSR[ 251 ][ 353 ],
   alphaCSR[ 251 ][ 354 ],
   alphaCSR[ 251 ][ 355 ],
   alphaCSR[ 251 ][ 356 ],
   alphaCSR[ 251 ][ 357 ],
   alphaCSR[ 251 ][ 358 ],
   alphaCSR[ 251 ][ 359 ],
   alphaCSR[ 251 ][ 360 ],
   alphaCSR[ 251 ][ 361 ],
   alphaCSR[ 251 ][ 362 ],
   alphaCSR[ 251 ][ 363 ],
   alphaCSR[ 251 ][ 364 ],
   alphaCSR[ 251 ][ 365 ],
   alphaCSR[ 251 ][ 366 ],
   alphaCSR[ 251 ][ 367 ],
   alphaCSR[ 251 ][ 368 ],
   alphaCSR[ 251 ][ 369 ],
   alphaCSR[ 251 ][ 370 ],
   alphaCSR[ 251 ][ 371 ],
   alphaCSR[ 251 ][ 372 ],
   alphaCSR[ 251 ][ 373 ],
   alphaCSR[ 251 ][ 374 ],
   alphaCSR[ 251 ][ 375 ],
   alphaCSR[ 251 ][ 376 ],
   alphaCSR[ 251 ][ 377 ],
   alphaCSR[ 251 ][ 378 ],
   alphaCSR[ 251 ][ 379 ],
   alphaCSR[ 251 ][ 380 ],
   alphaCSR[ 251 ][ 381 ],
   alphaCSR[ 251 ][ 382 ],
   alphaCSR[ 251 ][ 383 ],
   alphaCSR[ 252 ][ 0 ],
   alphaCSR[ 252 ][ 1 ],
   alphaCSR[ 252 ][ 2 ],
   alphaCSR[ 252 ][ 3 ],
   alphaCSR[ 252 ][ 4 ],
   alphaCSR[ 252 ][ 5 ],
   alphaCSR[ 252 ][ 6 ],
   alphaCSR[ 252 ][ 7 ],
   alphaCSR[ 252 ][ 8 ],
   alphaCSR[ 252 ][ 9 ],
   alphaCSR[ 252 ][ 10 ],
   alphaCSR[ 252 ][ 11 ],
   alphaCSR[ 252 ][ 12 ],
   alphaCSR[ 252 ][ 13 ],
   alphaCSR[ 252 ][ 14 ],
   alphaCSR[ 252 ][ 15 ],
   alphaCSR[ 252 ][ 16 ],
   alphaCSR[ 252 ][ 17 ],
   alphaCSR[ 252 ][ 18 ],
   alphaCSR[ 252 ][ 19 ],
   alphaCSR[ 252 ][ 20 ],
   alphaCSR[ 252 ][ 21 ],
   alphaCSR[ 252 ][ 22 ],
   alphaCSR[ 252 ][ 23 ],
   alphaCSR[ 252 ][ 24 ],
   alphaCSR[ 252 ][ 25 ],
   alphaCSR[ 252 ][ 26 ],
   alphaCSR[ 252 ][ 27 ],
   alphaCSR[ 252 ][ 28 ],
   alphaCSR[ 252 ][ 29 ],
   alphaCSR[ 252 ][ 30 ],
   alphaCSR[ 252 ][ 31 ],
   alphaCSR[ 252 ][ 32 ],
   alphaCSR[ 252 ][ 33 ],
   alphaCSR[ 252 ][ 34 ],
   alphaCSR[ 252 ][ 35 ],
   alphaCSR[ 252 ][ 36 ],
   alphaCSR[ 252 ][ 37 ],
   alphaCSR[ 252 ][ 38 ],
   alphaCSR[ 252 ][ 39 ],
   alphaCSR[ 252 ][ 40 ],
   alphaCSR[ 252 ][ 41 ],
   alphaCSR[ 252 ][ 42 ],
   alphaCSR[ 252 ][ 43 ],
   alphaCSR[ 252 ][ 44 ],
   alphaCSR[ 252 ][ 45 ],
   alphaCSR[ 252 ][ 46 ],
   alphaCSR[ 252 ][ 47 ],
   alphaCSR[ 252 ][ 48 ],
   alphaCSR[ 252 ][ 49 ],
   alphaCSR[ 252 ][ 50 ],
   alphaCSR[ 252 ][ 51 ],
   alphaCSR[ 252 ][ 52 ],
   alphaCSR[ 252 ][ 53 ],
   alphaCSR[ 252 ][ 54 ],
   alphaCSR[ 252 ][ 55 ],
   alphaCSR[ 252 ][ 56 ],
   alphaCSR[ 252 ][ 57 ],
   alphaCSR[ 252 ][ 58 ],
   alphaCSR[ 252 ][ 59 ],
   alphaCSR[ 252 ][ 60 ],
   alphaCSR[ 252 ][ 61 ],
   alphaCSR[ 252 ][ 62 ],
   alphaCSR[ 252 ][ 63 ],
   alphaCSR[ 252 ][ 64 ],
   alphaCSR[ 252 ][ 65 ],
   alphaCSR[ 252 ][ 66 ],
   alphaCSR[ 252 ][ 67 ],
   alphaCSR[ 252 ][ 68 ],
   alphaCSR[ 252 ][ 69 ],
   alphaCSR[ 252 ][ 70 ],
   alphaCSR[ 252 ][ 71 ],
   alphaCSR[ 252 ][ 72 ],
   alphaCSR[ 252 ][ 73 ],
   alphaCSR[ 252 ][ 74 ],
   alphaCSR[ 252 ][ 75 ],
   alphaCSR[ 252 ][ 76 ],
   alphaCSR[ 252 ][ 77 ],
   alphaCSR[ 252 ][ 78 ],
   alphaCSR[ 252 ][ 79 ],
   alphaCSR[ 252 ][ 80 ],
   alphaCSR[ 252 ][ 81 ],
   alphaCSR[ 252 ][ 82 ],
   alphaCSR[ 252 ][ 83 ],
   alphaCSR[ 252 ][ 84 ],
   alphaCSR[ 252 ][ 85 ],
   alphaCSR[ 252 ][ 86 ],
   alphaCSR[ 252 ][ 87 ],
   alphaCSR[ 252 ][ 88 ],
   alphaCSR[ 252 ][ 89 ],
   alphaCSR[ 252 ][ 90 ],
   alphaCSR[ 252 ][ 91 ],
   alphaCSR[ 252 ][ 92 ],
   alphaCSR[ 252 ][ 93 ],
   alphaCSR[ 252 ][ 94 ],
   alphaCSR[ 252 ][ 95 ],
   alphaCSR[ 252 ][ 96 ],
   alphaCSR[ 252 ][ 97 ],
   alphaCSR[ 252 ][ 98 ],
   alphaCSR[ 252 ][ 99 ],
   alphaCSR[ 252 ][ 100 ],
   alphaCSR[ 252 ][ 101 ],
   alphaCSR[ 252 ][ 102 ],
   alphaCSR[ 252 ][ 103 ],
   alphaCSR[ 252 ][ 104 ],
   alphaCSR[ 252 ][ 105 ],
   alphaCSR[ 252 ][ 106 ],
   alphaCSR[ 252 ][ 107 ],
   alphaCSR[ 252 ][ 108 ],
   alphaCSR[ 252 ][ 109 ],
   alphaCSR[ 252 ][ 110 ],
   alphaCSR[ 252 ][ 111 ],
   alphaCSR[ 252 ][ 112 ],
   alphaCSR[ 252 ][ 113 ],
   alphaCSR[ 252 ][ 114 ],
   alphaCSR[ 252 ][ 115 ],
   alphaCSR[ 252 ][ 116 ],
   alphaCSR[ 252 ][ 117 ],
   alphaCSR[ 252 ][ 118 ],
   alphaCSR[ 252 ][ 119 ],
   alphaCSR[ 252 ][ 120 ],
   alphaCSR[ 252 ][ 121 ],
   alphaCSR[ 252 ][ 122 ],
   alphaCSR[ 252 ][ 123 ],
   alphaCSR[ 252 ][ 124 ],
   alphaCSR[ 252 ][ 125 ],
   alphaCSR[ 252 ][ 126 ],
   alphaCSR[ 252 ][ 127 ],
   alphaCSR[ 252 ][ 128 ],
   alphaCSR[ 252 ][ 129 ],
   alphaCSR[ 252 ][ 130 ],
   alphaCSR[ 252 ][ 131 ],
   alphaCSR[ 252 ][ 132 ],
   alphaCSR[ 252 ][ 133 ],
   alphaCSR[ 252 ][ 134 ],
   alphaCSR[ 252 ][ 135 ],
   alphaCSR[ 252 ][ 136 ],
   alphaCSR[ 252 ][ 137 ],
   alphaCSR[ 252 ][ 138 ],
   alphaCSR[ 252 ][ 139 ],
   alphaCSR[ 252 ][ 140 ],
   alphaCSR[ 252 ][ 141 ],
   alphaCSR[ 252 ][ 142 ],
   alphaCSR[ 252 ][ 143 ],
   alphaCSR[ 252 ][ 144 ],
   alphaCSR[ 252 ][ 145 ],
   alphaCSR[ 252 ][ 146 ],
   alphaCSR[ 252 ][ 147 ],
   alphaCSR[ 252 ][ 148 ],
   alphaCSR[ 252 ][ 149 ],
   alphaCSR[ 252 ][ 150 ],
   alphaCSR[ 252 ][ 151 ],
   alphaCSR[ 252 ][ 152 ],
   alphaCSR[ 252 ][ 153 ],
   alphaCSR[ 252 ][ 154 ],
   alphaCSR[ 252 ][ 155 ],
   alphaCSR[ 252 ][ 156 ],
   alphaCSR[ 252 ][ 157 ],
   alphaCSR[ 252 ][ 158 ],
   alphaCSR[ 252 ][ 159 ],
   alphaCSR[ 252 ][ 160 ],
   alphaCSR[ 252 ][ 161 ],
   alphaCSR[ 252 ][ 162 ],
   alphaCSR[ 252 ][ 163 ],
   alphaCSR[ 252 ][ 164 ],
   alphaCSR[ 252 ][ 165 ],
   alphaCSR[ 252 ][ 166 ],
   alphaCSR[ 252 ][ 167 ],
   alphaCSR[ 252 ][ 168 ],
   alphaCSR[ 252 ][ 169 ],
   alphaCSR[ 252 ][ 170 ],
   alphaCSR[ 252 ][ 171 ],
   alphaCSR[ 252 ][ 172 ],
   alphaCSR[ 252 ][ 173 ],
   alphaCSR[ 252 ][ 174 ],
   alphaCSR[ 252 ][ 175 ],
   alphaCSR[ 252 ][ 176 ],
   alphaCSR[ 252 ][ 177 ],
   alphaCSR[ 252 ][ 178 ],
   alphaCSR[ 252 ][ 179 ],
   alphaCSR[ 252 ][ 180 ],
   alphaCSR[ 252 ][ 181 ],
   alphaCSR[ 252 ][ 182 ],
   alphaCSR[ 252 ][ 183 ],
   alphaCSR[ 252 ][ 184 ],
   alphaCSR[ 252 ][ 185 ],
   alphaCSR[ 252 ][ 186 ],
   alphaCSR[ 252 ][ 187 ],
   alphaCSR[ 252 ][ 188 ],
   alphaCSR[ 252 ][ 189 ],
   alphaCSR[ 252 ][ 190 ],
   alphaCSR[ 252 ][ 191 ],
   alphaCSR[ 252 ][ 192 ],
   alphaCSR[ 252 ][ 193 ],
   alphaCSR[ 252 ][ 194 ],
   alphaCSR[ 252 ][ 195 ],
   alphaCSR[ 252 ][ 196 ],
   alphaCSR[ 252 ][ 197 ],
   alphaCSR[ 252 ][ 198 ],
   alphaCSR[ 252 ][ 199 ],
   alphaCSR[ 252 ][ 200 ],
   alphaCSR[ 252 ][ 201 ],
   alphaCSR[ 252 ][ 202 ],
   alphaCSR[ 252 ][ 203 ],
   alphaCSR[ 252 ][ 204 ],
   alphaCSR[ 252 ][ 205 ],
   alphaCSR[ 252 ][ 206 ],
   alphaCSR[ 252 ][ 207 ],
   alphaCSR[ 252 ][ 208 ],
   alphaCSR[ 252 ][ 209 ],
   alphaCSR[ 252 ][ 210 ],
   alphaCSR[ 252 ][ 211 ],
   alphaCSR[ 252 ][ 212 ],
   alphaCSR[ 252 ][ 213 ],
   alphaCSR[ 252 ][ 214 ],
   alphaCSR[ 252 ][ 215 ],
   alphaCSR[ 252 ][ 216 ],
   alphaCSR[ 252 ][ 217 ],
   alphaCSR[ 252 ][ 218 ],
   alphaCSR[ 252 ][ 219 ],
   alphaCSR[ 252 ][ 220 ],
   alphaCSR[ 252 ][ 221 ],
   alphaCSR[ 252 ][ 222 ],
   alphaCSR[ 252 ][ 223 ],
   alphaCSR[ 252 ][ 224 ],
   alphaCSR[ 252 ][ 225 ],
   alphaCSR[ 252 ][ 226 ],
   alphaCSR[ 252 ][ 227 ],
   alphaCSR[ 252 ][ 228 ],
   alphaCSR[ 252 ][ 229 ],
   alphaCSR[ 252 ][ 230 ],
   alphaCSR[ 252 ][ 231 ],
   alphaCSR[ 252 ][ 232 ],
   alphaCSR[ 252 ][ 233 ],
   alphaCSR[ 252 ][ 234 ],
   alphaCSR[ 252 ][ 235 ],
   alphaCSR[ 252 ][ 236 ],
   alphaCSR[ 252 ][ 237 ],
   alphaCSR[ 252 ][ 238 ],
   alphaCSR[ 252 ][ 239 ],
   alphaCSR[ 252 ][ 240 ],
   alphaCSR[ 252 ][ 241 ],
   alphaCSR[ 252 ][ 242 ],
   alphaCSR[ 252 ][ 243 ],
   alphaCSR[ 252 ][ 244 ],
   alphaCSR[ 252 ][ 245 ],
   alphaCSR[ 252 ][ 246 ],
   alphaCSR[ 252 ][ 247 ],
   alphaCSR[ 252 ][ 248 ],
   alphaCSR[ 252 ][ 249 ],
   alphaCSR[ 252 ][ 250 ],
   alphaCSR[ 252 ][ 251 ],
   alphaCSR[ 252 ][ 252 ],
   alphaCSR[ 252 ][ 253 ],
   alphaCSR[ 252 ][ 254 ],
   alphaCSR[ 252 ][ 255 ],
   alphaCSR[ 252 ][ 256 ],
   alphaCSR[ 252 ][ 257 ],
   alphaCSR[ 252 ][ 258 ],
   alphaCSR[ 252 ][ 259 ],
   alphaCSR[ 252 ][ 260 ],
   alphaCSR[ 252 ][ 261 ],
   alphaCSR[ 252 ][ 262 ],
   alphaCSR[ 252 ][ 263 ],
   alphaCSR[ 252 ][ 264 ],
   alphaCSR[ 252 ][ 265 ],
   alphaCSR[ 252 ][ 266 ],
   alphaCSR[ 252 ][ 267 ],
   alphaCSR[ 252 ][ 268 ],
   alphaCSR[ 252 ][ 269 ],
   alphaCSR[ 252 ][ 270 ],
   alphaCSR[ 252 ][ 271 ],
   alphaCSR[ 252 ][ 272 ],
   alphaCSR[ 252 ][ 273 ],
   alphaCSR[ 252 ][ 274 ],
   alphaCSR[ 252 ][ 275 ],
   alphaCSR[ 252 ][ 276 ],
   alphaCSR[ 252 ][ 277 ],
   alphaCSR[ 252 ][ 278 ],
   alphaCSR[ 252 ][ 279 ],
   alphaCSR[ 252 ][ 280 ],
   alphaCSR[ 252 ][ 281 ],
   alphaCSR[ 252 ][ 282 ],
   alphaCSR[ 252 ][ 283 ],
   alphaCSR[ 252 ][ 284 ],
   alphaCSR[ 252 ][ 285 ],
   alphaCSR[ 252 ][ 286 ],
   alphaCSR[ 252 ][ 287 ],
   alphaCSR[ 252 ][ 288 ],
   alphaCSR[ 252 ][ 289 ],
   alphaCSR[ 252 ][ 290 ],
   alphaCSR[ 252 ][ 291 ],
   alphaCSR[ 252 ][ 292 ],
   alphaCSR[ 252 ][ 293 ],
   alphaCSR[ 252 ][ 294 ],
   alphaCSR[ 252 ][ 295 ],
   alphaCSR[ 252 ][ 296 ],
   alphaCSR[ 252 ][ 297 ],
   alphaCSR[ 252 ][ 298 ],
   alphaCSR[ 252 ][ 299 ],
   alphaCSR[ 252 ][ 300 ],
   alphaCSR[ 252 ][ 301 ],
   alphaCSR[ 252 ][ 302 ],
   alphaCSR[ 252 ][ 303 ],
   alphaCSR[ 252 ][ 304 ],
   alphaCSR[ 252 ][ 305 ],
   alphaCSR[ 252 ][ 306 ],
   alphaCSR[ 252 ][ 307 ],
   alphaCSR[ 252 ][ 308 ],
   alphaCSR[ 252 ][ 309 ],
   alphaCSR[ 252 ][ 310 ],
   alphaCSR[ 252 ][ 311 ],
   alphaCSR[ 252 ][ 312 ],
   alphaCSR[ 252 ][ 313 ],
   alphaCSR[ 252 ][ 314 ],
   alphaCSR[ 252 ][ 315 ],
   alphaCSR[ 252 ][ 316 ],
   alphaCSR[ 252 ][ 317 ],
   alphaCSR[ 252 ][ 318 ],
   alphaCSR[ 252 ][ 319 ],
   alphaCSR[ 252 ][ 320 ],
   alphaCSR[ 252 ][ 321 ],
   alphaCSR[ 252 ][ 322 ],
   alphaCSR[ 252 ][ 323 ],
   alphaCSR[ 252 ][ 324 ],
   alphaCSR[ 252 ][ 325 ],
   alphaCSR[ 252 ][ 326 ],
   alphaCSR[ 252 ][ 327 ],
   alphaCSR[ 252 ][ 328 ],
   alphaCSR[ 252 ][ 329 ],
   alphaCSR[ 252 ][ 330 ],
   alphaCSR[ 252 ][ 331 ],
   alphaCSR[ 252 ][ 332 ],
   alphaCSR[ 252 ][ 333 ],
   alphaCSR[ 252 ][ 334 ],
   alphaCSR[ 252 ][ 335 ],
   alphaCSR[ 252 ][ 336 ],
   alphaCSR[ 252 ][ 337 ],
   alphaCSR[ 252 ][ 338 ],
   alphaCSR[ 252 ][ 339 ],
   alphaCSR[ 252 ][ 340 ],
   alphaCSR[ 252 ][ 341 ],
   alphaCSR[ 252 ][ 342 ],
   alphaCSR[ 252 ][ 343 ],
   alphaCSR[ 252 ][ 344 ],
   alphaCSR[ 252 ][ 345 ],
   alphaCSR[ 252 ][ 346 ],
   alphaCSR[ 252 ][ 347 ],
   alphaCSR[ 252 ][ 348 ],
   alphaCSR[ 252 ][ 349 ],
   alphaCSR[ 252 ][ 350 ],
   alphaCSR[ 252 ][ 351 ],
   alphaCSR[ 252 ][ 352 ],
   alphaCSR[ 252 ][ 353 ],
   alphaCSR[ 252 ][ 354 ],
   alphaCSR[ 252 ][ 355 ],
   alphaCSR[ 252 ][ 356 ],
   alphaCSR[ 252 ][ 357 ],
   alphaCSR[ 252 ][ 358 ],
   alphaCSR[ 252 ][ 359 ],
   alphaCSR[ 252 ][ 360 ],
   alphaCSR[ 252 ][ 361 ],
   alphaCSR[ 252 ][ 362 ],
   alphaCSR[ 252 ][ 363 ],
   alphaCSR[ 252 ][ 364 ],
   alphaCSR[ 252 ][ 365 ],
   alphaCSR[ 252 ][ 366 ],
   alphaCSR[ 252 ][ 367 ],
   alphaCSR[ 252 ][ 368 ],
   alphaCSR[ 252 ][ 369 ],
   alphaCSR[ 252 ][ 370 ],
   alphaCSR[ 252 ][ 371 ],
   alphaCSR[ 252 ][ 372 ],
   alphaCSR[ 252 ][ 373 ],
   alphaCSR[ 252 ][ 374 ],
   alphaCSR[ 252 ][ 375 ],
   alphaCSR[ 252 ][ 376 ],
   alphaCSR[ 252 ][ 377 ],
   alphaCSR[ 252 ][ 378 ],
   alphaCSR[ 252 ][ 379 ],
   alphaCSR[ 252 ][ 380 ],
   alphaCSR[ 252 ][ 381 ],
   alphaCSR[ 252 ][ 382 ],
   alphaCSR[ 252 ][ 383 ],
   alphaCSR[ 253 ][ 0 ],
   alphaCSR[ 253 ][ 1 ],
   alphaCSR[ 253 ][ 2 ],
   alphaCSR[ 253 ][ 3 ],
   alphaCSR[ 253 ][ 4 ],
   alphaCSR[ 253 ][ 5 ],
   alphaCSR[ 253 ][ 6 ],
   alphaCSR[ 253 ][ 7 ],
   alphaCSR[ 253 ][ 8 ],
   alphaCSR[ 253 ][ 9 ],
   alphaCSR[ 253 ][ 10 ],
   alphaCSR[ 253 ][ 11 ],
   alphaCSR[ 253 ][ 12 ],
   alphaCSR[ 253 ][ 13 ],
   alphaCSR[ 253 ][ 14 ],
   alphaCSR[ 253 ][ 15 ],
   alphaCSR[ 253 ][ 16 ],
   alphaCSR[ 253 ][ 17 ],
   alphaCSR[ 253 ][ 18 ],
   alphaCSR[ 253 ][ 19 ],
   alphaCSR[ 253 ][ 20 ],
   alphaCSR[ 253 ][ 21 ],
   alphaCSR[ 253 ][ 22 ],
   alphaCSR[ 253 ][ 23 ],
   alphaCSR[ 253 ][ 24 ],
   alphaCSR[ 253 ][ 25 ],
   alphaCSR[ 253 ][ 26 ],
   alphaCSR[ 253 ][ 27 ],
   alphaCSR[ 253 ][ 28 ],
   alphaCSR[ 253 ][ 29 ],
   alphaCSR[ 253 ][ 30 ],
   alphaCSR[ 253 ][ 31 ],
   alphaCSR[ 253 ][ 32 ],
   alphaCSR[ 253 ][ 33 ],
   alphaCSR[ 253 ][ 34 ],
   alphaCSR[ 253 ][ 35 ],
   alphaCSR[ 253 ][ 36 ],
   alphaCSR[ 253 ][ 37 ],
   alphaCSR[ 253 ][ 38 ],
   alphaCSR[ 253 ][ 39 ],
   alphaCSR[ 253 ][ 40 ],
   alphaCSR[ 253 ][ 41 ],
   alphaCSR[ 253 ][ 42 ],
   alphaCSR[ 253 ][ 43 ],
   alphaCSR[ 253 ][ 44 ],
   alphaCSR[ 253 ][ 45 ],
   alphaCSR[ 253 ][ 46 ],
   alphaCSR[ 253 ][ 47 ],
   alphaCSR[ 253 ][ 48 ],
   alphaCSR[ 253 ][ 49 ],
   alphaCSR[ 253 ][ 50 ],
   alphaCSR[ 253 ][ 51 ],
   alphaCSR[ 253 ][ 52 ],
   alphaCSR[ 253 ][ 53 ],
   alphaCSR[ 253 ][ 54 ],
   alphaCSR[ 253 ][ 55 ],
   alphaCSR[ 253 ][ 56 ],
   alphaCSR[ 253 ][ 57 ],
   alphaCSR[ 253 ][ 58 ],
   alphaCSR[ 253 ][ 59 ],
   alphaCSR[ 253 ][ 60 ],
   alphaCSR[ 253 ][ 61 ],
   alphaCSR[ 253 ][ 62 ],
   alphaCSR[ 253 ][ 63 ],
   alphaCSR[ 253 ][ 64 ],
   alphaCSR[ 253 ][ 65 ],
   alphaCSR[ 253 ][ 66 ],
   alphaCSR[ 253 ][ 67 ],
   alphaCSR[ 253 ][ 68 ],
   alphaCSR[ 253 ][ 69 ],
   alphaCSR[ 253 ][ 70 ],
   alphaCSR[ 253 ][ 71 ],
   alphaCSR[ 253 ][ 72 ],
   alphaCSR[ 253 ][ 73 ],
   alphaCSR[ 253 ][ 74 ],
   alphaCSR[ 253 ][ 75 ],
   alphaCSR[ 253 ][ 76 ],
   alphaCSR[ 253 ][ 77 ],
   alphaCSR[ 253 ][ 78 ],
   alphaCSR[ 253 ][ 79 ],
   alphaCSR[ 253 ][ 80 ],
   alphaCSR[ 253 ][ 81 ],
   alphaCSR[ 253 ][ 82 ],
   alphaCSR[ 253 ][ 83 ],
   alphaCSR[ 253 ][ 84 ],
   alphaCSR[ 253 ][ 85 ],
   alphaCSR[ 253 ][ 86 ],
   alphaCSR[ 253 ][ 87 ],
   alphaCSR[ 253 ][ 88 ],
   alphaCSR[ 253 ][ 89 ],
   alphaCSR[ 253 ][ 90 ],
   alphaCSR[ 253 ][ 91 ],
   alphaCSR[ 253 ][ 92 ],
   alphaCSR[ 253 ][ 93 ],
   alphaCSR[ 253 ][ 94 ],
   alphaCSR[ 253 ][ 95 ],
   alphaCSR[ 253 ][ 96 ],
   alphaCSR[ 253 ][ 97 ],
   alphaCSR[ 253 ][ 98 ],
   alphaCSR[ 253 ][ 99 ],
   alphaCSR[ 253 ][ 100 ],
   alphaCSR[ 253 ][ 101 ],
   alphaCSR[ 253 ][ 102 ],
   alphaCSR[ 253 ][ 103 ],
   alphaCSR[ 253 ][ 104 ],
   alphaCSR[ 253 ][ 105 ],
   alphaCSR[ 253 ][ 106 ],
   alphaCSR[ 253 ][ 107 ],
   alphaCSR[ 253 ][ 108 ],
   alphaCSR[ 253 ][ 109 ],
   alphaCSR[ 253 ][ 110 ],
   alphaCSR[ 253 ][ 111 ],
   alphaCSR[ 253 ][ 112 ],
   alphaCSR[ 253 ][ 113 ],
   alphaCSR[ 253 ][ 114 ],
   alphaCSR[ 253 ][ 115 ],
   alphaCSR[ 253 ][ 116 ],
   alphaCSR[ 253 ][ 117 ],
   alphaCSR[ 253 ][ 118 ],
   alphaCSR[ 253 ][ 119 ],
   alphaCSR[ 253 ][ 120 ],
   alphaCSR[ 253 ][ 121 ],
   alphaCSR[ 253 ][ 122 ],
   alphaCSR[ 253 ][ 123 ],
   alphaCSR[ 253 ][ 124 ],
   alphaCSR[ 253 ][ 125 ],
   alphaCSR[ 253 ][ 126 ],
   alphaCSR[ 253 ][ 127 ],
   alphaCSR[ 253 ][ 128 ],
   alphaCSR[ 253 ][ 129 ],
   alphaCSR[ 253 ][ 130 ],
   alphaCSR[ 253 ][ 131 ],
   alphaCSR[ 253 ][ 132 ],
   alphaCSR[ 253 ][ 133 ],
   alphaCSR[ 253 ][ 134 ],
   alphaCSR[ 253 ][ 135 ],
   alphaCSR[ 253 ][ 136 ],
   alphaCSR[ 253 ][ 137 ],
   alphaCSR[ 253 ][ 138 ],
   alphaCSR[ 253 ][ 139 ],
   alphaCSR[ 253 ][ 140 ],
   alphaCSR[ 253 ][ 141 ],
   alphaCSR[ 253 ][ 142 ],
   alphaCSR[ 253 ][ 143 ],
   alphaCSR[ 253 ][ 144 ],
   alphaCSR[ 253 ][ 145 ],
   alphaCSR[ 253 ][ 146 ],
   alphaCSR[ 253 ][ 147 ],
   alphaCSR[ 253 ][ 148 ],
   alphaCSR[ 253 ][ 149 ],
   alphaCSR[ 253 ][ 150 ],
   alphaCSR[ 253 ][ 151 ],
   alphaCSR[ 253 ][ 152 ],
   alphaCSR[ 253 ][ 153 ],
   alphaCSR[ 253 ][ 154 ],
   alphaCSR[ 253 ][ 155 ],
   alphaCSR[ 253 ][ 156 ],
   alphaCSR[ 253 ][ 157 ],
   alphaCSR[ 253 ][ 158 ],
   alphaCSR[ 253 ][ 159 ],
   alphaCSR[ 253 ][ 160 ],
   alphaCSR[ 253 ][ 161 ],
   alphaCSR[ 253 ][ 162 ],
   alphaCSR[ 253 ][ 163 ],
   alphaCSR[ 253 ][ 164 ],
   alphaCSR[ 253 ][ 165 ],
   alphaCSR[ 253 ][ 166 ],
   alphaCSR[ 253 ][ 167 ],
   alphaCSR[ 253 ][ 168 ],
   alphaCSR[ 253 ][ 169 ],
   alphaCSR[ 253 ][ 170 ],
   alphaCSR[ 253 ][ 171 ],
   alphaCSR[ 253 ][ 172 ],
   alphaCSR[ 253 ][ 173 ],
   alphaCSR[ 253 ][ 174 ],
   alphaCSR[ 253 ][ 175 ],
   alphaCSR[ 253 ][ 176 ],
   alphaCSR[ 253 ][ 177 ],
   alphaCSR[ 253 ][ 178 ],
   alphaCSR[ 253 ][ 179 ],
   alphaCSR[ 253 ][ 180 ],
   alphaCSR[ 253 ][ 181 ],
   alphaCSR[ 253 ][ 182 ],
   alphaCSR[ 253 ][ 183 ],
   alphaCSR[ 253 ][ 184 ],
   alphaCSR[ 253 ][ 185 ],
   alphaCSR[ 253 ][ 186 ],
   alphaCSR[ 253 ][ 187 ],
   alphaCSR[ 253 ][ 188 ],
   alphaCSR[ 253 ][ 189 ],
   alphaCSR[ 253 ][ 190 ],
   alphaCSR[ 253 ][ 191 ],
   alphaCSR[ 253 ][ 192 ],
   alphaCSR[ 253 ][ 193 ],
   alphaCSR[ 253 ][ 194 ],
   alphaCSR[ 253 ][ 195 ],
   alphaCSR[ 253 ][ 196 ],
   alphaCSR[ 253 ][ 197 ],
   alphaCSR[ 253 ][ 198 ],
   alphaCSR[ 253 ][ 199 ],
   alphaCSR[ 253 ][ 200 ],
   alphaCSR[ 253 ][ 201 ],
   alphaCSR[ 253 ][ 202 ],
   alphaCSR[ 253 ][ 203 ],
   alphaCSR[ 253 ][ 204 ],
   alphaCSR[ 253 ][ 205 ],
   alphaCSR[ 253 ][ 206 ],
   alphaCSR[ 253 ][ 207 ],
   alphaCSR[ 253 ][ 208 ],
   alphaCSR[ 253 ][ 209 ],
   alphaCSR[ 253 ][ 210 ],
   alphaCSR[ 253 ][ 211 ],
   alphaCSR[ 253 ][ 212 ],
   alphaCSR[ 253 ][ 213 ],
   alphaCSR[ 253 ][ 214 ],
   alphaCSR[ 253 ][ 215 ],
   alphaCSR[ 253 ][ 216 ],
   alphaCSR[ 253 ][ 217 ],
   alphaCSR[ 253 ][ 218 ],
   alphaCSR[ 253 ][ 219 ],
   alphaCSR[ 253 ][ 220 ],
   alphaCSR[ 253 ][ 221 ],
   alphaCSR[ 253 ][ 222 ],
   alphaCSR[ 253 ][ 223 ],
   alphaCSR[ 253 ][ 224 ],
   alphaCSR[ 253 ][ 225 ],
   alphaCSR[ 253 ][ 226 ],
   alphaCSR[ 253 ][ 227 ],
   alphaCSR[ 253 ][ 228 ],
   alphaCSR[ 253 ][ 229 ],
   alphaCSR[ 253 ][ 230 ],
   alphaCSR[ 253 ][ 231 ],
   alphaCSR[ 253 ][ 232 ],
   alphaCSR[ 253 ][ 233 ],
   alphaCSR[ 253 ][ 234 ],
   alphaCSR[ 253 ][ 235 ],
   alphaCSR[ 253 ][ 236 ],
   alphaCSR[ 253 ][ 237 ],
   alphaCSR[ 253 ][ 238 ],
   alphaCSR[ 253 ][ 239 ],
   alphaCSR[ 253 ][ 240 ],
   alphaCSR[ 253 ][ 241 ],
   alphaCSR[ 253 ][ 242 ],
   alphaCSR[ 253 ][ 243 ],
   alphaCSR[ 253 ][ 244 ],
   alphaCSR[ 253 ][ 245 ],
   alphaCSR[ 253 ][ 246 ],
   alphaCSR[ 253 ][ 247 ],
   alphaCSR[ 253 ][ 248 ],
   alphaCSR[ 253 ][ 249 ],
   alphaCSR[ 253 ][ 250 ],
   alphaCSR[ 253 ][ 251 ],
   alphaCSR[ 253 ][ 252 ],
   alphaCSR[ 253 ][ 253 ],
   alphaCSR[ 253 ][ 254 ],
   alphaCSR[ 253 ][ 255 ],
   alphaCSR[ 253 ][ 256 ],
   alphaCSR[ 253 ][ 257 ],
   alphaCSR[ 253 ][ 258 ],
   alphaCSR[ 253 ][ 259 ],
   alphaCSR[ 253 ][ 260 ],
   alphaCSR[ 253 ][ 261 ],
   alphaCSR[ 253 ][ 262 ],
   alphaCSR[ 253 ][ 263 ],
   alphaCSR[ 253 ][ 264 ],
   alphaCSR[ 253 ][ 265 ],
   alphaCSR[ 253 ][ 266 ],
   alphaCSR[ 253 ][ 267 ],
   alphaCSR[ 253 ][ 268 ],
   alphaCSR[ 253 ][ 269 ],
   alphaCSR[ 253 ][ 270 ],
   alphaCSR[ 253 ][ 271 ],
   alphaCSR[ 253 ][ 272 ],
   alphaCSR[ 253 ][ 273 ],
   alphaCSR[ 253 ][ 274 ],
   alphaCSR[ 253 ][ 275 ],
   alphaCSR[ 253 ][ 276 ],
   alphaCSR[ 253 ][ 277 ],
   alphaCSR[ 253 ][ 278 ],
   alphaCSR[ 253 ][ 279 ],
   alphaCSR[ 253 ][ 280 ],
   alphaCSR[ 253 ][ 281 ],
   alphaCSR[ 253 ][ 282 ],
   alphaCSR[ 253 ][ 283 ],
   alphaCSR[ 253 ][ 284 ],
   alphaCSR[ 253 ][ 285 ],
   alphaCSR[ 253 ][ 286 ],
   alphaCSR[ 253 ][ 287 ],
   alphaCSR[ 253 ][ 288 ],
   alphaCSR[ 253 ][ 289 ],
   alphaCSR[ 253 ][ 290 ],
   alphaCSR[ 253 ][ 291 ],
   alphaCSR[ 253 ][ 292 ],
   alphaCSR[ 253 ][ 293 ],
   alphaCSR[ 253 ][ 294 ],
   alphaCSR[ 253 ][ 295 ],
   alphaCSR[ 253 ][ 296 ],
   alphaCSR[ 253 ][ 297 ],
   alphaCSR[ 253 ][ 298 ],
   alphaCSR[ 253 ][ 299 ],
   alphaCSR[ 253 ][ 300 ],
   alphaCSR[ 253 ][ 301 ],
   alphaCSR[ 253 ][ 302 ],
   alphaCSR[ 253 ][ 303 ],
   alphaCSR[ 253 ][ 304 ],
   alphaCSR[ 253 ][ 305 ],
   alphaCSR[ 253 ][ 306 ],
   alphaCSR[ 253 ][ 307 ],
   alphaCSR[ 253 ][ 308 ],
   alphaCSR[ 253 ][ 309 ],
   alphaCSR[ 253 ][ 310 ],
   alphaCSR[ 253 ][ 311 ],
   alphaCSR[ 253 ][ 312 ],
   alphaCSR[ 253 ][ 313 ],
   alphaCSR[ 253 ][ 314 ],
   alphaCSR[ 253 ][ 315 ],
   alphaCSR[ 253 ][ 316 ],
   alphaCSR[ 253 ][ 317 ],
   alphaCSR[ 253 ][ 318 ],
   alphaCSR[ 253 ][ 319 ],
   alphaCSR[ 253 ][ 320 ],
   alphaCSR[ 253 ][ 321 ],
   alphaCSR[ 253 ][ 322 ],
   alphaCSR[ 253 ][ 323 ],
   alphaCSR[ 253 ][ 324 ],
   alphaCSR[ 253 ][ 325 ],
   alphaCSR[ 253 ][ 326 ],
   alphaCSR[ 253 ][ 327 ],
   alphaCSR[ 253 ][ 328 ],
   alphaCSR[ 253 ][ 329 ],
   alphaCSR[ 253 ][ 330 ],
   alphaCSR[ 253 ][ 331 ],
   alphaCSR[ 253 ][ 332 ],
   alphaCSR[ 253 ][ 333 ],
   alphaCSR[ 253 ][ 334 ],
   alphaCSR[ 253 ][ 335 ],
   alphaCSR[ 253 ][ 336 ],
   alphaCSR[ 253 ][ 337 ],
   alphaCSR[ 253 ][ 338 ],
   alphaCSR[ 253 ][ 339 ],
   alphaCSR[ 253 ][ 340 ],
   alphaCSR[ 253 ][ 341 ],
   alphaCSR[ 253 ][ 342 ],
   alphaCSR[ 253 ][ 343 ],
   alphaCSR[ 253 ][ 344 ],
   alphaCSR[ 253 ][ 345 ],
   alphaCSR[ 253 ][ 346 ],
   alphaCSR[ 253 ][ 347 ],
   alphaCSR[ 253 ][ 348 ],
   alphaCSR[ 253 ][ 349 ],
   alphaCSR[ 253 ][ 350 ],
   alphaCSR[ 253 ][ 351 ],
   alphaCSR[ 253 ][ 352 ],
   alphaCSR[ 253 ][ 353 ],
   alphaCSR[ 253 ][ 354 ],
   alphaCSR[ 253 ][ 355 ],
   alphaCSR[ 253 ][ 356 ],
   alphaCSR[ 253 ][ 357 ],
   alphaCSR[ 253 ][ 358 ],
   alphaCSR[ 253 ][ 359 ],
   alphaCSR[ 253 ][ 360 ],
   alphaCSR[ 253 ][ 361 ],
   alphaCSR[ 253 ][ 362 ],
   alphaCSR[ 253 ][ 363 ],
   alphaCSR[ 253 ][ 364 ],
   alphaCSR[ 253 ][ 365 ],
   alphaCSR[ 253 ][ 366 ],
   alphaCSR[ 253 ][ 367 ],
   alphaCSR[ 253 ][ 368 ],
   alphaCSR[ 253 ][ 369 ],
   alphaCSR[ 253 ][ 370 ],
   alphaCSR[ 253 ][ 371 ],
   alphaCSR[ 253 ][ 372 ],
   alphaCSR[ 253 ][ 373 ],
   alphaCSR[ 253 ][ 374 ],
   alphaCSR[ 253 ][ 375 ],
   alphaCSR[ 253 ][ 376 ],
   alphaCSR[ 253 ][ 377 ],
   alphaCSR[ 253 ][ 378 ],
   alphaCSR[ 253 ][ 379 ],
   alphaCSR[ 253 ][ 380 ],
   alphaCSR[ 253 ][ 381 ],
   alphaCSR[ 253 ][ 382 ],
   alphaCSR[ 253 ][ 383 ],
   alphaCSR[ 254 ][ 0 ],
   alphaCSR[ 254 ][ 1 ],
   alphaCSR[ 254 ][ 2 ],
   alphaCSR[ 254 ][ 3 ],
   alphaCSR[ 254 ][ 4 ],
   alphaCSR[ 254 ][ 5 ],
   alphaCSR[ 254 ][ 6 ],
   alphaCSR[ 254 ][ 7 ],
   alphaCSR[ 254 ][ 8 ],
   alphaCSR[ 254 ][ 9 ],
   alphaCSR[ 254 ][ 10 ],
   alphaCSR[ 254 ][ 11 ],
   alphaCSR[ 254 ][ 12 ],
   alphaCSR[ 254 ][ 13 ],
   alphaCSR[ 254 ][ 14 ],
   alphaCSR[ 254 ][ 15 ],
   alphaCSR[ 254 ][ 16 ],
   alphaCSR[ 254 ][ 17 ],
   alphaCSR[ 254 ][ 18 ],
   alphaCSR[ 254 ][ 19 ],
   alphaCSR[ 254 ][ 20 ],
   alphaCSR[ 254 ][ 21 ],
   alphaCSR[ 254 ][ 22 ],
   alphaCSR[ 254 ][ 23 ],
   alphaCSR[ 254 ][ 24 ],
   alphaCSR[ 254 ][ 25 ],
   alphaCSR[ 254 ][ 26 ],
   alphaCSR[ 254 ][ 27 ],
   alphaCSR[ 254 ][ 28 ],
   alphaCSR[ 254 ][ 29 ],
   alphaCSR[ 254 ][ 30 ],
   alphaCSR[ 254 ][ 31 ],
   alphaCSR[ 254 ][ 32 ],
   alphaCSR[ 254 ][ 33 ],
   alphaCSR[ 254 ][ 34 ],
   alphaCSR[ 254 ][ 35 ],
   alphaCSR[ 254 ][ 36 ],
   alphaCSR[ 254 ][ 37 ],
   alphaCSR[ 254 ][ 38 ],
   alphaCSR[ 254 ][ 39 ],
   alphaCSR[ 254 ][ 40 ],
   alphaCSR[ 254 ][ 41 ],
   alphaCSR[ 254 ][ 42 ],
   alphaCSR[ 254 ][ 43 ],
   alphaCSR[ 254 ][ 44 ],
   alphaCSR[ 254 ][ 45 ],
   alphaCSR[ 254 ][ 46 ],
   alphaCSR[ 254 ][ 47 ],
   alphaCSR[ 254 ][ 48 ],
   alphaCSR[ 254 ][ 49 ],
   alphaCSR[ 254 ][ 50 ],
   alphaCSR[ 254 ][ 51 ],
   alphaCSR[ 254 ][ 52 ],
   alphaCSR[ 254 ][ 53 ],
   alphaCSR[ 254 ][ 54 ],
   alphaCSR[ 254 ][ 55 ],
   alphaCSR[ 254 ][ 56 ],
   alphaCSR[ 254 ][ 57 ],
   alphaCSR[ 254 ][ 58 ],
   alphaCSR[ 254 ][ 59 ],
   alphaCSR[ 254 ][ 60 ],
   alphaCSR[ 254 ][ 61 ],
   alphaCSR[ 254 ][ 62 ],
   alphaCSR[ 254 ][ 63 ],
   alphaCSR[ 254 ][ 64 ],
   alphaCSR[ 254 ][ 65 ],
   alphaCSR[ 254 ][ 66 ],
   alphaCSR[ 254 ][ 67 ],
   alphaCSR[ 254 ][ 68 ],
   alphaCSR[ 254 ][ 69 ],
   alphaCSR[ 254 ][ 70 ],
   alphaCSR[ 254 ][ 71 ],
   alphaCSR[ 254 ][ 72 ],
   alphaCSR[ 254 ][ 73 ],
   alphaCSR[ 254 ][ 74 ],
   alphaCSR[ 254 ][ 75 ],
   alphaCSR[ 254 ][ 76 ],
   alphaCSR[ 254 ][ 77 ],
   alphaCSR[ 254 ][ 78 ],
   alphaCSR[ 254 ][ 79 ],
   alphaCSR[ 254 ][ 80 ],
   alphaCSR[ 254 ][ 81 ],
   alphaCSR[ 254 ][ 82 ],
   alphaCSR[ 254 ][ 83 ],
   alphaCSR[ 254 ][ 84 ],
   alphaCSR[ 254 ][ 85 ],
   alphaCSR[ 254 ][ 86 ],
   alphaCSR[ 254 ][ 87 ],
   alphaCSR[ 254 ][ 88 ],
   alphaCSR[ 254 ][ 89 ],
   alphaCSR[ 254 ][ 90 ],
   alphaCSR[ 254 ][ 91 ],
   alphaCSR[ 254 ][ 92 ],
   alphaCSR[ 254 ][ 93 ],
   alphaCSR[ 254 ][ 94 ],
   alphaCSR[ 254 ][ 95 ],
   alphaCSR[ 254 ][ 96 ],
   alphaCSR[ 254 ][ 97 ],
   alphaCSR[ 254 ][ 98 ],
   alphaCSR[ 254 ][ 99 ],
   alphaCSR[ 254 ][ 100 ],
   alphaCSR[ 254 ][ 101 ],
   alphaCSR[ 254 ][ 102 ],
   alphaCSR[ 254 ][ 103 ],
   alphaCSR[ 254 ][ 104 ],
   alphaCSR[ 254 ][ 105 ],
   alphaCSR[ 254 ][ 106 ],
   alphaCSR[ 254 ][ 107 ],
   alphaCSR[ 254 ][ 108 ],
   alphaCSR[ 254 ][ 109 ],
   alphaCSR[ 254 ][ 110 ],
   alphaCSR[ 254 ][ 111 ],
   alphaCSR[ 254 ][ 112 ],
   alphaCSR[ 254 ][ 113 ],
   alphaCSR[ 254 ][ 114 ],
   alphaCSR[ 254 ][ 115 ],
   alphaCSR[ 254 ][ 116 ],
   alphaCSR[ 254 ][ 117 ],
   alphaCSR[ 254 ][ 118 ],
   alphaCSR[ 254 ][ 119 ],
   alphaCSR[ 254 ][ 120 ],
   alphaCSR[ 254 ][ 121 ],
   alphaCSR[ 254 ][ 122 ],
   alphaCSR[ 254 ][ 123 ],
   alphaCSR[ 254 ][ 124 ],
   alphaCSR[ 254 ][ 125 ],
   alphaCSR[ 254 ][ 126 ],
   alphaCSR[ 254 ][ 127 ],
   alphaCSR[ 254 ][ 128 ],
   alphaCSR[ 254 ][ 129 ],
   alphaCSR[ 254 ][ 130 ],
   alphaCSR[ 254 ][ 131 ],
   alphaCSR[ 254 ][ 132 ],
   alphaCSR[ 254 ][ 133 ],
   alphaCSR[ 254 ][ 134 ],
   alphaCSR[ 254 ][ 135 ],
   alphaCSR[ 254 ][ 136 ],
   alphaCSR[ 254 ][ 137 ],
   alphaCSR[ 254 ][ 138 ],
   alphaCSR[ 254 ][ 139 ],
   alphaCSR[ 254 ][ 140 ],
   alphaCSR[ 254 ][ 141 ],
   alphaCSR[ 254 ][ 142 ],
   alphaCSR[ 254 ][ 143 ],
   alphaCSR[ 254 ][ 144 ],
   alphaCSR[ 254 ][ 145 ],
   alphaCSR[ 254 ][ 146 ],
   alphaCSR[ 254 ][ 147 ],
   alphaCSR[ 254 ][ 148 ],
   alphaCSR[ 254 ][ 149 ],
   alphaCSR[ 254 ][ 150 ],
   alphaCSR[ 254 ][ 151 ],
   alphaCSR[ 254 ][ 152 ],
   alphaCSR[ 254 ][ 153 ],
   alphaCSR[ 254 ][ 154 ],
   alphaCSR[ 254 ][ 155 ],
   alphaCSR[ 254 ][ 156 ],
   alphaCSR[ 254 ][ 157 ],
   alphaCSR[ 254 ][ 158 ],
   alphaCSR[ 254 ][ 159 ],
   alphaCSR[ 254 ][ 160 ],
   alphaCSR[ 254 ][ 161 ],
   alphaCSR[ 254 ][ 162 ],
   alphaCSR[ 254 ][ 163 ],
   alphaCSR[ 254 ][ 164 ],
   alphaCSR[ 254 ][ 165 ],
   alphaCSR[ 254 ][ 166 ],
   alphaCSR[ 254 ][ 167 ],
   alphaCSR[ 254 ][ 168 ],
   alphaCSR[ 254 ][ 169 ],
   alphaCSR[ 254 ][ 170 ],
   alphaCSR[ 254 ][ 171 ],
   alphaCSR[ 254 ][ 172 ],
   alphaCSR[ 254 ][ 173 ],
   alphaCSR[ 254 ][ 174 ],
   alphaCSR[ 254 ][ 175 ],
   alphaCSR[ 254 ][ 176 ],
   alphaCSR[ 254 ][ 177 ],
   alphaCSR[ 254 ][ 178 ],
   alphaCSR[ 254 ][ 179 ],
   alphaCSR[ 254 ][ 180 ],
   alphaCSR[ 254 ][ 181 ],
   alphaCSR[ 254 ][ 182 ],
   alphaCSR[ 254 ][ 183 ],
   alphaCSR[ 254 ][ 184 ],
   alphaCSR[ 254 ][ 185 ],
   alphaCSR[ 254 ][ 186 ],
   alphaCSR[ 254 ][ 187 ],
   alphaCSR[ 254 ][ 188 ],
   alphaCSR[ 254 ][ 189 ],
   alphaCSR[ 254 ][ 190 ],
   alphaCSR[ 254 ][ 191 ],
   alphaCSR[ 254 ][ 192 ],
   alphaCSR[ 254 ][ 193 ],
   alphaCSR[ 254 ][ 194 ],
   alphaCSR[ 254 ][ 195 ],
   alphaCSR[ 254 ][ 196 ],
   alphaCSR[ 254 ][ 197 ],
   alphaCSR[ 254 ][ 198 ],
   alphaCSR[ 254 ][ 199 ],
   alphaCSR[ 254 ][ 200 ],
   alphaCSR[ 254 ][ 201 ],
   alphaCSR[ 254 ][ 202 ],
   alphaCSR[ 254 ][ 203 ],
   alphaCSR[ 254 ][ 204 ],
   alphaCSR[ 254 ][ 205 ],
   alphaCSR[ 254 ][ 206 ],
   alphaCSR[ 254 ][ 207 ],
   alphaCSR[ 254 ][ 208 ],
   alphaCSR[ 254 ][ 209 ],
   alphaCSR[ 254 ][ 210 ],
   alphaCSR[ 254 ][ 211 ],
   alphaCSR[ 254 ][ 212 ],
   alphaCSR[ 254 ][ 213 ],
   alphaCSR[ 254 ][ 214 ],
   alphaCSR[ 254 ][ 215 ],
   alphaCSR[ 254 ][ 216 ],
   alphaCSR[ 254 ][ 217 ],
   alphaCSR[ 254 ][ 218 ],
   alphaCSR[ 254 ][ 219 ],
   alphaCSR[ 254 ][ 220 ],
   alphaCSR[ 254 ][ 221 ],
   alphaCSR[ 254 ][ 222 ],
   alphaCSR[ 254 ][ 223 ],
   alphaCSR[ 254 ][ 224 ],
   alphaCSR[ 254 ][ 225 ],
   alphaCSR[ 254 ][ 226 ],
   alphaCSR[ 254 ][ 227 ],
   alphaCSR[ 254 ][ 228 ],
   alphaCSR[ 254 ][ 229 ],
   alphaCSR[ 254 ][ 230 ],
   alphaCSR[ 254 ][ 231 ],
   alphaCSR[ 254 ][ 232 ],
   alphaCSR[ 254 ][ 233 ],
   alphaCSR[ 254 ][ 234 ],
   alphaCSR[ 254 ][ 235 ],
   alphaCSR[ 254 ][ 236 ],
   alphaCSR[ 254 ][ 237 ],
   alphaCSR[ 254 ][ 238 ],
   alphaCSR[ 254 ][ 239 ],
   alphaCSR[ 254 ][ 240 ],
   alphaCSR[ 254 ][ 241 ],
   alphaCSR[ 254 ][ 242 ],
   alphaCSR[ 254 ][ 243 ],
   alphaCSR[ 254 ][ 244 ],
   alphaCSR[ 254 ][ 245 ],
   alphaCSR[ 254 ][ 246 ],
   alphaCSR[ 254 ][ 247 ],
   alphaCSR[ 254 ][ 248 ],
   alphaCSR[ 254 ][ 249 ],
   alphaCSR[ 254 ][ 250 ],
   alphaCSR[ 254 ][ 251 ],
   alphaCSR[ 254 ][ 252 ],
   alphaCSR[ 254 ][ 253 ],
   alphaCSR[ 254 ][ 254 ],
   alphaCSR[ 254 ][ 255 ],
   alphaCSR[ 254 ][ 256 ],
   alphaCSR[ 254 ][ 257 ],
   alphaCSR[ 254 ][ 258 ],
   alphaCSR[ 254 ][ 259 ],
   alphaCSR[ 254 ][ 260 ],
   alphaCSR[ 254 ][ 261 ],
   alphaCSR[ 254 ][ 262 ],
   alphaCSR[ 254 ][ 263 ],
   alphaCSR[ 254 ][ 264 ],
   alphaCSR[ 254 ][ 265 ],
   alphaCSR[ 254 ][ 266 ],
   alphaCSR[ 254 ][ 267 ],
   alphaCSR[ 254 ][ 268 ],
   alphaCSR[ 254 ][ 269 ],
   alphaCSR[ 254 ][ 270 ],
   alphaCSR[ 254 ][ 271 ],
   alphaCSR[ 254 ][ 272 ],
   alphaCSR[ 254 ][ 273 ],
   alphaCSR[ 254 ][ 274 ],
   alphaCSR[ 254 ][ 275 ],
   alphaCSR[ 254 ][ 276 ],
   alphaCSR[ 254 ][ 277 ],
   alphaCSR[ 254 ][ 278 ],
   alphaCSR[ 254 ][ 279 ],
   alphaCSR[ 254 ][ 280 ],
   alphaCSR[ 254 ][ 281 ],
   alphaCSR[ 254 ][ 282 ],
   alphaCSR[ 254 ][ 283 ],
   alphaCSR[ 254 ][ 284 ],
   alphaCSR[ 254 ][ 285 ],
   alphaCSR[ 254 ][ 286 ],
   alphaCSR[ 254 ][ 287 ],
   alphaCSR[ 254 ][ 288 ],
   alphaCSR[ 254 ][ 289 ],
   alphaCSR[ 254 ][ 290 ],
   alphaCSR[ 254 ][ 291 ],
   alphaCSR[ 254 ][ 292 ],
   alphaCSR[ 254 ][ 293 ],
   alphaCSR[ 254 ][ 294 ],
   alphaCSR[ 254 ][ 295 ],
   alphaCSR[ 254 ][ 296 ],
   alphaCSR[ 254 ][ 297 ],
   alphaCSR[ 254 ][ 298 ],
   alphaCSR[ 254 ][ 299 ],
   alphaCSR[ 254 ][ 300 ],
   alphaCSR[ 254 ][ 301 ],
   alphaCSR[ 254 ][ 302 ],
   alphaCSR[ 254 ][ 303 ],
   alphaCSR[ 254 ][ 304 ],
   alphaCSR[ 254 ][ 305 ],
   alphaCSR[ 254 ][ 306 ],
   alphaCSR[ 254 ][ 307 ],
   alphaCSR[ 254 ][ 308 ],
   alphaCSR[ 254 ][ 309 ],
   alphaCSR[ 254 ][ 310 ],
   alphaCSR[ 254 ][ 311 ],
   alphaCSR[ 254 ][ 312 ],
   alphaCSR[ 254 ][ 313 ],
   alphaCSR[ 254 ][ 314 ],
   alphaCSR[ 254 ][ 315 ],
   alphaCSR[ 254 ][ 316 ],
   alphaCSR[ 254 ][ 317 ],
   alphaCSR[ 254 ][ 318 ],
   alphaCSR[ 254 ][ 319 ],
   alphaCSR[ 254 ][ 320 ],
   alphaCSR[ 254 ][ 321 ],
   alphaCSR[ 254 ][ 322 ],
   alphaCSR[ 254 ][ 323 ],
   alphaCSR[ 254 ][ 324 ],
   alphaCSR[ 254 ][ 325 ],
   alphaCSR[ 254 ][ 326 ],
   alphaCSR[ 254 ][ 327 ],
   alphaCSR[ 254 ][ 328 ],
   alphaCSR[ 254 ][ 329 ],
   alphaCSR[ 254 ][ 330 ],
   alphaCSR[ 254 ][ 331 ],
   alphaCSR[ 254 ][ 332 ],
   alphaCSR[ 254 ][ 333 ],
   alphaCSR[ 254 ][ 334 ],
   alphaCSR[ 254 ][ 335 ],
   alphaCSR[ 254 ][ 336 ],
   alphaCSR[ 254 ][ 337 ],
   alphaCSR[ 254 ][ 338 ],
   alphaCSR[ 254 ][ 339 ],
   alphaCSR[ 254 ][ 340 ],
   alphaCSR[ 254 ][ 341 ],
   alphaCSR[ 254 ][ 342 ],
   alphaCSR[ 254 ][ 343 ],
   alphaCSR[ 254 ][ 344 ],
   alphaCSR[ 254 ][ 345 ],
   alphaCSR[ 254 ][ 346 ],
   alphaCSR[ 254 ][ 347 ],
   alphaCSR[ 254 ][ 348 ],
   alphaCSR[ 254 ][ 349 ],
   alphaCSR[ 254 ][ 350 ],
   alphaCSR[ 254 ][ 351 ],
   alphaCSR[ 254 ][ 352 ],
   alphaCSR[ 254 ][ 353 ],
   alphaCSR[ 254 ][ 354 ],
   alphaCSR[ 254 ][ 355 ],
   alphaCSR[ 254 ][ 356 ],
   alphaCSR[ 254 ][ 357 ],
   alphaCSR[ 254 ][ 358 ],
   alphaCSR[ 254 ][ 359 ],
   alphaCSR[ 254 ][ 360 ],
   alphaCSR[ 254 ][ 361 ],
   alphaCSR[ 254 ][ 362 ],
   alphaCSR[ 254 ][ 363 ],
   alphaCSR[ 254 ][ 364 ],
   alphaCSR[ 254 ][ 365 ],
   alphaCSR[ 254 ][ 366 ],
   alphaCSR[ 254 ][ 367 ],
   alphaCSR[ 254 ][ 368 ],
   alphaCSR[ 254 ][ 369 ],
   alphaCSR[ 254 ][ 370 ],
   alphaCSR[ 254 ][ 371 ],
   alphaCSR[ 254 ][ 372 ],
   alphaCSR[ 254 ][ 373 ],
   alphaCSR[ 254 ][ 374 ],
   alphaCSR[ 254 ][ 375 ],
   alphaCSR[ 254 ][ 376 ],
   alphaCSR[ 254 ][ 377 ],
   alphaCSR[ 254 ][ 378 ],
   alphaCSR[ 254 ][ 379 ],
   alphaCSR[ 254 ][ 380 ],
   alphaCSR[ 254 ][ 381 ],
   alphaCSR[ 254 ][ 382 ],
   alphaCSR[ 254 ][ 383 ],
   alphaCSR[ 255 ][ 0 ],
   alphaCSR[ 255 ][ 1 ],
   alphaCSR[ 255 ][ 2 ],
   alphaCSR[ 255 ][ 3 ],
   alphaCSR[ 255 ][ 4 ],
   alphaCSR[ 255 ][ 5 ],
   alphaCSR[ 255 ][ 6 ],
   alphaCSR[ 255 ][ 7 ],
   alphaCSR[ 255 ][ 8 ],
   alphaCSR[ 255 ][ 9 ],
   alphaCSR[ 255 ][ 10 ],
   alphaCSR[ 255 ][ 11 ],
   alphaCSR[ 255 ][ 12 ],
   alphaCSR[ 255 ][ 13 ],
   alphaCSR[ 255 ][ 14 ],
   alphaCSR[ 255 ][ 15 ],
   alphaCSR[ 255 ][ 16 ],
   alphaCSR[ 255 ][ 17 ],
   alphaCSR[ 255 ][ 18 ],
   alphaCSR[ 255 ][ 19 ],
   alphaCSR[ 255 ][ 20 ],
   alphaCSR[ 255 ][ 21 ],
   alphaCSR[ 255 ][ 22 ],
   alphaCSR[ 255 ][ 23 ],
   alphaCSR[ 255 ][ 24 ],
   alphaCSR[ 255 ][ 25 ],
   alphaCSR[ 255 ][ 26 ],
   alphaCSR[ 255 ][ 27 ],
   alphaCSR[ 255 ][ 28 ],
   alphaCSR[ 255 ][ 29 ],
   alphaCSR[ 255 ][ 30 ],
   alphaCSR[ 255 ][ 31 ],
   alphaCSR[ 255 ][ 32 ],
   alphaCSR[ 255 ][ 33 ],
   alphaCSR[ 255 ][ 34 ],
   alphaCSR[ 255 ][ 35 ],
   alphaCSR[ 255 ][ 36 ],
   alphaCSR[ 255 ][ 37 ],
   alphaCSR[ 255 ][ 38 ],
   alphaCSR[ 255 ][ 39 ],
   alphaCSR[ 255 ][ 40 ],
   alphaCSR[ 255 ][ 41 ],
   alphaCSR[ 255 ][ 42 ],
   alphaCSR[ 255 ][ 43 ],
   alphaCSR[ 255 ][ 44 ],
   alphaCSR[ 255 ][ 45 ],
   alphaCSR[ 255 ][ 46 ],
   alphaCSR[ 255 ][ 47 ],
   alphaCSR[ 255 ][ 48 ],
   alphaCSR[ 255 ][ 49 ],
   alphaCSR[ 255 ][ 50 ],
   alphaCSR[ 255 ][ 51 ],
   alphaCSR[ 255 ][ 52 ],
   alphaCSR[ 255 ][ 53 ],
   alphaCSR[ 255 ][ 54 ],
   alphaCSR[ 255 ][ 55 ],
   alphaCSR[ 255 ][ 56 ],
   alphaCSR[ 255 ][ 57 ],
   alphaCSR[ 255 ][ 58 ],
   alphaCSR[ 255 ][ 59 ],
   alphaCSR[ 255 ][ 60 ],
   alphaCSR[ 255 ][ 61 ],
   alphaCSR[ 255 ][ 62 ],
   alphaCSR[ 255 ][ 63 ],
   alphaCSR[ 255 ][ 64 ],
   alphaCSR[ 255 ][ 65 ],
   alphaCSR[ 255 ][ 66 ],
   alphaCSR[ 255 ][ 67 ],
   alphaCSR[ 255 ][ 68 ],
   alphaCSR[ 255 ][ 69 ],
   alphaCSR[ 255 ][ 70 ],
   alphaCSR[ 255 ][ 71 ],
   alphaCSR[ 255 ][ 72 ],
   alphaCSR[ 255 ][ 73 ],
   alphaCSR[ 255 ][ 74 ],
   alphaCSR[ 255 ][ 75 ],
   alphaCSR[ 255 ][ 76 ],
   alphaCSR[ 255 ][ 77 ],
   alphaCSR[ 255 ][ 78 ],
   alphaCSR[ 255 ][ 79 ],
   alphaCSR[ 255 ][ 80 ],
   alphaCSR[ 255 ][ 81 ],
   alphaCSR[ 255 ][ 82 ],
   alphaCSR[ 255 ][ 83 ],
   alphaCSR[ 255 ][ 84 ],
   alphaCSR[ 255 ][ 85 ],
   alphaCSR[ 255 ][ 86 ],
   alphaCSR[ 255 ][ 87 ],
   alphaCSR[ 255 ][ 88 ],
   alphaCSR[ 255 ][ 89 ],
   alphaCSR[ 255 ][ 90 ],
   alphaCSR[ 255 ][ 91 ],
   alphaCSR[ 255 ][ 92 ],
   alphaCSR[ 255 ][ 93 ],
   alphaCSR[ 255 ][ 94 ],
   alphaCSR[ 255 ][ 95 ],
   alphaCSR[ 255 ][ 96 ],
   alphaCSR[ 255 ][ 97 ],
   alphaCSR[ 255 ][ 98 ],
   alphaCSR[ 255 ][ 99 ],
   alphaCSR[ 255 ][ 100 ],
   alphaCSR[ 255 ][ 101 ],
   alphaCSR[ 255 ][ 102 ],
   alphaCSR[ 255 ][ 103 ],
   alphaCSR[ 255 ][ 104 ],
   alphaCSR[ 255 ][ 105 ],
   alphaCSR[ 255 ][ 106 ],
   alphaCSR[ 255 ][ 107 ],
   alphaCSR[ 255 ][ 108 ],
   alphaCSR[ 255 ][ 109 ],
   alphaCSR[ 255 ][ 110 ],
   alphaCSR[ 255 ][ 111 ],
   alphaCSR[ 255 ][ 112 ],
   alphaCSR[ 255 ][ 113 ],
   alphaCSR[ 255 ][ 114 ],
   alphaCSR[ 255 ][ 115 ],
   alphaCSR[ 255 ][ 116 ],
   alphaCSR[ 255 ][ 117 ],
   alphaCSR[ 255 ][ 118 ],
   alphaCSR[ 255 ][ 119 ],
   alphaCSR[ 255 ][ 120 ],
   alphaCSR[ 255 ][ 121 ],
   alphaCSR[ 255 ][ 122 ],
   alphaCSR[ 255 ][ 123 ],
   alphaCSR[ 255 ][ 124 ],
   alphaCSR[ 255 ][ 125 ],
   alphaCSR[ 255 ][ 126 ],
   alphaCSR[ 255 ][ 127 ],
   alphaCSR[ 255 ][ 128 ],
   alphaCSR[ 255 ][ 129 ],
   alphaCSR[ 255 ][ 130 ],
   alphaCSR[ 255 ][ 131 ],
   alphaCSR[ 255 ][ 132 ],
   alphaCSR[ 255 ][ 133 ],
   alphaCSR[ 255 ][ 134 ],
   alphaCSR[ 255 ][ 135 ],
   alphaCSR[ 255 ][ 136 ],
   alphaCSR[ 255 ][ 137 ],
   alphaCSR[ 255 ][ 138 ],
   alphaCSR[ 255 ][ 139 ],
   alphaCSR[ 255 ][ 140 ],
   alphaCSR[ 255 ][ 141 ],
   alphaCSR[ 255 ][ 142 ],
   alphaCSR[ 255 ][ 143 ],
   alphaCSR[ 255 ][ 144 ],
   alphaCSR[ 255 ][ 145 ],
   alphaCSR[ 255 ][ 146 ],
   alphaCSR[ 255 ][ 147 ],
   alphaCSR[ 255 ][ 148 ],
   alphaCSR[ 255 ][ 149 ],
   alphaCSR[ 255 ][ 150 ],
   alphaCSR[ 255 ][ 151 ],
   alphaCSR[ 255 ][ 152 ],
   alphaCSR[ 255 ][ 153 ],
   alphaCSR[ 255 ][ 154 ],
   alphaCSR[ 255 ][ 155 ],
   alphaCSR[ 255 ][ 156 ],
   alphaCSR[ 255 ][ 157 ],
   alphaCSR[ 255 ][ 158 ],
   alphaCSR[ 255 ][ 159 ],
   alphaCSR[ 255 ][ 160 ],
   alphaCSR[ 255 ][ 161 ],
   alphaCSR[ 255 ][ 162 ],
   alphaCSR[ 255 ][ 163 ],
   alphaCSR[ 255 ][ 164 ],
   alphaCSR[ 255 ][ 165 ],
   alphaCSR[ 255 ][ 166 ],
   alphaCSR[ 255 ][ 167 ],
   alphaCSR[ 255 ][ 168 ],
   alphaCSR[ 255 ][ 169 ],
   alphaCSR[ 255 ][ 170 ],
   alphaCSR[ 255 ][ 171 ],
   alphaCSR[ 255 ][ 172 ],
   alphaCSR[ 255 ][ 173 ],
   alphaCSR[ 255 ][ 174 ],
   alphaCSR[ 255 ][ 175 ],
   alphaCSR[ 255 ][ 176 ],
   alphaCSR[ 255 ][ 177 ],
   alphaCSR[ 255 ][ 178 ],
   alphaCSR[ 255 ][ 179 ],
   alphaCSR[ 255 ][ 180 ],
   alphaCSR[ 255 ][ 181 ],
   alphaCSR[ 255 ][ 182 ],
   alphaCSR[ 255 ][ 183 ],
   alphaCSR[ 255 ][ 184 ],
   alphaCSR[ 255 ][ 185 ],
   alphaCSR[ 255 ][ 186 ],
   alphaCSR[ 255 ][ 187 ],
   alphaCSR[ 255 ][ 188 ],
   alphaCSR[ 255 ][ 189 ],
   alphaCSR[ 255 ][ 190 ],
   alphaCSR[ 255 ][ 191 ],
   alphaCSR[ 255 ][ 192 ],
   alphaCSR[ 255 ][ 193 ],
   alphaCSR[ 255 ][ 194 ],
   alphaCSR[ 255 ][ 195 ],
   alphaCSR[ 255 ][ 196 ],
   alphaCSR[ 255 ][ 197 ],
   alphaCSR[ 255 ][ 198 ],
   alphaCSR[ 255 ][ 199 ],
   alphaCSR[ 255 ][ 200 ],
   alphaCSR[ 255 ][ 201 ],
   alphaCSR[ 255 ][ 202 ],
   alphaCSR[ 255 ][ 203 ],
   alphaCSR[ 255 ][ 204 ],
   alphaCSR[ 255 ][ 205 ],
   alphaCSR[ 255 ][ 206 ],
   alphaCSR[ 255 ][ 207 ],
   alphaCSR[ 255 ][ 208 ],
   alphaCSR[ 255 ][ 209 ],
   alphaCSR[ 255 ][ 210 ],
   alphaCSR[ 255 ][ 211 ],
   alphaCSR[ 255 ][ 212 ],
   alphaCSR[ 255 ][ 213 ],
   alphaCSR[ 255 ][ 214 ],
   alphaCSR[ 255 ][ 215 ],
   alphaCSR[ 255 ][ 216 ],
   alphaCSR[ 255 ][ 217 ],
   alphaCSR[ 255 ][ 218 ],
   alphaCSR[ 255 ][ 219 ],
   alphaCSR[ 255 ][ 220 ],
   alphaCSR[ 255 ][ 221 ],
   alphaCSR[ 255 ][ 222 ],
   alphaCSR[ 255 ][ 223 ],
   alphaCSR[ 255 ][ 224 ],
   alphaCSR[ 255 ][ 225 ],
   alphaCSR[ 255 ][ 226 ],
   alphaCSR[ 255 ][ 227 ],
   alphaCSR[ 255 ][ 228 ],
   alphaCSR[ 255 ][ 229 ],
   alphaCSR[ 255 ][ 230 ],
   alphaCSR[ 255 ][ 231 ],
   alphaCSR[ 255 ][ 232 ],
   alphaCSR[ 255 ][ 233 ],
   alphaCSR[ 255 ][ 234 ],
   alphaCSR[ 255 ][ 235 ],
   alphaCSR[ 255 ][ 236 ],
   alphaCSR[ 255 ][ 237 ],
   alphaCSR[ 255 ][ 238 ],
   alphaCSR[ 255 ][ 239 ],
   alphaCSR[ 255 ][ 240 ],
   alphaCSR[ 255 ][ 241 ],
   alphaCSR[ 255 ][ 242 ],
   alphaCSR[ 255 ][ 243 ],
   alphaCSR[ 255 ][ 244 ],
   alphaCSR[ 255 ][ 245 ],
   alphaCSR[ 255 ][ 246 ],
   alphaCSR[ 255 ][ 247 ],
   alphaCSR[ 255 ][ 248 ],
   alphaCSR[ 255 ][ 249 ],
   alphaCSR[ 255 ][ 250 ],
   alphaCSR[ 255 ][ 251 ],
   alphaCSR[ 255 ][ 252 ],
   alphaCSR[ 255 ][ 253 ],
   alphaCSR[ 255 ][ 254 ],
   alphaCSR[ 255 ][ 255 ],
   alphaCSR[ 255 ][ 256 ],
   alphaCSR[ 255 ][ 257 ],
   alphaCSR[ 255 ][ 258 ],
   alphaCSR[ 255 ][ 259 ],
   alphaCSR[ 255 ][ 260 ],
   alphaCSR[ 255 ][ 261 ],
   alphaCSR[ 255 ][ 262 ],
   alphaCSR[ 255 ][ 263 ],
   alphaCSR[ 255 ][ 264 ],
   alphaCSR[ 255 ][ 265 ],
   alphaCSR[ 255 ][ 266 ],
   alphaCSR[ 255 ][ 267 ],
   alphaCSR[ 255 ][ 268 ],
   alphaCSR[ 255 ][ 269 ],
   alphaCSR[ 255 ][ 270 ],
   alphaCSR[ 255 ][ 271 ],
   alphaCSR[ 255 ][ 272 ],
   alphaCSR[ 255 ][ 273 ],
   alphaCSR[ 255 ][ 274 ],
   alphaCSR[ 255 ][ 275 ],
   alphaCSR[ 255 ][ 276 ],
   alphaCSR[ 255 ][ 277 ],
   alphaCSR[ 255 ][ 278 ],
   alphaCSR[ 255 ][ 279 ],
   alphaCSR[ 255 ][ 280 ],
   alphaCSR[ 255 ][ 281 ],
   alphaCSR[ 255 ][ 282 ],
   alphaCSR[ 255 ][ 283 ],
   alphaCSR[ 255 ][ 284 ],
   alphaCSR[ 255 ][ 285 ],
   alphaCSR[ 255 ][ 286 ],
   alphaCSR[ 255 ][ 287 ],
   alphaCSR[ 255 ][ 288 ],
   alphaCSR[ 255 ][ 289 ],
   alphaCSR[ 255 ][ 290 ],
   alphaCSR[ 255 ][ 291 ],
   alphaCSR[ 255 ][ 292 ],
   alphaCSR[ 255 ][ 293 ],
   alphaCSR[ 255 ][ 294 ],
   alphaCSR[ 255 ][ 295 ],
   alphaCSR[ 255 ][ 296 ],
   alphaCSR[ 255 ][ 297 ],
   alphaCSR[ 255 ][ 298 ],
   alphaCSR[ 255 ][ 299 ],
   alphaCSR[ 255 ][ 300 ],
   alphaCSR[ 255 ][ 301 ],
   alphaCSR[ 255 ][ 302 ],
   alphaCSR[ 255 ][ 303 ],
   alphaCSR[ 255 ][ 304 ],
   alphaCSR[ 255 ][ 305 ],
   alphaCSR[ 255 ][ 306 ],
   alphaCSR[ 255 ][ 307 ],
   alphaCSR[ 255 ][ 308 ],
   alphaCSR[ 255 ][ 309 ],
   alphaCSR[ 255 ][ 310 ],
   alphaCSR[ 255 ][ 311 ],
   alphaCSR[ 255 ][ 312 ],
   alphaCSR[ 255 ][ 313 ],
   alphaCSR[ 255 ][ 314 ],
   alphaCSR[ 255 ][ 315 ],
   alphaCSR[ 255 ][ 316 ],
   alphaCSR[ 255 ][ 317 ],
   alphaCSR[ 255 ][ 318 ],
   alphaCSR[ 255 ][ 319 ],
   alphaCSR[ 255 ][ 320 ],
   alphaCSR[ 255 ][ 321 ],
   alphaCSR[ 255 ][ 322 ],
   alphaCSR[ 255 ][ 323 ],
   alphaCSR[ 255 ][ 324 ],
   alphaCSR[ 255 ][ 325 ],
   alphaCSR[ 255 ][ 326 ],
   alphaCSR[ 255 ][ 327 ],
   alphaCSR[ 255 ][ 328 ],
   alphaCSR[ 255 ][ 329 ],
   alphaCSR[ 255 ][ 330 ],
   alphaCSR[ 255 ][ 331 ],
   alphaCSR[ 255 ][ 332 ],
   alphaCSR[ 255 ][ 333 ],
   alphaCSR[ 255 ][ 334 ],
   alphaCSR[ 255 ][ 335 ],
   alphaCSR[ 255 ][ 336 ],
   alphaCSR[ 255 ][ 337 ],
   alphaCSR[ 255 ][ 338 ],
   alphaCSR[ 255 ][ 339 ],
   alphaCSR[ 255 ][ 340 ],
   alphaCSR[ 255 ][ 341 ],
   alphaCSR[ 255 ][ 342 ],
   alphaCSR[ 255 ][ 343 ],
   alphaCSR[ 255 ][ 344 ],
   alphaCSR[ 255 ][ 345 ],
   alphaCSR[ 255 ][ 346 ],
   alphaCSR[ 255 ][ 347 ],
   alphaCSR[ 255 ][ 348 ],
   alphaCSR[ 255 ][ 349 ],
   alphaCSR[ 255 ][ 350 ],
   alphaCSR[ 255 ][ 351 ],
   alphaCSR[ 255 ][ 352 ],
   alphaCSR[ 255 ][ 353 ],
   alphaCSR[ 255 ][ 354 ],
   alphaCSR[ 255 ][ 355 ],
   alphaCSR[ 255 ][ 356 ],
   alphaCSR[ 255 ][ 357 ],
   alphaCSR[ 255 ][ 358 ],
   alphaCSR[ 255 ][ 359 ],
   alphaCSR[ 255 ][ 360 ],
   alphaCSR[ 255 ][ 361 ],
   alphaCSR[ 255 ][ 362 ],
   alphaCSR[ 255 ][ 363 ],
   alphaCSR[ 255 ][ 364 ],
   alphaCSR[ 255 ][ 365 ],
   alphaCSR[ 255 ][ 366 ],
   alphaCSR[ 255 ][ 367 ],
   alphaCSR[ 255 ][ 368 ],
   alphaCSR[ 255 ][ 369 ],
   alphaCSR[ 255 ][ 370 ],
   alphaCSR[ 255 ][ 371 ],
   alphaCSR[ 255 ][ 372 ],
   alphaCSR[ 255 ][ 373 ],
   alphaCSR[ 255 ][ 374 ],
   alphaCSR[ 255 ][ 375 ],
   alphaCSR[ 255 ][ 376 ],
   alphaCSR[ 255 ][ 377 ],
   alphaCSR[ 255 ][ 378 ],
   alphaCSR[ 255 ][ 379 ],
   alphaCSR[ 255 ][ 380 ],
   alphaCSR[ 255 ][ 381 ],
   alphaCSR[ 255 ][ 382 ],
   alphaCSR[ 255 ][ 383 ],


 doutA1[0],
doutA1[1],
doutA1[2],
doutA1[3],
doutA1[4],
doutA1[5],
doutA1[6],
doutA1[7],
doutA1[8],
doutA1[9],
doutA1[10],
doutA1[11],
doutA1[12],
doutA1[13],
doutA1[14],
doutA1[15],
doutA1[16],
doutA1[17],
doutA1[18],
doutA1[19],
doutA1[20],
doutA1[21],
doutA1[22],
doutA1[23],
doutA1[24],
doutA1[25],
doutA1[26],
doutA1[27],
doutA1[28],
doutA1[29],
doutA1[30],
doutA1[31],
doutA1[32],
doutA1[33],
doutA1[34],
doutA1[35],
doutA1[36],
doutA1[37],
doutA1[38],
doutA1[39],
doutA1[40],
doutA1[41],
doutA1[42],
doutA1[43],
doutA1[44],
doutA1[45],
doutA1[46],
doutA1[47],
doutA1[48],
doutA1[49],
doutA1[50],
doutA1[51],
doutA1[52],
doutA1[53],
doutA1[54],
doutA1[55],
doutA1[56],
doutA1[57],
doutA1[58],
doutA1[59],
doutA1[60],
doutA1[61],
doutA1[62],
doutA1[63],
doutA1[64],
doutA1[65],
doutA1[66],
doutA1[67],
doutA1[68],
doutA1[69],
doutA1[70],
doutA1[71],
doutA1[72],
doutA1[73],
doutA1[74],
doutA1[75],
doutA1[76],
doutA1[77],
doutA1[78],
doutA1[79],
doutA1[80],
doutA1[81],
doutA1[82],
doutA1[83],
doutA1[84],
doutA1[85],
doutA1[86],
doutA1[87],
doutA1[88],
doutA1[89],
doutA1[90],
doutA1[91],
doutA1[92],
doutA1[93],
doutA1[94],
doutA1[95],
doutA1[96],
doutA1[97],
doutA1[98],
doutA1[99],
doutA1[100],
doutA1[101],
doutA1[102],
doutA1[103],
doutA1[104],
doutA1[105],
doutA1[106],
doutA1[107],
doutA1[108],
doutA1[109],
doutA1[110],
doutA1[111],
doutA1[112],
doutA1[113],
doutA1[114],
doutA1[115],
doutA1[116],
doutA1[117],
doutA1[118],
doutA1[119],
doutA1[120],
doutA1[121],
doutA1[122],
doutA1[123],
doutA1[124],
doutA1[125],
doutA1[126],
doutA1[127],
doutA1[128],
doutA1[129],
doutA1[130],
doutA1[131],
doutA1[132],
doutA1[133],
doutA1[134],
doutA1[135],
doutA1[136],
doutA1[137],
doutA1[138],
doutA1[139],
doutA1[140],
doutA1[141],
doutA1[142],
doutA1[143],
doutA1[144],
doutA1[145],
doutA1[146],
doutA1[147],
doutA1[148],
doutA1[149],
doutA1[150],
doutA1[151],
doutA1[152],
doutA1[153],
doutA1[154],
doutA1[155],
doutA1[156],
doutA1[157],
doutA1[158],
doutA1[159],
doutA1[160],
doutA1[161],
doutA1[162],
doutA1[163],
doutA1[164],
doutA1[165],
doutA1[166],
doutA1[167],
doutA1[168],
doutA1[169],
doutA1[170],
doutA1[171],
doutA1[172],
doutA1[173],
doutA1[174],
doutA1[175],
doutA1[176],
doutA1[177],
doutA1[178],
doutA1[179],
doutA1[180],
doutA1[181],
doutA1[182],
doutA1[183],
doutA1[184],
doutA1[185],
doutA1[186],
doutA1[187],
doutA1[188],
doutA1[189],
doutA1[190],
doutA1[191],
doutA1[192],
doutA1[193],
doutA1[194],
doutA1[195],
doutA1[196],
doutA1[197],
doutA1[198],
doutA1[199],
doutA1[200],
doutA1[201],
doutA1[202],
doutA1[203],
doutA1[204],
doutA1[205],
doutA1[206],
doutA1[207],
doutA1[208],
doutA1[209],
doutA1[210],
doutA1[211],
doutA1[212],
doutA1[213],
doutA1[214],
doutA1[215],
doutA1[216],
doutA1[217],
doutA1[218],
doutA1[219],
doutA1[220],
doutA1[221],
doutA1[222],
doutA1[223],
doutA1[224],
doutA1[225],
doutA1[226],
doutA1[227],
doutA1[228],
doutA1[229],
doutA1[230],
doutA1[231],
doutA1[232],
doutA1[233],
doutA1[234],
doutA1[235],
doutA1[236],
doutA1[237],
doutA1[238],
doutA1[239],
doutA1[240],
doutA1[241],
doutA1[242],
doutA1[243],
doutA1[244],
doutA1[245],
doutA1[246],
doutA1[247],
doutA1[248],
doutA1[249],
doutA1[250],
doutA1[251],
doutA1[252],
doutA1[253],
doutA1[254],
doutA1[255],
doutA1[256],
doutA1[257],
doutA1[258],
doutA1[259],
doutA1[260],
doutA1[261],
doutA1[262],
doutA1[263],
doutA1[264],
doutA1[265],
doutA1[266],
doutA1[267],
doutA1[268],
doutA1[269],
doutA1[270],
doutA1[271],
doutA1[272],
doutA1[273],
doutA1[274],
doutA1[275],
doutA1[276],
doutA1[277],
doutA1[278],
doutA1[279],
doutA1[280],
doutA1[281],
doutA1[282],
doutA1[283],
doutA1[284],
doutA1[285],
doutA1[286],
doutA1[287],
doutA1[288],
doutA1[289],
doutA1[290],
doutA1[291],
doutA1[292],
doutA1[293],
doutA1[294],
doutA1[295],
doutA1[296],
doutA1[297],
doutA1[298],
doutA1[299],
doutA1[300],
doutA1[301],
doutA1[302],
doutA1[303],
doutA1[304],
doutA1[305],
doutA1[306],
doutA1[307],
doutA1[308],
doutA1[309],
doutA1[310],
doutA1[311],
doutA1[312],
doutA1[313],
doutA1[314],
doutA1[315],
doutA1[316],
doutA1[317],
doutA1[318],
doutA1[319],
doutA1[320],
doutA1[321],
doutA1[322],
doutA1[323],
doutA1[324],
doutA1[325],
doutA1[326],
doutA1[327],
doutA1[328],
doutA1[329],
doutA1[330],
doutA1[331],
doutA1[332],
doutA1[333],
doutA1[334],
doutA1[335],
doutA1[336],
doutA1[337],
doutA1[338],
doutA1[339],
doutA1[340],
doutA1[341],
doutA1[342],
doutA1[343],
doutA1[344],
doutA1[345],
doutA1[346],
doutA1[347],
doutA1[348],
doutA1[349],
doutA1[350],
doutA1[351],
doutA1[352],
doutA1[353],
doutA1[354],
doutA1[355],
doutA1[356],
doutA1[357],
doutA1[358],
doutA1[359],
doutA1[360],
doutA1[361],
doutA1[362],
doutA1[363],
doutA1[364],
doutA1[365],
doutA1[366],
doutA1[367],
doutA1[368],
doutA1[369],
doutA1[370],
doutA1[371],
doutA1[372],
doutA1[373],
doutA1[374],
doutA1[375],
doutA1[376],
doutA1[377],
doutA1[378],
doutA1[379],
doutA1[380],
doutA1[381],
doutA1[382],
doutA1[383],
doutA1[384],
doutA1[385],
doutA1[386],
doutA1[387],
doutA1[388],
doutA1[389],
doutA1[390],
doutA1[391],
doutA1[392],
doutA1[393],
doutA1[394],
doutA1[395],
doutA1[396],
doutA1[397],
doutA1[398],
doutA1[399],
doutA1[400],
doutA1[401],
doutA1[402],
doutA1[403],
doutA1[404],
doutA1[405],
doutA1[406],
doutA1[407],
doutA1[408],
doutA1[409],
doutA1[410],
doutA1[411],
doutA1[412],
doutA1[413],
doutA1[414],
doutA1[415],
doutA1[416],
doutA1[417],
doutA1[418],
doutA1[419],
doutA1[420],
doutA1[421],
doutA1[422],
doutA1[423],
doutA1[424],
doutA1[425],
doutA1[426],
doutA1[427],
doutA1[428],
doutA1[429],
doutA1[430],
doutA1[431],
doutA1[432],
doutA1[433],
doutA1[434],
doutA1[435],
doutA1[436],
doutA1[437],
doutA1[438],
doutA1[439],
doutA1[440],
doutA1[441],
doutA1[442],
doutA1[443],
doutA1[444],
doutA1[445],
doutA1[446],
doutA1[447],
doutA1[448],
doutA1[449],
doutA1[450],
doutA1[451],
doutA1[452],
doutA1[453],
doutA1[454],
doutA1[455],
doutA1[456],
doutA1[457],
doutA1[458],
doutA1[459],
doutA1[460],
doutA1[461],
doutA1[462],
doutA1[463],
doutA1[464],
doutA1[465],
doutA1[466],
doutA1[467],
doutA1[468],
doutA1[469],
doutA1[470],
doutA1[471],
doutA1[472],
doutA1[473],
doutA1[474],
doutA1[475],
doutA1[476],
doutA1[477],
doutA1[478],
doutA1[479],
doutA1[480],
doutA1[481],
doutA1[482],
doutA1[483],
doutA1[484],
doutA1[485],
doutA1[486],
doutA1[487],
doutA1[488],
doutA1[489],
doutA1[490],
doutA1[491],
doutA1[492],
doutA1[493],
doutA1[494],
doutA1[495],
doutA1[496],
doutA1[497],
doutA1[498],
doutA1[499],
doutA1[500],
doutA1[501],
doutA1[502],
doutA1[503],
doutA1[504],
doutA1[505],
doutA1[506],
doutA1[507],
doutA1[508],
doutA1[509],
doutA1[510],
doutA1[511],
doutA1[512],
doutA1[513],
doutA1[514],
doutA1[515],
doutA1[516],
doutA1[517],
doutA1[518],
doutA1[519],
doutA1[520],
doutA1[521],
doutA1[522],
doutA1[523],
doutA1[524],
doutA1[525],
doutA1[526],
doutA1[527],
doutA1[528],
doutA1[529],
doutA1[530],
doutA1[531],
doutA1[532],
doutA1[533],
doutA1[534],
doutA1[535],
doutA1[536],
doutA1[537],
doutA1[538],
doutA1[539],
doutA1[540],
doutA1[541],
doutA1[542],
doutA1[543],
doutA1[544],
doutA1[545],
doutA1[546],
doutA1[547],
doutA1[548],
doutA1[549],
doutA1[550],
doutA1[551],
doutA1[552],
doutA1[553],
doutA1[554],
doutA1[555],
doutA1[556],
doutA1[557],
doutA1[558],
doutA1[559],
doutA1[560],
doutA1[561],
doutA1[562],
doutA1[563],
doutA1[564],
doutA1[565],
doutA1[566],
doutA1[567],
doutA1[568],
doutA1[569],
doutA1[570],
doutA1[571],
doutA1[572],
doutA1[573],
doutA1[574],
doutA1[575],
doutA1[576],
doutA1[577],
doutA1[578],
doutA1[579],
doutA1[580],
doutA1[581],
doutA1[582],
doutA1[583],
doutA1[584],
doutA1[585],
doutA1[586],
doutA1[587],
doutA1[588],
doutA1[589],
doutA1[590],
doutA1[591],
doutA1[592],
doutA1[593],
doutA1[594],
doutA1[595],
doutA1[596],
doutA1[597],
doutA1[598],
doutA1[599],
doutA1[600],
doutA1[601],
doutA1[602],
doutA1[603],
doutA1[604],
doutA1[605],
doutA1[606],
doutA1[607],
doutA1[608],
doutA1[609],
doutA1[610],
doutA1[611],
doutA1[612],
doutA1[613],
doutA1[614],
doutA1[615],
doutA1[616],
doutA1[617],
doutA1[618],
doutA1[619],
doutA1[620],
doutA1[621],
doutA1[622],
doutA1[623],
doutA1[624],
doutA1[625],
doutA1[626],
doutA1[627],
doutA1[628],
doutA1[629],
doutA1[630],
doutA1[631],
doutA1[632],
doutA1[633],
doutA1[634],
doutA1[635],
doutA1[636],
doutA1[637],
doutA1[638],
doutA1[639],
doutA1[640],
doutA1[641],
doutA1[642],
doutA1[643],
doutA1[644],
doutA1[645],
doutA1[646],
doutA1[647],
doutA1[648],
doutA1[649],
doutA1[650],
doutA1[651],
doutA1[652],
doutA1[653],
doutA1[654],
doutA1[655],
doutA1[656],
doutA1[657],
doutA1[658],
doutA1[659],
doutA1[660],
doutA1[661],
doutA1[662],
doutA1[663],
doutA1[664],
doutA1[665],
doutA1[666],
doutA1[667],
doutA1[668],
doutA1[669],
doutA1[670],
doutA1[671],
doutA1[672],
doutA1[673],
doutA1[674],
doutA1[675],
doutA1[676],
doutA1[677],
doutA1[678],
doutA1[679],
doutA1[680],
doutA1[681],
doutA1[682],
doutA1[683],
doutA1[684],
doutA1[685],
doutA1[686],
doutA1[687],
doutA1[688],
doutA1[689],
doutA1[690],
doutA1[691],
doutA1[692],
doutA1[693],
doutA1[694],
doutA1[695],
doutA1[696],
doutA1[697],
doutA1[698],
doutA1[699],
doutA1[700],
doutA1[701],
doutA1[702],
doutA1[703],
doutA1[704],
doutA1[705],
doutA1[706],
doutA1[707],
doutA1[708],
doutA1[709],
doutA1[710],
doutA1[711],
doutA1[712],
doutA1[713],
doutA1[714],
doutA1[715],
doutA1[716],
doutA1[717],
doutA1[718],
doutA1[719],
doutA1[720],
doutA1[721],
doutA1[722],
doutA1[723],
doutA1[724],
doutA1[725],
doutA1[726],
doutA1[727],
doutA1[728],
doutA1[729],
doutA1[730],
doutA1[731],
doutA1[732],
doutA1[733],
doutA1[734],
doutA1[735],
doutA1[736],
doutA1[737],
doutA1[738],
doutA1[739],
doutA1[740],
doutA1[741],
doutA1[742],
doutA1[743],
doutA1[744],
doutA1[745],
doutA1[746],
doutA1[747],
doutA1[748],
doutA1[749],
doutA1[750],
doutA1[751],
doutA1[752],
doutA1[753],
doutA1[754],
doutA1[755],
doutA1[756],
doutA1[757],
doutA1[758],
doutA1[759],
doutA1[760],
doutA1[761],
doutA1[762],
doutA1[763],
doutA1[764],
doutA1[765],
doutA1[766],
doutA1[767],

B_[0][0][0],
B_[0][1][0],
B_[0][2][0],
B_[1][0][0],
B_[1][1][0],
B_[1][2][0],
B_[2][0][0],
B_[2][1][0],
B_[2][2][0],
B_[3][0][0],
B_[3][1][0],
B_[3][2][0],
B_[4][0][0],
B_[4][1][0],
B_[4][2][0],
B_[5][0][0],
B_[5][1][0],
B_[5][2][0],
B_[6][0][0],
B_[6][1][0],
B_[6][2][0],
B_[7][0][0],
B_[7][1][0],
B_[7][2][0],
B_[8][0][0],
B_[8][1][0],
B_[8][2][0],
B_[9][0][0],
B_[9][1][0],
B_[9][2][0],
B_[10][0][0],
B_[10][1][0],
B_[10][2][0],
B_[11][0][0],
B_[11][1][0],
B_[11][2][0],
B_[12][0][0],
B_[12][1][0],
B_[12][2][0],
B_[13][0][0],
B_[13][1][0],
B_[13][2][0],
B_[14][0][0],
B_[14][1][0],
B_[14][2][0],
B_[15][0][0],
B_[15][1][0],
B_[15][2][0],
B_[0][0][1],
B_[0][1][1],
B_[0][2][1],
B_[1][0][1],
B_[1][1][1],
B_[1][2][1],
B_[2][0][1],
B_[2][1][1],
B_[2][2][1],
B_[3][0][1],
B_[3][1][1],
B_[3][2][1],
B_[4][0][1],
B_[4][1][1],
B_[4][2][1],
B_[5][0][1],
B_[5][1][1],
B_[5][2][1],
B_[6][0][1],
B_[6][1][1],
B_[6][2][1],
B_[7][0][1],
B_[7][1][1],
B_[7][2][1],
B_[8][0][1],
B_[8][1][1],
B_[8][2][1],
B_[9][0][1],
B_[9][1][1],
B_[9][2][1],
B_[10][0][1],
B_[10][1][1],
B_[10][2][1],
B_[11][0][1],
B_[11][1][1],
B_[11][2][1],
B_[12][0][1],
B_[12][1][1],
B_[12][2][1],
B_[13][0][1],
B_[13][1][1],
B_[13][2][1],
B_[14][0][1],
B_[14][1][1],
B_[14][2][1],
B_[15][0][1],
B_[15][1][1],
B_[15][2][1],
B_[0][0][2],
B_[0][1][2],
B_[0][2][2],
B_[1][0][2],
B_[1][1][2],
B_[1][2][2],
B_[2][0][2],
B_[2][1][2],
B_[2][2][2],
B_[3][0][2],
B_[3][1][2],
B_[3][2][2],
B_[4][0][2],
B_[4][1][2],
B_[4][2][2],
B_[5][0][2],
B_[5][1][2],
B_[5][2][2],
B_[6][0][2],
B_[6][1][2],
B_[6][2][2],
B_[7][0][2],
B_[7][1][2],
B_[7][2][2],
B_[8][0][2],
B_[8][1][2],
B_[8][2][2],
B_[9][0][2],
B_[9][1][2],
B_[9][2][2],
B_[10][0][2],
B_[10][1][2],
B_[10][2][2],
B_[11][0][2],
B_[11][1][2],
B_[11][2][2],
B_[12][0][2],
B_[12][1][2],
B_[12][2][2],
B_[13][0][2],
B_[13][1][2],
B_[13][2][2],
B_[14][0][2],
B_[14][1][2],
B_[14][2][2],
B_[15][0][2],
B_[15][1][2],
B_[15][2][2],
B_[0][0][3],
B_[0][1][3],
B_[0][2][3],
B_[1][0][3],
B_[1][1][3],
B_[1][2][3],
B_[2][0][3],
B_[2][1][3],
B_[2][2][3],
B_[3][0][3],
B_[3][1][3],
B_[3][2][3],
B_[4][0][3],
B_[4][1][3],
B_[4][2][3],
B_[5][0][3],
B_[5][1][3],
B_[5][2][3],
B_[6][0][3],
B_[6][1][3],
B_[6][2][3],
B_[7][0][3],
B_[7][1][3],
B_[7][2][3],
B_[8][0][3],
B_[8][1][3],
B_[8][2][3],
B_[9][0][3],
B_[9][1][3],
B_[9][2][3],
B_[10][0][3],
B_[10][1][3],
B_[10][2][3],
B_[11][0][3],
B_[11][1][3],
B_[11][2][3],
B_[12][0][3],
B_[12][1][3],
B_[12][2][3],
B_[13][0][3],
B_[13][1][3],
B_[13][2][3],
B_[14][0][3],
B_[14][1][3],
B_[14][2][3],
B_[15][0][3],
B_[15][1][3],
B_[15][2][3],
B_[0][0][4],
B_[0][1][4],
B_[0][2][4],
B_[1][0][4],
B_[1][1][4],
B_[1][2][4],
B_[2][0][4],
B_[2][1][4],
B_[2][2][4],
B_[3][0][4],
B_[3][1][4],
B_[3][2][4],
B_[4][0][4],
B_[4][1][4],
B_[4][2][4],
B_[5][0][4],
B_[5][1][4],
B_[5][2][4],
B_[6][0][4],
B_[6][1][4],
B_[6][2][4],
B_[7][0][4],
B_[7][1][4],
B_[7][2][4],
B_[8][0][4],
B_[8][1][4],
B_[8][2][4],
B_[9][0][4],
B_[9][1][4],
B_[9][2][4],
B_[10][0][4],
B_[10][1][4],
B_[10][2][4],
B_[11][0][4],
B_[11][1][4],
B_[11][2][4],
B_[12][0][4],
B_[12][1][4],
B_[12][2][4],
B_[13][0][4],
B_[13][1][4],
B_[13][2][4],
B_[14][0][4],
B_[14][1][4],
B_[14][2][4],
B_[15][0][4],
B_[15][1][4],
B_[15][2][4],
B_[0][0][5],
B_[0][1][5],
B_[0][2][5],
B_[1][0][5],
B_[1][1][5],
B_[1][2][5],
B_[2][0][5],
B_[2][1][5],
B_[2][2][5],
B_[3][0][5],
B_[3][1][5],
B_[3][2][5],
B_[4][0][5],
B_[4][1][5],
B_[4][2][5],
B_[5][0][5],
B_[5][1][5],
B_[5][2][5],
B_[6][0][5],
B_[6][1][5],
B_[6][2][5],
B_[7][0][5],
B_[7][1][5],
B_[7][2][5],
B_[8][0][5],
B_[8][1][5],
B_[8][2][5],
B_[9][0][5],
B_[9][1][5],
B_[9][2][5],
B_[10][0][5],
B_[10][1][5],
B_[10][2][5],
B_[11][0][5],
B_[11][1][5],
B_[11][2][5],
B_[12][0][5],
B_[12][1][5],
B_[12][2][5],
B_[13][0][5],
B_[13][1][5],
B_[13][2][5],
B_[14][0][5],
B_[14][1][5],
B_[14][2][5],
B_[15][0][5],
B_[15][1][5],
B_[15][2][5],
B_[0][0][6],
B_[0][1][6],
B_[0][2][6],
B_[1][0][6],
B_[1][1][6],
B_[1][2][6],
B_[2][0][6],
B_[2][1][6],
B_[2][2][6],
B_[3][0][6],
B_[3][1][6],
B_[3][2][6],
B_[4][0][6],
B_[4][1][6],
B_[4][2][6],
B_[5][0][6],
B_[5][1][6],
B_[5][2][6],
B_[6][0][6],
B_[6][1][6],
B_[6][2][6],
B_[7][0][6],
B_[7][1][6],
B_[7][2][6],
B_[8][0][6],
B_[8][1][6],
B_[8][2][6],
B_[9][0][6],
B_[9][1][6],
B_[9][2][6],
B_[10][0][6],
B_[10][1][6],
B_[10][2][6],
B_[11][0][6],
B_[11][1][6],
B_[11][2][6],
B_[12][0][6],
B_[12][1][6],
B_[12][2][6],
B_[13][0][6],
B_[13][1][6],
B_[13][2][6],
B_[14][0][6],
B_[14][1][6],
B_[14][2][6],
B_[15][0][6],
B_[15][1][6],
B_[15][2][6],
B_[0][0][7],
B_[0][1][7],
B_[0][2][7],
B_[1][0][7],
B_[1][1][7],
B_[1][2][7],
B_[2][0][7],
B_[2][1][7],
B_[2][2][7],
B_[3][0][7],
B_[3][1][7],
B_[3][2][7],
B_[4][0][7],
B_[4][1][7],
B_[4][2][7],
B_[5][0][7],
B_[5][1][7],
B_[5][2][7],
B_[6][0][7],
B_[6][1][7],
B_[6][2][7],
B_[7][0][7],
B_[7][1][7],
B_[7][2][7],
B_[8][0][7],
B_[8][1][7],
B_[8][2][7],
B_[9][0][7],
B_[9][1][7],
B_[9][2][7],
B_[10][0][7],
B_[10][1][7],
B_[10][2][7],
B_[11][0][7],
B_[11][1][7],
B_[11][2][7],
B_[12][0][7],
B_[12][1][7],
B_[12][2][7],
B_[13][0][7],
B_[13][1][7],
B_[13][2][7],
B_[14][0][7],
B_[14][1][7],
B_[14][2][7],
B_[15][0][7],
B_[15][1][7],
B_[15][2][7],
B_[0][0][8],
B_[0][1][8],
B_[0][2][8],
B_[1][0][8],
B_[1][1][8],
B_[1][2][8],
B_[2][0][8],
B_[2][1][8],
B_[2][2][8],
B_[3][0][8],
B_[3][1][8],
B_[3][2][8],
B_[4][0][8],
B_[4][1][8],
B_[4][2][8],
B_[5][0][8],
B_[5][1][8],
B_[5][2][8],
B_[6][0][8],
B_[6][1][8],
B_[6][2][8],
B_[7][0][8],
B_[7][1][8],
B_[7][2][8],
B_[8][0][8],
B_[8][1][8],
B_[8][2][8],
B_[9][0][8],
B_[9][1][8],
B_[9][2][8],
B_[10][0][8],
B_[10][1][8],
B_[10][2][8],
B_[11][0][8],
B_[11][1][8],
B_[11][2][8],
B_[12][0][8],
B_[12][1][8],
B_[12][2][8],
B_[13][0][8],
B_[13][1][8],
B_[13][2][8],
B_[14][0][8],
B_[14][1][8],
B_[14][2][8],
B_[15][0][8],
B_[15][1][8],
B_[15][2][8],
B_[0][0][9],
B_[0][1][9],
B_[0][2][9],
B_[1][0][9],
B_[1][1][9],
B_[1][2][9],
B_[2][0][9],
B_[2][1][9],
B_[2][2][9],
B_[3][0][9],
B_[3][1][9],
B_[3][2][9],
B_[4][0][9],
B_[4][1][9],
B_[4][2][9],
B_[5][0][9],
B_[5][1][9],
B_[5][2][9],
B_[6][0][9],
B_[6][1][9],
B_[6][2][9],
B_[7][0][9],
B_[7][1][9],
B_[7][2][9],
B_[8][0][9],
B_[8][1][9],
B_[8][2][9],
B_[9][0][9],
B_[9][1][9],
B_[9][2][9],
B_[10][0][9],
B_[10][1][9],
B_[10][2][9],
B_[11][0][9],
B_[11][1][9],
B_[11][2][9],
B_[12][0][9],
B_[12][1][9],
B_[12][2][9],
B_[13][0][9],
B_[13][1][9],
B_[13][2][9],
B_[14][0][9],
B_[14][1][9],
B_[14][2][9],
B_[15][0][9],
B_[15][1][9],
B_[15][2][9],
B_[0][0][10],
B_[0][1][10],
B_[0][2][10],
B_[1][0][10],
B_[1][1][10],
B_[1][2][10],
B_[2][0][10],
B_[2][1][10],
B_[2][2][10],
B_[3][0][10],
B_[3][1][10],
B_[3][2][10],
B_[4][0][10],
B_[4][1][10],
B_[4][2][10],
B_[5][0][10],
B_[5][1][10],
B_[5][2][10],
B_[6][0][10],
B_[6][1][10],
B_[6][2][10],
B_[7][0][10],
B_[7][1][10],
B_[7][2][10],
B_[8][0][10],
B_[8][1][10],
B_[8][2][10],
B_[9][0][10],
B_[9][1][10],
B_[9][2][10],
B_[10][0][10],
B_[10][1][10],
B_[10][2][10],
B_[11][0][10],
B_[11][1][10],
B_[11][2][10],
B_[12][0][10],
B_[12][1][10],
B_[12][2][10],
B_[13][0][10],
B_[13][1][10],
B_[13][2][10],
B_[14][0][10],
B_[14][1][10],
B_[14][2][10],
B_[15][0][10],
B_[15][1][10],
B_[15][2][10],
B_[0][0][11],
B_[0][1][11],
B_[0][2][11],
B_[1][0][11],
B_[1][1][11],
B_[1][2][11],
B_[2][0][11],
B_[2][1][11],
B_[2][2][11],
B_[3][0][11],
B_[3][1][11],
B_[3][2][11],
B_[4][0][11],
B_[4][1][11],
B_[4][2][11],
B_[5][0][11],
B_[5][1][11],
B_[5][2][11],
B_[6][0][11],
B_[6][1][11],
B_[6][2][11],
B_[7][0][11],
B_[7][1][11],
B_[7][2][11],
B_[8][0][11],
B_[8][1][11],
B_[8][2][11],
B_[9][0][11],
B_[9][1][11],
B_[9][2][11],
B_[10][0][11],
B_[10][1][11],
B_[10][2][11],
B_[11][0][11],
B_[11][1][11],
B_[11][2][11],
B_[12][0][11],
B_[12][1][11],
B_[12][2][11],
B_[13][0][11],
B_[13][1][11],
B_[13][2][11],
B_[14][0][11],
B_[14][1][11],
B_[14][2][11],
B_[15][0][11],
B_[15][1][11],
B_[15][2][11],
B_[0][0][12],
B_[0][1][12],
B_[0][2][12],
B_[1][0][12],
B_[1][1][12],
B_[1][2][12],
B_[2][0][12],
B_[2][1][12],
B_[2][2][12],
B_[3][0][12],
B_[3][1][12],
B_[3][2][12],
B_[4][0][12],
B_[4][1][12],
B_[4][2][12],
B_[5][0][12],
B_[5][1][12],
B_[5][2][12],
B_[6][0][12],
B_[6][1][12],
B_[6][2][12],
B_[7][0][12],
B_[7][1][12],
B_[7][2][12],
B_[8][0][12],
B_[8][1][12],
B_[8][2][12],
B_[9][0][12],
B_[9][1][12],
B_[9][2][12],
B_[10][0][12],
B_[10][1][12],
B_[10][2][12],
B_[11][0][12],
B_[11][1][12],
B_[11][2][12],
B_[12][0][12],
B_[12][1][12],
B_[12][2][12],
B_[13][0][12],
B_[13][1][12],
B_[13][2][12],
B_[14][0][12],
B_[14][1][12],
B_[14][2][12],
B_[15][0][12],
B_[15][1][12],
B_[15][2][12],
B_[0][0][13],
B_[0][1][13],
B_[0][2][13],
B_[1][0][13],
B_[1][1][13],
B_[1][2][13],
B_[2][0][13],
B_[2][1][13],
B_[2][2][13],
B_[3][0][13],
B_[3][1][13],
B_[3][2][13],
B_[4][0][13],
B_[4][1][13],
B_[4][2][13],
B_[5][0][13],
B_[5][1][13],
B_[5][2][13],
B_[6][0][13],
B_[6][1][13],
B_[6][2][13],
B_[7][0][13],
B_[7][1][13],
B_[7][2][13],
B_[8][0][13],
B_[8][1][13],
B_[8][2][13],
B_[9][0][13],
B_[9][1][13],
B_[9][2][13],
B_[10][0][13],
B_[10][1][13],
B_[10][2][13],
B_[11][0][13],
B_[11][1][13],
B_[11][2][13],
B_[12][0][13],
B_[12][1][13],
B_[12][2][13],
B_[13][0][13],
B_[13][1][13],
B_[13][2][13],
B_[14][0][13],
B_[14][1][13],
B_[14][2][13],
B_[15][0][13],
B_[15][1][13],
B_[15][2][13],
B_[0][0][14],
B_[0][1][14],
B_[0][2][14],
B_[1][0][14],
B_[1][1][14],
B_[1][2][14],
B_[2][0][14],
B_[2][1][14],
B_[2][2][14],
B_[3][0][14],
B_[3][1][14],
B_[3][2][14],
B_[4][0][14],
B_[4][1][14],
B_[4][2][14],
B_[5][0][14],
B_[5][1][14],
B_[5][2][14],
B_[6][0][14],
B_[6][1][14],
B_[6][2][14],
B_[7][0][14],
B_[7][1][14],
B_[7][2][14],
B_[8][0][14],
B_[8][1][14],
B_[8][2][14],
B_[9][0][14],
B_[9][1][14],
B_[9][2][14],
B_[10][0][14],
B_[10][1][14],
B_[10][2][14],
B_[11][0][14],
B_[11][1][14],
B_[11][2][14],
B_[12][0][14],
B_[12][1][14],
B_[12][2][14],
B_[13][0][14],
B_[13][1][14],
B_[13][2][14],
B_[14][0][14],
B_[14][1][14],
B_[14][2][14],
B_[15][0][14],
B_[15][1][14],
B_[15][2][14],
B_[0][0][15],
B_[0][1][15],
B_[0][2][15],
B_[1][0][15],
B_[1][1][15],
B_[1][2][15],
B_[2][0][15],
B_[2][1][15],
B_[2][2][15],
B_[3][0][15],
B_[3][1][15],
B_[3][2][15],
B_[4][0][15],
B_[4][1][15],
B_[4][2][15],
B_[5][0][15],
B_[5][1][15],
B_[5][2][15],
B_[6][0][15],
B_[6][1][15],
B_[6][2][15],
B_[7][0][15],
B_[7][1][15],
B_[7][2][15],
B_[8][0][15],
B_[8][1][15],
B_[8][2][15],
B_[9][0][15],
B_[9][1][15],
B_[9][2][15],
B_[10][0][15],
B_[10][1][15],
B_[10][2][15],
B_[11][0][15],
B_[11][1][15],
B_[11][2][15],
B_[12][0][15],
B_[12][1][15],
B_[12][2][15],
B_[13][0][15],
B_[13][1][15],
B_[13][2][15],
B_[14][0][15],
B_[14][1][15],
B_[14][2][15],
B_[15][0][15],
B_[15][1][15],
B_[15][2][15],
B_[0][0][16],
B_[0][1][16],
B_[0][2][16],
B_[1][0][16],
B_[1][1][16],
B_[1][2][16],
B_[2][0][16],
B_[2][1][16],
B_[2][2][16],
B_[3][0][16],
B_[3][1][16],
B_[3][2][16],
B_[4][0][16],
B_[4][1][16],
B_[4][2][16],
B_[5][0][16],
B_[5][1][16],
B_[5][2][16],
B_[6][0][16],
B_[6][1][16],
B_[6][2][16],
B_[7][0][16],
B_[7][1][16],
B_[7][2][16],
B_[8][0][16],
B_[8][1][16],
B_[8][2][16],
B_[9][0][16],
B_[9][1][16],
B_[9][2][16],
B_[10][0][16],
B_[10][1][16],
B_[10][2][16],
B_[11][0][16],
B_[11][1][16],
B_[11][2][16],
B_[12][0][16],
B_[12][1][16],
B_[12][2][16],
B_[13][0][16],
B_[13][1][16],
B_[13][2][16],
B_[14][0][16],
B_[14][1][16],
B_[14][2][16],
B_[15][0][16],
B_[15][1][16],
B_[15][2][16],
B_[0][0][17],
B_[0][1][17],
B_[0][2][17],
B_[1][0][17],
B_[1][1][17],
B_[1][2][17],
B_[2][0][17],
B_[2][1][17],
B_[2][2][17],
B_[3][0][17],
B_[3][1][17],
B_[3][2][17],
B_[4][0][17],
B_[4][1][17],
B_[4][2][17],
B_[5][0][17],
B_[5][1][17],
B_[5][2][17],
B_[6][0][17],
B_[6][1][17],
B_[6][2][17],
B_[7][0][17],
B_[7][1][17],
B_[7][2][17],
B_[8][0][17],
B_[8][1][17],
B_[8][2][17],
B_[9][0][17],
B_[9][1][17],
B_[9][2][17],
B_[10][0][17],
B_[10][1][17],
B_[10][2][17],
B_[11][0][17],
B_[11][1][17],
B_[11][2][17],
B_[12][0][17],
B_[12][1][17],
B_[12][2][17],
B_[13][0][17],
B_[13][1][17],
B_[13][2][17],
B_[14][0][17],
B_[14][1][17],
B_[14][2][17],
B_[15][0][17],
B_[15][1][17],
B_[15][2][17],
B_[0][0][18],
B_[0][1][18],
B_[0][2][18],
B_[1][0][18],
B_[1][1][18],
B_[1][2][18],
B_[2][0][18],
B_[2][1][18],
B_[2][2][18],
B_[3][0][18],
B_[3][1][18],
B_[3][2][18],
B_[4][0][18],
B_[4][1][18],
B_[4][2][18],
B_[5][0][18],
B_[5][1][18],
B_[5][2][18],
B_[6][0][18],
B_[6][1][18],
B_[6][2][18],
B_[7][0][18],
B_[7][1][18],
B_[7][2][18],
B_[8][0][18],
B_[8][1][18],
B_[8][2][18],
B_[9][0][18],
B_[9][1][18],
B_[9][2][18],
B_[10][0][18],
B_[10][1][18],
B_[10][2][18],
B_[11][0][18],
B_[11][1][18],
B_[11][2][18],
B_[12][0][18],
B_[12][1][18],
B_[12][2][18],
B_[13][0][18],
B_[13][1][18],
B_[13][2][18],
B_[14][0][18],
B_[14][1][18],
B_[14][2][18],
B_[15][0][18],
B_[15][1][18],
B_[15][2][18],
B_[0][0][19],
B_[0][1][19],
B_[0][2][19],
B_[1][0][19],
B_[1][1][19],
B_[1][2][19],
B_[2][0][19],
B_[2][1][19],
B_[2][2][19],
B_[3][0][19],
B_[3][1][19],
B_[3][2][19],
B_[4][0][19],
B_[4][1][19],
B_[4][2][19],
B_[5][0][19],
B_[5][1][19],
B_[5][2][19],
B_[6][0][19],
B_[6][1][19],
B_[6][2][19],
B_[7][0][19],
B_[7][1][19],
B_[7][2][19],
B_[8][0][19],
B_[8][1][19],
B_[8][2][19],
B_[9][0][19],
B_[9][1][19],
B_[9][2][19],
B_[10][0][19],
B_[10][1][19],
B_[10][2][19],
B_[11][0][19],
B_[11][1][19],
B_[11][2][19],
B_[12][0][19],
B_[12][1][19],
B_[12][2][19],
B_[13][0][19],
B_[13][1][19],
B_[13][2][19],
B_[14][0][19],
B_[14][1][19],
B_[14][2][19],
B_[15][0][19],
B_[15][1][19],
B_[15][2][19],
B_[0][0][20],
B_[0][1][20],
B_[0][2][20],
B_[1][0][20],
B_[1][1][20],
B_[1][2][20],
B_[2][0][20],
B_[2][1][20],
B_[2][2][20],
B_[3][0][20],
B_[3][1][20],
B_[3][2][20],
B_[4][0][20],
B_[4][1][20],
B_[4][2][20],
B_[5][0][20],
B_[5][1][20],
B_[5][2][20],
B_[6][0][20],
B_[6][1][20],
B_[6][2][20],
B_[7][0][20],
B_[7][1][20],
B_[7][2][20],
B_[8][0][20],
B_[8][1][20],
B_[8][2][20],
B_[9][0][20],
B_[9][1][20],
B_[9][2][20],
B_[10][0][20],
B_[10][1][20],
B_[10][2][20],
B_[11][0][20],
B_[11][1][20],
B_[11][2][20],
B_[12][0][20],
B_[12][1][20],
B_[12][2][20],
B_[13][0][20],
B_[13][1][20],
B_[13][2][20],
B_[14][0][20],
B_[14][1][20],
B_[14][2][20],
B_[15][0][20],
B_[15][1][20],
B_[15][2][20],
B_[0][0][21],
B_[0][1][21],
B_[0][2][21],
B_[1][0][21],
B_[1][1][21],
B_[1][2][21],
B_[2][0][21],
B_[2][1][21],
B_[2][2][21],
B_[3][0][21],
B_[3][1][21],
B_[3][2][21],
B_[4][0][21],
B_[4][1][21],
B_[4][2][21],
B_[5][0][21],
B_[5][1][21],
B_[5][2][21],
B_[6][0][21],
B_[6][1][21],
B_[6][2][21],
B_[7][0][21],
B_[7][1][21],
B_[7][2][21],
B_[8][0][21],
B_[8][1][21],
B_[8][2][21],
B_[9][0][21],
B_[9][1][21],
B_[9][2][21],
B_[10][0][21],
B_[10][1][21],
B_[10][2][21],
B_[11][0][21],
B_[11][1][21],
B_[11][2][21],
B_[12][0][21],
B_[12][1][21],
B_[12][2][21],
B_[13][0][21],
B_[13][1][21],
B_[13][2][21],
B_[14][0][21],
B_[14][1][21],
B_[14][2][21],
B_[15][0][21],
B_[15][1][21],
B_[15][2][21],
B_[0][0][22],
B_[0][1][22],
B_[0][2][22],
B_[1][0][22],
B_[1][1][22],
B_[1][2][22],
B_[2][0][22],
B_[2][1][22],
B_[2][2][22],
B_[3][0][22],
B_[3][1][22],
B_[3][2][22],
B_[4][0][22],
B_[4][1][22],
B_[4][2][22],
B_[5][0][22],
B_[5][1][22],
B_[5][2][22],
B_[6][0][22],
B_[6][1][22],
B_[6][2][22],
B_[7][0][22],
B_[7][1][22],
B_[7][2][22],
B_[8][0][22],
B_[8][1][22],
B_[8][2][22],
B_[9][0][22],
B_[9][1][22],
B_[9][2][22],
B_[10][0][22],
B_[10][1][22],
B_[10][2][22],
B_[11][0][22],
B_[11][1][22],
B_[11][2][22],
B_[12][0][22],
B_[12][1][22],
B_[12][2][22],
B_[13][0][22],
B_[13][1][22],
B_[13][2][22],
B_[14][0][22],
B_[14][1][22],
B_[14][2][22],
B_[15][0][22],
B_[15][1][22],
B_[15][2][22],
B_[0][0][23],
B_[0][1][23],
B_[0][2][23],
B_[1][0][23],
B_[1][1][23],
B_[1][2][23],
B_[2][0][23],
B_[2][1][23],
B_[2][2][23],
B_[3][0][23],
B_[3][1][23],
B_[3][2][23],
B_[4][0][23],
B_[4][1][23],
B_[4][2][23],
B_[5][0][23],
B_[5][1][23],
B_[5][2][23],
B_[6][0][23],
B_[6][1][23],
B_[6][2][23],
B_[7][0][23],
B_[7][1][23],
B_[7][2][23],
B_[8][0][23],
B_[8][1][23],
B_[8][2][23],
B_[9][0][23],
B_[9][1][23],
B_[9][2][23],
B_[10][0][23],
B_[10][1][23],
B_[10][2][23],
B_[11][0][23],
B_[11][1][23],
B_[11][2][23],
B_[12][0][23],
B_[12][1][23],
B_[12][2][23],
B_[13][0][23],
B_[13][1][23],
B_[13][2][23],
B_[14][0][23],
B_[14][1][23],
B_[14][2][23],
B_[15][0][23],
B_[15][1][23],
B_[15][2][23],
B_[0][0][24],
B_[0][1][24],
B_[0][2][24],
B_[1][0][24],
B_[1][1][24],
B_[1][2][24],
B_[2][0][24],
B_[2][1][24],
B_[2][2][24],
B_[3][0][24],
B_[3][1][24],
B_[3][2][24],
B_[4][0][24],
B_[4][1][24],
B_[4][2][24],
B_[5][0][24],
B_[5][1][24],
B_[5][2][24],
B_[6][0][24],
B_[6][1][24],
B_[6][2][24],
B_[7][0][24],
B_[7][1][24],
B_[7][2][24],
B_[8][0][24],
B_[8][1][24],
B_[8][2][24],
B_[9][0][24],
B_[9][1][24],
B_[9][2][24],
B_[10][0][24],
B_[10][1][24],
B_[10][2][24],
B_[11][0][24],
B_[11][1][24],
B_[11][2][24],
B_[12][0][24],
B_[12][1][24],
B_[12][2][24],
B_[13][0][24],
B_[13][1][24],
B_[13][2][24],
B_[14][0][24],
B_[14][1][24],
B_[14][2][24],
B_[15][0][24],
B_[15][1][24],
B_[15][2][24],
B_[0][0][25],
B_[0][1][25],
B_[0][2][25],
B_[1][0][25],
B_[1][1][25],
B_[1][2][25],
B_[2][0][25],
B_[2][1][25],
B_[2][2][25],
B_[3][0][25],
B_[3][1][25],
B_[3][2][25],
B_[4][0][25],
B_[4][1][25],
B_[4][2][25],
B_[5][0][25],
B_[5][1][25],
B_[5][2][25],
B_[6][0][25],
B_[6][1][25],
B_[6][2][25],
B_[7][0][25],
B_[7][1][25],
B_[7][2][25],
B_[8][0][25],
B_[8][1][25],
B_[8][2][25],
B_[9][0][25],
B_[9][1][25],
B_[9][2][25],
B_[10][0][25],
B_[10][1][25],
B_[10][2][25],
B_[11][0][25],
B_[11][1][25],
B_[11][2][25],
B_[12][0][25],
B_[12][1][25],
B_[12][2][25],
B_[13][0][25],
B_[13][1][25],
B_[13][2][25],
B_[14][0][25],
B_[14][1][25],
B_[14][2][25],
B_[15][0][25],
B_[15][1][25],
B_[15][2][25],
B_[0][0][26],
B_[0][1][26],
B_[0][2][26],
B_[1][0][26],
B_[1][1][26],
B_[1][2][26],
B_[2][0][26],
B_[2][1][26],
B_[2][2][26],
B_[3][0][26],
B_[3][1][26],
B_[3][2][26],
B_[4][0][26],
B_[4][1][26],
B_[4][2][26],
B_[5][0][26],
B_[5][1][26],
B_[5][2][26],
B_[6][0][26],
B_[6][1][26],
B_[6][2][26],
B_[7][0][26],
B_[7][1][26],
B_[7][2][26],
B_[8][0][26],
B_[8][1][26],
B_[8][2][26],
B_[9][0][26],
B_[9][1][26],
B_[9][2][26],
B_[10][0][26],
B_[10][1][26],
B_[10][2][26],
B_[11][0][26],
B_[11][1][26],
B_[11][2][26],
B_[12][0][26],
B_[12][1][26],
B_[12][2][26],
B_[13][0][26],
B_[13][1][26],
B_[13][2][26],
B_[14][0][26],
B_[14][1][26],
B_[14][2][26],
B_[15][0][26],
B_[15][1][26],
B_[15][2][26],
B_[0][0][27],
B_[0][1][27],
B_[0][2][27],
B_[1][0][27],
B_[1][1][27],
B_[1][2][27],
B_[2][0][27],
B_[2][1][27],
B_[2][2][27],
B_[3][0][27],
B_[3][1][27],
B_[3][2][27],
B_[4][0][27],
B_[4][1][27],
B_[4][2][27],
B_[5][0][27],
B_[5][1][27],
B_[5][2][27],
B_[6][0][27],
B_[6][1][27],
B_[6][2][27],
B_[7][0][27],
B_[7][1][27],
B_[7][2][27],
B_[8][0][27],
B_[8][1][27],
B_[8][2][27],
B_[9][0][27],
B_[9][1][27],
B_[9][2][27],
B_[10][0][27],
B_[10][1][27],
B_[10][2][27],
B_[11][0][27],
B_[11][1][27],
B_[11][2][27],
B_[12][0][27],
B_[12][1][27],
B_[12][2][27],
B_[13][0][27],
B_[13][1][27],
B_[13][2][27],
B_[14][0][27],
B_[14][1][27],
B_[14][2][27],
B_[15][0][27],
B_[15][1][27],
B_[15][2][27],
B_[0][0][28],
B_[0][1][28],
B_[0][2][28],
B_[1][0][28],
B_[1][1][28],
B_[1][2][28],
B_[2][0][28],
B_[2][1][28],
B_[2][2][28],
B_[3][0][28],
B_[3][1][28],
B_[3][2][28],
B_[4][0][28],
B_[4][1][28],
B_[4][2][28],
B_[5][0][28],
B_[5][1][28],
B_[5][2][28],
B_[6][0][28],
B_[6][1][28],
B_[6][2][28],
B_[7][0][28],
B_[7][1][28],
B_[7][2][28],
B_[8][0][28],
B_[8][1][28],
B_[8][2][28],
B_[9][0][28],
B_[9][1][28],
B_[9][2][28],
B_[10][0][28],
B_[10][1][28],
B_[10][2][28],
B_[11][0][28],
B_[11][1][28],
B_[11][2][28],
B_[12][0][28],
B_[12][1][28],
B_[12][2][28],
B_[13][0][28],
B_[13][1][28],
B_[13][2][28],
B_[14][0][28],
B_[14][1][28],
B_[14][2][28],
B_[15][0][28],
B_[15][1][28],
B_[15][2][28],
B_[0][0][29],
B_[0][1][29],
B_[0][2][29],
B_[1][0][29],
B_[1][1][29],
B_[1][2][29],
B_[2][0][29],
B_[2][1][29],
B_[2][2][29],
B_[3][0][29],
B_[3][1][29],
B_[3][2][29],
B_[4][0][29],
B_[4][1][29],
B_[4][2][29],
B_[5][0][29],
B_[5][1][29],
B_[5][2][29],
B_[6][0][29],
B_[6][1][29],
B_[6][2][29],
B_[7][0][29],
B_[7][1][29],
B_[7][2][29],
B_[8][0][29],
B_[8][1][29],
B_[8][2][29],
B_[9][0][29],
B_[9][1][29],
B_[9][2][29],
B_[10][0][29],
B_[10][1][29],
B_[10][2][29],
B_[11][0][29],
B_[11][1][29],
B_[11][2][29],
B_[12][0][29],
B_[12][1][29],
B_[12][2][29],
B_[13][0][29],
B_[13][1][29],
B_[13][2][29],
B_[14][0][29],
B_[14][1][29],
B_[14][2][29],
B_[15][0][29],
B_[15][1][29],
B_[15][2][29],
B_[0][0][30],
B_[0][1][30],
B_[0][2][30],
B_[1][0][30],
B_[1][1][30],
B_[1][2][30],
B_[2][0][30],
B_[2][1][30],
B_[2][2][30],
B_[3][0][30],
B_[3][1][30],
B_[3][2][30],
B_[4][0][30],
B_[4][1][30],
B_[4][2][30],
B_[5][0][30],
B_[5][1][30],
B_[5][2][30],
B_[6][0][30],
B_[6][1][30],
B_[6][2][30],
B_[7][0][30],
B_[7][1][30],
B_[7][2][30],
B_[8][0][30],
B_[8][1][30],
B_[8][2][30],
B_[9][0][30],
B_[9][1][30],
B_[9][2][30],
B_[10][0][30],
B_[10][1][30],
B_[10][2][30],
B_[11][0][30],
B_[11][1][30],
B_[11][2][30],
B_[12][0][30],
B_[12][1][30],
B_[12][2][30],
B_[13][0][30],
B_[13][1][30],
B_[13][2][30],
B_[14][0][30],
B_[14][1][30],
B_[14][2][30],
B_[15][0][30],
B_[15][1][30],
B_[15][2][30],
B_[0][0][31],
B_[0][1][31],
B_[0][2][31],
B_[1][0][31],
B_[1][1][31],
B_[1][2][31],
B_[2][0][31],
B_[2][1][31],
B_[2][2][31],
B_[3][0][31],
B_[3][1][31],
B_[3][2][31],
B_[4][0][31],
B_[4][1][31],
B_[4][2][31],
B_[5][0][31],
B_[5][1][31],
B_[5][2][31],
B_[6][0][31],
B_[6][1][31],
B_[6][2][31],
B_[7][0][31],
B_[7][1][31],
B_[7][2][31],
B_[8][0][31],
B_[8][1][31],
B_[8][2][31],
B_[9][0][31],
B_[9][1][31],
B_[9][2][31],
B_[10][0][31],
B_[10][1][31],
B_[10][2][31],
B_[11][0][31],
B_[11][1][31],
B_[11][2][31],
B_[12][0][31],
B_[12][1][31],
B_[12][2][31],
B_[13][0][31],
B_[13][1][31],
B_[13][2][31],
B_[14][0][31],
B_[14][1][31],
B_[14][2][31],
B_[15][0][31],
B_[15][1][31],
B_[15][2][31],
B_[0][0][32],
B_[0][1][32],
B_[0][2][32],
B_[1][0][32],
B_[1][1][32],
B_[1][2][32],
B_[2][0][32],
B_[2][1][32],
B_[2][2][32],
B_[3][0][32],
B_[3][1][32],
B_[3][2][32],
B_[4][0][32],
B_[4][1][32],
B_[4][2][32],
B_[5][0][32],
B_[5][1][32],
B_[5][2][32],
B_[6][0][32],
B_[6][1][32],
B_[6][2][32],
B_[7][0][32],
B_[7][1][32],
B_[7][2][32],
B_[8][0][32],
B_[8][1][32],
B_[8][2][32],
B_[9][0][32],
B_[9][1][32],
B_[9][2][32],
B_[10][0][32],
B_[10][1][32],
B_[10][2][32],
B_[11][0][32],
B_[11][1][32],
B_[11][2][32],
B_[12][0][32],
B_[12][1][32],
B_[12][2][32],
B_[13][0][32],
B_[13][1][32],
B_[13][2][32],
B_[14][0][32],
B_[14][1][32],
B_[14][2][32],
B_[15][0][32],
B_[15][1][32],
B_[15][2][32],
B_[0][0][33],
B_[0][1][33],
B_[0][2][33],
B_[1][0][33],
B_[1][1][33],
B_[1][2][33],
B_[2][0][33],
B_[2][1][33],
B_[2][2][33],
B_[3][0][33],
B_[3][1][33],
B_[3][2][33],
B_[4][0][33],
B_[4][1][33],
B_[4][2][33],
B_[5][0][33],
B_[5][1][33],
B_[5][2][33],
B_[6][0][33],
B_[6][1][33],
B_[6][2][33],
B_[7][0][33],
B_[7][1][33],
B_[7][2][33],
B_[8][0][33],
B_[8][1][33],
B_[8][2][33],
B_[9][0][33],
B_[9][1][33],
B_[9][2][33],
B_[10][0][33],
B_[10][1][33],
B_[10][2][33],
B_[11][0][33],
B_[11][1][33],
B_[11][2][33],
B_[12][0][33],
B_[12][1][33],
B_[12][2][33],
B_[13][0][33],
B_[13][1][33],
B_[13][2][33],
B_[14][0][33],
B_[14][1][33],
B_[14][2][33],
B_[15][0][33],
B_[15][1][33],
B_[15][2][33],
B_[0][0][34],
B_[0][1][34],
B_[0][2][34],
B_[1][0][34],
B_[1][1][34],
B_[1][2][34],
B_[2][0][34],
B_[2][1][34],
B_[2][2][34],
B_[3][0][34],
B_[3][1][34],
B_[3][2][34],
B_[4][0][34],
B_[4][1][34],
B_[4][2][34],
B_[5][0][34],
B_[5][1][34],
B_[5][2][34],
B_[6][0][34],
B_[6][1][34],
B_[6][2][34],
B_[7][0][34],
B_[7][1][34],
B_[7][2][34],
B_[8][0][34],
B_[8][1][34],
B_[8][2][34],
B_[9][0][34],
B_[9][1][34],
B_[9][2][34],
B_[10][0][34],
B_[10][1][34],
B_[10][2][34],
B_[11][0][34],
B_[11][1][34],
B_[11][2][34],
B_[12][0][34],
B_[12][1][34],
B_[12][2][34],
B_[13][0][34],
B_[13][1][34],
B_[13][2][34],
B_[14][0][34],
B_[14][1][34],
B_[14][2][34],
B_[15][0][34],
B_[15][1][34],
B_[15][2][34],
B_[0][0][35],
B_[0][1][35],
B_[0][2][35],
B_[1][0][35],
B_[1][1][35],
B_[1][2][35],
B_[2][0][35],
B_[2][1][35],
B_[2][2][35],
B_[3][0][35],
B_[3][1][35],
B_[3][2][35],
B_[4][0][35],
B_[4][1][35],
B_[4][2][35],
B_[5][0][35],
B_[5][1][35],
B_[5][2][35],
B_[6][0][35],
B_[6][1][35],
B_[6][2][35],
B_[7][0][35],
B_[7][1][35],
B_[7][2][35],
B_[8][0][35],
B_[8][1][35],
B_[8][2][35],
B_[9][0][35],
B_[9][1][35],
B_[9][2][35],
B_[10][0][35],
B_[10][1][35],
B_[10][2][35],
B_[11][0][35],
B_[11][1][35],
B_[11][2][35],
B_[12][0][35],
B_[12][1][35],
B_[12][2][35],
B_[13][0][35],
B_[13][1][35],
B_[13][2][35],
B_[14][0][35],
B_[14][1][35],
B_[14][2][35],
B_[15][0][35],
B_[15][1][35],
B_[15][2][35],
B_[0][0][36],
B_[0][1][36],
B_[0][2][36],
B_[1][0][36],
B_[1][1][36],
B_[1][2][36],
B_[2][0][36],
B_[2][1][36],
B_[2][2][36],
B_[3][0][36],
B_[3][1][36],
B_[3][2][36],
B_[4][0][36],
B_[4][1][36],
B_[4][2][36],
B_[5][0][36],
B_[5][1][36],
B_[5][2][36],
B_[6][0][36],
B_[6][1][36],
B_[6][2][36],
B_[7][0][36],
B_[7][1][36],
B_[7][2][36],
B_[8][0][36],
B_[8][1][36],
B_[8][2][36],
B_[9][0][36],
B_[9][1][36],
B_[9][2][36],
B_[10][0][36],
B_[10][1][36],
B_[10][2][36],
B_[11][0][36],
B_[11][1][36],
B_[11][2][36],
B_[12][0][36],
B_[12][1][36],
B_[12][2][36],
B_[13][0][36],
B_[13][1][36],
B_[13][2][36],
B_[14][0][36],
B_[14][1][36],
B_[14][2][36],
B_[15][0][36],
B_[15][1][36],
B_[15][2][36],
B_[0][0][37],
B_[0][1][37],
B_[0][2][37],
B_[1][0][37],
B_[1][1][37],
B_[1][2][37],
B_[2][0][37],
B_[2][1][37],
B_[2][2][37],
B_[3][0][37],
B_[3][1][37],
B_[3][2][37],
B_[4][0][37],
B_[4][1][37],
B_[4][2][37],
B_[5][0][37],
B_[5][1][37],
B_[5][2][37],
B_[6][0][37],
B_[6][1][37],
B_[6][2][37],
B_[7][0][37],
B_[7][1][37],
B_[7][2][37],
B_[8][0][37],
B_[8][1][37],
B_[8][2][37],
B_[9][0][37],
B_[9][1][37],
B_[9][2][37],
B_[10][0][37],
B_[10][1][37],
B_[10][2][37],
B_[11][0][37],
B_[11][1][37],
B_[11][2][37],
B_[12][0][37],
B_[12][1][37],
B_[12][2][37],
B_[13][0][37],
B_[13][1][37],
B_[13][2][37],
B_[14][0][37],
B_[14][1][37],
B_[14][2][37],
B_[15][0][37],
B_[15][1][37],
B_[15][2][37],
B_[0][0][38],
B_[0][1][38],
B_[0][2][38],
B_[1][0][38],
B_[1][1][38],
B_[1][2][38],
B_[2][0][38],
B_[2][1][38],
B_[2][2][38],
B_[3][0][38],
B_[3][1][38],
B_[3][2][38],
B_[4][0][38],
B_[4][1][38],
B_[4][2][38],
B_[5][0][38],
B_[5][1][38],
B_[5][2][38],
B_[6][0][38],
B_[6][1][38],
B_[6][2][38],
B_[7][0][38],
B_[7][1][38],
B_[7][2][38],
B_[8][0][38],
B_[8][1][38],
B_[8][2][38],
B_[9][0][38],
B_[9][1][38],
B_[9][2][38],
B_[10][0][38],
B_[10][1][38],
B_[10][2][38],
B_[11][0][38],
B_[11][1][38],
B_[11][2][38],
B_[12][0][38],
B_[12][1][38],
B_[12][2][38],
B_[13][0][38],
B_[13][1][38],
B_[13][2][38],
B_[14][0][38],
B_[14][1][38],
B_[14][2][38],
B_[15][0][38],
B_[15][1][38],
B_[15][2][38],
B_[0][0][39],
B_[0][1][39],
B_[0][2][39],
B_[1][0][39],
B_[1][1][39],
B_[1][2][39],
B_[2][0][39],
B_[2][1][39],
B_[2][2][39],
B_[3][0][39],
B_[3][1][39],
B_[3][2][39],
B_[4][0][39],
B_[4][1][39],
B_[4][2][39],
B_[5][0][39],
B_[5][1][39],
B_[5][2][39],
B_[6][0][39],
B_[6][1][39],
B_[6][2][39],
B_[7][0][39],
B_[7][1][39],
B_[7][2][39],
B_[8][0][39],
B_[8][1][39],
B_[8][2][39],
B_[9][0][39],
B_[9][1][39],
B_[9][2][39],
B_[10][0][39],
B_[10][1][39],
B_[10][2][39],
B_[11][0][39],
B_[11][1][39],
B_[11][2][39],
B_[12][0][39],
B_[12][1][39],
B_[12][2][39],
B_[13][0][39],
B_[13][1][39],
B_[13][2][39],
B_[14][0][39],
B_[14][1][39],
B_[14][2][39],
B_[15][0][39],
B_[15][1][39],
B_[15][2][39],
B_[0][0][40],
B_[0][1][40],
B_[0][2][40],
B_[1][0][40],
B_[1][1][40],
B_[1][2][40],
B_[2][0][40],
B_[2][1][40],
B_[2][2][40],
B_[3][0][40],
B_[3][1][40],
B_[3][2][40],
B_[4][0][40],
B_[4][1][40],
B_[4][2][40],
B_[5][0][40],
B_[5][1][40],
B_[5][2][40],
B_[6][0][40],
B_[6][1][40],
B_[6][2][40],
B_[7][0][40],
B_[7][1][40],
B_[7][2][40],
B_[8][0][40],
B_[8][1][40],
B_[8][2][40],
B_[9][0][40],
B_[9][1][40],
B_[9][2][40],
B_[10][0][40],
B_[10][1][40],
B_[10][2][40],
B_[11][0][40],
B_[11][1][40],
B_[11][2][40],
B_[12][0][40],
B_[12][1][40],
B_[12][2][40],
B_[13][0][40],
B_[13][1][40],
B_[13][2][40],
B_[14][0][40],
B_[14][1][40],
B_[14][2][40],
B_[15][0][40],
B_[15][1][40],
B_[15][2][40],
B_[0][0][41],
B_[0][1][41],
B_[0][2][41],
B_[1][0][41],
B_[1][1][41],
B_[1][2][41],
B_[2][0][41],
B_[2][1][41],
B_[2][2][41],
B_[3][0][41],
B_[3][1][41],
B_[3][2][41],
B_[4][0][41],
B_[4][1][41],
B_[4][2][41],
B_[5][0][41],
B_[5][1][41],
B_[5][2][41],
B_[6][0][41],
B_[6][1][41],
B_[6][2][41],
B_[7][0][41],
B_[7][1][41],
B_[7][2][41],
B_[8][0][41],
B_[8][1][41],
B_[8][2][41],
B_[9][0][41],
B_[9][1][41],
B_[9][2][41],
B_[10][0][41],
B_[10][1][41],
B_[10][2][41],
B_[11][0][41],
B_[11][1][41],
B_[11][2][41],
B_[12][0][41],
B_[12][1][41],
B_[12][2][41],
B_[13][0][41],
B_[13][1][41],
B_[13][2][41],
B_[14][0][41],
B_[14][1][41],
B_[14][2][41],
B_[15][0][41],
B_[15][1][41],
B_[15][2][41],
B_[0][0][42],
B_[0][1][42],
B_[0][2][42],
B_[1][0][42],
B_[1][1][42],
B_[1][2][42],
B_[2][0][42],
B_[2][1][42],
B_[2][2][42],
B_[3][0][42],
B_[3][1][42],
B_[3][2][42],
B_[4][0][42],
B_[4][1][42],
B_[4][2][42],
B_[5][0][42],
B_[5][1][42],
B_[5][2][42],
B_[6][0][42],
B_[6][1][42],
B_[6][2][42],
B_[7][0][42],
B_[7][1][42],
B_[7][2][42],
B_[8][0][42],
B_[8][1][42],
B_[8][2][42],
B_[9][0][42],
B_[9][1][42],
B_[9][2][42],
B_[10][0][42],
B_[10][1][42],
B_[10][2][42],
B_[11][0][42],
B_[11][1][42],
B_[11][2][42],
B_[12][0][42],
B_[12][1][42],
B_[12][2][42],
B_[13][0][42],
B_[13][1][42],
B_[13][2][42],
B_[14][0][42],
B_[14][1][42],
B_[14][2][42],
B_[15][0][42],
B_[15][1][42],
B_[15][2][42],
B_[0][0][43],
B_[0][1][43],
B_[0][2][43],
B_[1][0][43],
B_[1][1][43],
B_[1][2][43],
B_[2][0][43],
B_[2][1][43],
B_[2][2][43],
B_[3][0][43],
B_[3][1][43],
B_[3][2][43],
B_[4][0][43],
B_[4][1][43],
B_[4][2][43],
B_[5][0][43],
B_[5][1][43],
B_[5][2][43],
B_[6][0][43],
B_[6][1][43],
B_[6][2][43],
B_[7][0][43],
B_[7][1][43],
B_[7][2][43],
B_[8][0][43],
B_[8][1][43],
B_[8][2][43],
B_[9][0][43],
B_[9][1][43],
B_[9][2][43],
B_[10][0][43],
B_[10][1][43],
B_[10][2][43],
B_[11][0][43],
B_[11][1][43],
B_[11][2][43],
B_[12][0][43],
B_[12][1][43],
B_[12][2][43],
B_[13][0][43],
B_[13][1][43],
B_[13][2][43],
B_[14][0][43],
B_[14][1][43],
B_[14][2][43],
B_[15][0][43],
B_[15][1][43],
B_[15][2][43],
B_[0][0][44],
B_[0][1][44],
B_[0][2][44],
B_[1][0][44],
B_[1][1][44],
B_[1][2][44],
B_[2][0][44],
B_[2][1][44],
B_[2][2][44],
B_[3][0][44],
B_[3][1][44],
B_[3][2][44],
B_[4][0][44],
B_[4][1][44],
B_[4][2][44],
B_[5][0][44],
B_[5][1][44],
B_[5][2][44],
B_[6][0][44],
B_[6][1][44],
B_[6][2][44],
B_[7][0][44],
B_[7][1][44],
B_[7][2][44],
B_[8][0][44],
B_[8][1][44],
B_[8][2][44],
B_[9][0][44],
B_[9][1][44],
B_[9][2][44],
B_[10][0][44],
B_[10][1][44],
B_[10][2][44],
B_[11][0][44],
B_[11][1][44],
B_[11][2][44],
B_[12][0][44],
B_[12][1][44],
B_[12][2][44],
B_[13][0][44],
B_[13][1][44],
B_[13][2][44],
B_[14][0][44],
B_[14][1][44],
B_[14][2][44],
B_[15][0][44],
B_[15][1][44],
B_[15][2][44],
B_[0][0][45],
B_[0][1][45],
B_[0][2][45],
B_[1][0][45],
B_[1][1][45],
B_[1][2][45],
B_[2][0][45],
B_[2][1][45],
B_[2][2][45],
B_[3][0][45],
B_[3][1][45],
B_[3][2][45],
B_[4][0][45],
B_[4][1][45],
B_[4][2][45],
B_[5][0][45],
B_[5][1][45],
B_[5][2][45],
B_[6][0][45],
B_[6][1][45],
B_[6][2][45],
B_[7][0][45],
B_[7][1][45],
B_[7][2][45],
B_[8][0][45],
B_[8][1][45],
B_[8][2][45],
B_[9][0][45],
B_[9][1][45],
B_[9][2][45],
B_[10][0][45],
B_[10][1][45],
B_[10][2][45],
B_[11][0][45],
B_[11][1][45],
B_[11][2][45],
B_[12][0][45],
B_[12][1][45],
B_[12][2][45],
B_[13][0][45],
B_[13][1][45],
B_[13][2][45],
B_[14][0][45],
B_[14][1][45],
B_[14][2][45],
B_[15][0][45],
B_[15][1][45],
B_[15][2][45],
B_[0][0][46],
B_[0][1][46],
B_[0][2][46],
B_[1][0][46],
B_[1][1][46],
B_[1][2][46],
B_[2][0][46],
B_[2][1][46],
B_[2][2][46],
B_[3][0][46],
B_[3][1][46],
B_[3][2][46],
B_[4][0][46],
B_[4][1][46],
B_[4][2][46],
B_[5][0][46],
B_[5][1][46],
B_[5][2][46],
B_[6][0][46],
B_[6][1][46],
B_[6][2][46],
B_[7][0][46],
B_[7][1][46],
B_[7][2][46],
B_[8][0][46],
B_[8][1][46],
B_[8][2][46],
B_[9][0][46],
B_[9][1][46],
B_[9][2][46],
B_[10][0][46],
B_[10][1][46],
B_[10][2][46],
B_[11][0][46],
B_[11][1][46],
B_[11][2][46],
B_[12][0][46],
B_[12][1][46],
B_[12][2][46],
B_[13][0][46],
B_[13][1][46],
B_[13][2][46],
B_[14][0][46],
B_[14][1][46],
B_[14][2][46],
B_[15][0][46],
B_[15][1][46],
B_[15][2][46],
B_[0][0][47],
B_[0][1][47],
B_[0][2][47],
B_[1][0][47],
B_[1][1][47],
B_[1][2][47],
B_[2][0][47],
B_[2][1][47],
B_[2][2][47],
B_[3][0][47],
B_[3][1][47],
B_[3][2][47],
B_[4][0][47],
B_[4][1][47],
B_[4][2][47],
B_[5][0][47],
B_[5][1][47],
B_[5][2][47],
B_[6][0][47],
B_[6][1][47],
B_[6][2][47],
B_[7][0][47],
B_[7][1][47],
B_[7][2][47],
B_[8][0][47],
B_[8][1][47],
B_[8][2][47],
B_[9][0][47],
B_[9][1][47],
B_[9][2][47],
B_[10][0][47],
B_[10][1][47],
B_[10][2][47],
B_[11][0][47],
B_[11][1][47],
B_[11][2][47],
B_[12][0][47],
B_[12][1][47],
B_[12][2][47],
B_[13][0][47],
B_[13][1][47],
B_[13][2][47],
B_[14][0][47],
B_[14][1][47],
B_[14][2][47],
B_[15][0][47],
B_[15][1][47],
B_[15][2][47],
B_[0][0][48],
B_[0][1][48],
B_[0][2][48],
B_[1][0][48],
B_[1][1][48],
B_[1][2][48],
B_[2][0][48],
B_[2][1][48],
B_[2][2][48],
B_[3][0][48],
B_[3][1][48],
B_[3][2][48],
B_[4][0][48],
B_[4][1][48],
B_[4][2][48],
B_[5][0][48],
B_[5][1][48],
B_[5][2][48],
B_[6][0][48],
B_[6][1][48],
B_[6][2][48],
B_[7][0][48],
B_[7][1][48],
B_[7][2][48],
B_[8][0][48],
B_[8][1][48],
B_[8][2][48],
B_[9][0][48],
B_[9][1][48],
B_[9][2][48],
B_[10][0][48],
B_[10][1][48],
B_[10][2][48],
B_[11][0][48],
B_[11][1][48],
B_[11][2][48],
B_[12][0][48],
B_[12][1][48],
B_[12][2][48],
B_[13][0][48],
B_[13][1][48],
B_[13][2][48],
B_[14][0][48],
B_[14][1][48],
B_[14][2][48],
B_[15][0][48],
B_[15][1][48],
B_[15][2][48],
B_[0][0][49],
B_[0][1][49],
B_[0][2][49],
B_[1][0][49],
B_[1][1][49],
B_[1][2][49],
B_[2][0][49],
B_[2][1][49],
B_[2][2][49],
B_[3][0][49],
B_[3][1][49],
B_[3][2][49],
B_[4][0][49],
B_[4][1][49],
B_[4][2][49],
B_[5][0][49],
B_[5][1][49],
B_[5][2][49],
B_[6][0][49],
B_[6][1][49],
B_[6][2][49],
B_[7][0][49],
B_[7][1][49],
B_[7][2][49],
B_[8][0][49],
B_[8][1][49],
B_[8][2][49],
B_[9][0][49],
B_[9][1][49],
B_[9][2][49],
B_[10][0][49],
B_[10][1][49],
B_[10][2][49],
B_[11][0][49],
B_[11][1][49],
B_[11][2][49],
B_[12][0][49],
B_[12][1][49],
B_[12][2][49],
B_[13][0][49],
B_[13][1][49],
B_[13][2][49],
B_[14][0][49],
B_[14][1][49],
B_[14][2][49],
B_[15][0][49],
B_[15][1][49],
B_[15][2][49],
B_[0][0][50],
B_[0][1][50],
B_[0][2][50],
B_[1][0][50],
B_[1][1][50],
B_[1][2][50],
B_[2][0][50],
B_[2][1][50],
B_[2][2][50],
B_[3][0][50],
B_[3][1][50],
B_[3][2][50],
B_[4][0][50],
B_[4][1][50],
B_[4][2][50],
B_[5][0][50],
B_[5][1][50],
B_[5][2][50],
B_[6][0][50],
B_[6][1][50],
B_[6][2][50],
B_[7][0][50],
B_[7][1][50],
B_[7][2][50],
B_[8][0][50],
B_[8][1][50],
B_[8][2][50],
B_[9][0][50],
B_[9][1][50],
B_[9][2][50],
B_[10][0][50],
B_[10][1][50],
B_[10][2][50],
B_[11][0][50],
B_[11][1][50],
B_[11][2][50],
B_[12][0][50],
B_[12][1][50],
B_[12][2][50],
B_[13][0][50],
B_[13][1][50],
B_[13][2][50],
B_[14][0][50],
B_[14][1][50],
B_[14][2][50],
B_[15][0][50],
B_[15][1][50],
B_[15][2][50],
B_[0][0][51],
B_[0][1][51],
B_[0][2][51],
B_[1][0][51],
B_[1][1][51],
B_[1][2][51],
B_[2][0][51],
B_[2][1][51],
B_[2][2][51],
B_[3][0][51],
B_[3][1][51],
B_[3][2][51],
B_[4][0][51],
B_[4][1][51],
B_[4][2][51],
B_[5][0][51],
B_[5][1][51],
B_[5][2][51],
B_[6][0][51],
B_[6][1][51],
B_[6][2][51],
B_[7][0][51],
B_[7][1][51],
B_[7][2][51],
B_[8][0][51],
B_[8][1][51],
B_[8][2][51],
B_[9][0][51],
B_[9][1][51],
B_[9][2][51],
B_[10][0][51],
B_[10][1][51],
B_[10][2][51],
B_[11][0][51],
B_[11][1][51],
B_[11][2][51],
B_[12][0][51],
B_[12][1][51],
B_[12][2][51],
B_[13][0][51],
B_[13][1][51],
B_[13][2][51],
B_[14][0][51],
B_[14][1][51],
B_[14][2][51],
B_[15][0][51],
B_[15][1][51],
B_[15][2][51],
B_[0][0][52],
B_[0][1][52],
B_[0][2][52],
B_[1][0][52],
B_[1][1][52],
B_[1][2][52],
B_[2][0][52],
B_[2][1][52],
B_[2][2][52],
B_[3][0][52],
B_[3][1][52],
B_[3][2][52],
B_[4][0][52],
B_[4][1][52],
B_[4][2][52],
B_[5][0][52],
B_[5][1][52],
B_[5][2][52],
B_[6][0][52],
B_[6][1][52],
B_[6][2][52],
B_[7][0][52],
B_[7][1][52],
B_[7][2][52],
B_[8][0][52],
B_[8][1][52],
B_[8][2][52],
B_[9][0][52],
B_[9][1][52],
B_[9][2][52],
B_[10][0][52],
B_[10][1][52],
B_[10][2][52],
B_[11][0][52],
B_[11][1][52],
B_[11][2][52],
B_[12][0][52],
B_[12][1][52],
B_[12][2][52],
B_[13][0][52],
B_[13][1][52],
B_[13][2][52],
B_[14][0][52],
B_[14][1][52],
B_[14][2][52],
B_[15][0][52],
B_[15][1][52],
B_[15][2][52],
B_[0][0][53],
B_[0][1][53],
B_[0][2][53],
B_[1][0][53],
B_[1][1][53],
B_[1][2][53],
B_[2][0][53],
B_[2][1][53],
B_[2][2][53],
B_[3][0][53],
B_[3][1][53],
B_[3][2][53],
B_[4][0][53],
B_[4][1][53],
B_[4][2][53],
B_[5][0][53],
B_[5][1][53],
B_[5][2][53],
B_[6][0][53],
B_[6][1][53],
B_[6][2][53],
B_[7][0][53],
B_[7][1][53],
B_[7][2][53],
B_[8][0][53],
B_[8][1][53],
B_[8][2][53],
B_[9][0][53],
B_[9][1][53],
B_[9][2][53],
B_[10][0][53],
B_[10][1][53],
B_[10][2][53],
B_[11][0][53],
B_[11][1][53],
B_[11][2][53],
B_[12][0][53],
B_[12][1][53],
B_[12][2][53],
B_[13][0][53],
B_[13][1][53],
B_[13][2][53],
B_[14][0][53],
B_[14][1][53],
B_[14][2][53],
B_[15][0][53],
B_[15][1][53],
B_[15][2][53],
B_[0][0][54],
B_[0][1][54],
B_[0][2][54],
B_[1][0][54],
B_[1][1][54],
B_[1][2][54],
B_[2][0][54],
B_[2][1][54],
B_[2][2][54],
B_[3][0][54],
B_[3][1][54],
B_[3][2][54],
B_[4][0][54],
B_[4][1][54],
B_[4][2][54],
B_[5][0][54],
B_[5][1][54],
B_[5][2][54],
B_[6][0][54],
B_[6][1][54],
B_[6][2][54],
B_[7][0][54],
B_[7][1][54],
B_[7][2][54],
B_[8][0][54],
B_[8][1][54],
B_[8][2][54],
B_[9][0][54],
B_[9][1][54],
B_[9][2][54],
B_[10][0][54],
B_[10][1][54],
B_[10][2][54],
B_[11][0][54],
B_[11][1][54],
B_[11][2][54],
B_[12][0][54],
B_[12][1][54],
B_[12][2][54],
B_[13][0][54],
B_[13][1][54],
B_[13][2][54],
B_[14][0][54],
B_[14][1][54],
B_[14][2][54],
B_[15][0][54],
B_[15][1][54],
B_[15][2][54],
B_[0][0][55],
B_[0][1][55],
B_[0][2][55],
B_[1][0][55],
B_[1][1][55],
B_[1][2][55],
B_[2][0][55],
B_[2][1][55],
B_[2][2][55],
B_[3][0][55],
B_[3][1][55],
B_[3][2][55],
B_[4][0][55],
B_[4][1][55],
B_[4][2][55],
B_[5][0][55],
B_[5][1][55],
B_[5][2][55],
B_[6][0][55],
B_[6][1][55],
B_[6][2][55],
B_[7][0][55],
B_[7][1][55],
B_[7][2][55],
B_[8][0][55],
B_[8][1][55],
B_[8][2][55],
B_[9][0][55],
B_[9][1][55],
B_[9][2][55],
B_[10][0][55],
B_[10][1][55],
B_[10][2][55],
B_[11][0][55],
B_[11][1][55],
B_[11][2][55],
B_[12][0][55],
B_[12][1][55],
B_[12][2][55],
B_[13][0][55],
B_[13][1][55],
B_[13][2][55],
B_[14][0][55],
B_[14][1][55],
B_[14][2][55],
B_[15][0][55],
B_[15][1][55],
B_[15][2][55],
B_[0][0][56],
B_[0][1][56],
B_[0][2][56],
B_[1][0][56],
B_[1][1][56],
B_[1][2][56],
B_[2][0][56],
B_[2][1][56],
B_[2][2][56],
B_[3][0][56],
B_[3][1][56],
B_[3][2][56],
B_[4][0][56],
B_[4][1][56],
B_[4][2][56],
B_[5][0][56],
B_[5][1][56],
B_[5][2][56],
B_[6][0][56],
B_[6][1][56],
B_[6][2][56],
B_[7][0][56],
B_[7][1][56],
B_[7][2][56],
B_[8][0][56],
B_[8][1][56],
B_[8][2][56],
B_[9][0][56],
B_[9][1][56],
B_[9][2][56],
B_[10][0][56],
B_[10][1][56],
B_[10][2][56],
B_[11][0][56],
B_[11][1][56],
B_[11][2][56],
B_[12][0][56],
B_[12][1][56],
B_[12][2][56],
B_[13][0][56],
B_[13][1][56],
B_[13][2][56],
B_[14][0][56],
B_[14][1][56],
B_[14][2][56],
B_[15][0][56],
B_[15][1][56],
B_[15][2][56],
B_[0][0][57],
B_[0][1][57],
B_[0][2][57],
B_[1][0][57],
B_[1][1][57],
B_[1][2][57],
B_[2][0][57],
B_[2][1][57],
B_[2][2][57],
B_[3][0][57],
B_[3][1][57],
B_[3][2][57],
B_[4][0][57],
B_[4][1][57],
B_[4][2][57],
B_[5][0][57],
B_[5][1][57],
B_[5][2][57],
B_[6][0][57],
B_[6][1][57],
B_[6][2][57],
B_[7][0][57],
B_[7][1][57],
B_[7][2][57],
B_[8][0][57],
B_[8][1][57],
B_[8][2][57],
B_[9][0][57],
B_[9][1][57],
B_[9][2][57],
B_[10][0][57],
B_[10][1][57],
B_[10][2][57],
B_[11][0][57],
B_[11][1][57],
B_[11][2][57],
B_[12][0][57],
B_[12][1][57],
B_[12][2][57],
B_[13][0][57],
B_[13][1][57],
B_[13][2][57],
B_[14][0][57],
B_[14][1][57],
B_[14][2][57],
B_[15][0][57],
B_[15][1][57],
B_[15][2][57],
B_[0][0][58],
B_[0][1][58],
B_[0][2][58],
B_[1][0][58],
B_[1][1][58],
B_[1][2][58],
B_[2][0][58],
B_[2][1][58],
B_[2][2][58],
B_[3][0][58],
B_[3][1][58],
B_[3][2][58],
B_[4][0][58],
B_[4][1][58],
B_[4][2][58],
B_[5][0][58],
B_[5][1][58],
B_[5][2][58],
B_[6][0][58],
B_[6][1][58],
B_[6][2][58],
B_[7][0][58],
B_[7][1][58],
B_[7][2][58],
B_[8][0][58],
B_[8][1][58],
B_[8][2][58],
B_[9][0][58],
B_[9][1][58],
B_[9][2][58],
B_[10][0][58],
B_[10][1][58],
B_[10][2][58],
B_[11][0][58],
B_[11][1][58],
B_[11][2][58],
B_[12][0][58],
B_[12][1][58],
B_[12][2][58],
B_[13][0][58],
B_[13][1][58],
B_[13][2][58],
B_[14][0][58],
B_[14][1][58],
B_[14][2][58],
B_[15][0][58],
B_[15][1][58],
B_[15][2][58],
B_[0][0][59],
B_[0][1][59],
B_[0][2][59],
B_[1][0][59],
B_[1][1][59],
B_[1][2][59],
B_[2][0][59],
B_[2][1][59],
B_[2][2][59],
B_[3][0][59],
B_[3][1][59],
B_[3][2][59],
B_[4][0][59],
B_[4][1][59],
B_[4][2][59],
B_[5][0][59],
B_[5][1][59],
B_[5][2][59],
B_[6][0][59],
B_[6][1][59],
B_[6][2][59],
B_[7][0][59],
B_[7][1][59],
B_[7][2][59],
B_[8][0][59],
B_[8][1][59],
B_[8][2][59],
B_[9][0][59],
B_[9][1][59],
B_[9][2][59],
B_[10][0][59],
B_[10][1][59],
B_[10][2][59],
B_[11][0][59],
B_[11][1][59],
B_[11][2][59],
B_[12][0][59],
B_[12][1][59],
B_[12][2][59],
B_[13][0][59],
B_[13][1][59],
B_[13][2][59],
B_[14][0][59],
B_[14][1][59],
B_[14][2][59],
B_[15][0][59],
B_[15][1][59],
B_[15][2][59],
B_[0][0][60],
B_[0][1][60],
B_[0][2][60],
B_[1][0][60],
B_[1][1][60],
B_[1][2][60],
B_[2][0][60],
B_[2][1][60],
B_[2][2][60],
B_[3][0][60],
B_[3][1][60],
B_[3][2][60],
B_[4][0][60],
B_[4][1][60],
B_[4][2][60],
B_[5][0][60],
B_[5][1][60],
B_[5][2][60],
B_[6][0][60],
B_[6][1][60],
B_[6][2][60],
B_[7][0][60],
B_[7][1][60],
B_[7][2][60],
B_[8][0][60],
B_[8][1][60],
B_[8][2][60],
B_[9][0][60],
B_[9][1][60],
B_[9][2][60],
B_[10][0][60],
B_[10][1][60],
B_[10][2][60],
B_[11][0][60],
B_[11][1][60],
B_[11][2][60],
B_[12][0][60],
B_[12][1][60],
B_[12][2][60],
B_[13][0][60],
B_[13][1][60],
B_[13][2][60],
B_[14][0][60],
B_[14][1][60],
B_[14][2][60],
B_[15][0][60],
B_[15][1][60],
B_[15][2][60],
B_[0][0][61],
B_[0][1][61],
B_[0][2][61],
B_[1][0][61],
B_[1][1][61],
B_[1][2][61],
B_[2][0][61],
B_[2][1][61],
B_[2][2][61],
B_[3][0][61],
B_[3][1][61],
B_[3][2][61],
B_[4][0][61],
B_[4][1][61],
B_[4][2][61],
B_[5][0][61],
B_[5][1][61],
B_[5][2][61],
B_[6][0][61],
B_[6][1][61],
B_[6][2][61],
B_[7][0][61],
B_[7][1][61],
B_[7][2][61],
B_[8][0][61],
B_[8][1][61],
B_[8][2][61],
B_[9][0][61],
B_[9][1][61],
B_[9][2][61],
B_[10][0][61],
B_[10][1][61],
B_[10][2][61],
B_[11][0][61],
B_[11][1][61],
B_[11][2][61],
B_[12][0][61],
B_[12][1][61],
B_[12][2][61],
B_[13][0][61],
B_[13][1][61],
B_[13][2][61],
B_[14][0][61],
B_[14][1][61],
B_[14][2][61],
B_[15][0][61],
B_[15][1][61],
B_[15][2][61],
B_[0][0][62],
B_[0][1][62],
B_[0][2][62],
B_[1][0][62],
B_[1][1][62],
B_[1][2][62],
B_[2][0][62],
B_[2][1][62],
B_[2][2][62],
B_[3][0][62],
B_[3][1][62],
B_[3][2][62],
B_[4][0][62],
B_[4][1][62],
B_[4][2][62],
B_[5][0][62],
B_[5][1][62],
B_[5][2][62],
B_[6][0][62],
B_[6][1][62],
B_[6][2][62],
B_[7][0][62],
B_[7][1][62],
B_[7][2][62],
B_[8][0][62],
B_[8][1][62],
B_[8][2][62],
B_[9][0][62],
B_[9][1][62],
B_[9][2][62],
B_[10][0][62],
B_[10][1][62],
B_[10][2][62],
B_[11][0][62],
B_[11][1][62],
B_[11][2][62],
B_[12][0][62],
B_[12][1][62],
B_[12][2][62],
B_[13][0][62],
B_[13][1][62],
B_[13][2][62],
B_[14][0][62],
B_[14][1][62],
B_[14][2][62],
B_[15][0][62],
B_[15][1][62],
B_[15][2][62],
B_[0][0][63],
B_[0][1][63],
B_[0][2][63],
B_[1][0][63],
B_[1][1][63],
B_[1][2][63],
B_[2][0][63],
B_[2][1][63],
B_[2][2][63],
B_[3][0][63],
B_[3][1][63],
B_[3][2][63],
B_[4][0][63],
B_[4][1][63],
B_[4][2][63],
B_[5][0][63],
B_[5][1][63],
B_[5][2][63],
B_[6][0][63],
B_[6][1][63],
B_[6][2][63],
B_[7][0][63],
B_[7][1][63],
B_[7][2][63],
B_[8][0][63],
B_[8][1][63],
B_[8][2][63],
B_[9][0][63],
B_[9][1][63],
B_[9][2][63],
B_[10][0][63],
B_[10][1][63],
B_[10][2][63],
B_[11][0][63],
B_[11][1][63],
B_[11][2][63],
B_[12][0][63],
B_[12][1][63],
B_[12][2][63],
B_[13][0][63],
B_[13][1][63],
B_[13][2][63],
B_[14][0][63],
B_[14][1][63],
B_[14][2][63],
B_[15][0][63],
B_[15][1][63],
B_[15][2][63],
B_[0][0][64],
B_[0][1][64],
B_[0][2][64],
B_[1][0][64],
B_[1][1][64],
B_[1][2][64],
B_[2][0][64],
B_[2][1][64],
B_[2][2][64],
B_[3][0][64],
B_[3][1][64],
B_[3][2][64],
B_[4][0][64],
B_[4][1][64],
B_[4][2][64],
B_[5][0][64],
B_[5][1][64],
B_[5][2][64],
B_[6][0][64],
B_[6][1][64],
B_[6][2][64],
B_[7][0][64],
B_[7][1][64],
B_[7][2][64],
B_[8][0][64],
B_[8][1][64],
B_[8][2][64],
B_[9][0][64],
B_[9][1][64],
B_[9][2][64],
B_[10][0][64],
B_[10][1][64],
B_[10][2][64],
B_[11][0][64],
B_[11][1][64],
B_[11][2][64],
B_[12][0][64],
B_[12][1][64],
B_[12][2][64],
B_[13][0][64],
B_[13][1][64],
B_[13][2][64],
B_[14][0][64],
B_[14][1][64],
B_[14][2][64],
B_[15][0][64],
B_[15][1][64],
B_[15][2][64],
B_[0][0][65],
B_[0][1][65],
B_[0][2][65],
B_[1][0][65],
B_[1][1][65],
B_[1][2][65],
B_[2][0][65],
B_[2][1][65],
B_[2][2][65],
B_[3][0][65],
B_[3][1][65],
B_[3][2][65],
B_[4][0][65],
B_[4][1][65],
B_[4][2][65],
B_[5][0][65],
B_[5][1][65],
B_[5][2][65],
B_[6][0][65],
B_[6][1][65],
B_[6][2][65],
B_[7][0][65],
B_[7][1][65],
B_[7][2][65],
B_[8][0][65],
B_[8][1][65],
B_[8][2][65],
B_[9][0][65],
B_[9][1][65],
B_[9][2][65],
B_[10][0][65],
B_[10][1][65],
B_[10][2][65],
B_[11][0][65],
B_[11][1][65],
B_[11][2][65],
B_[12][0][65],
B_[12][1][65],
B_[12][2][65],
B_[13][0][65],
B_[13][1][65],
B_[13][2][65],
B_[14][0][65],
B_[14][1][65],
B_[14][2][65],
B_[15][0][65],
B_[15][1][65],
B_[15][2][65],
B_[0][0][66],
B_[0][1][66],
B_[0][2][66],
B_[1][0][66],
B_[1][1][66],
B_[1][2][66],
B_[2][0][66],
B_[2][1][66],
B_[2][2][66],
B_[3][0][66],
B_[3][1][66],
B_[3][2][66],
B_[4][0][66],
B_[4][1][66],
B_[4][2][66],
B_[5][0][66],
B_[5][1][66],
B_[5][2][66],
B_[6][0][66],
B_[6][1][66],
B_[6][2][66],
B_[7][0][66],
B_[7][1][66],
B_[7][2][66],
B_[8][0][66],
B_[8][1][66],
B_[8][2][66],
B_[9][0][66],
B_[9][1][66],
B_[9][2][66],
B_[10][0][66],
B_[10][1][66],
B_[10][2][66],
B_[11][0][66],
B_[11][1][66],
B_[11][2][66],
B_[12][0][66],
B_[12][1][66],
B_[12][2][66],
B_[13][0][66],
B_[13][1][66],
B_[13][2][66],
B_[14][0][66],
B_[14][1][66],
B_[14][2][66],
B_[15][0][66],
B_[15][1][66],
B_[15][2][66],
B_[0][0][67],
B_[0][1][67],
B_[0][2][67],
B_[1][0][67],
B_[1][1][67],
B_[1][2][67],
B_[2][0][67],
B_[2][1][67],
B_[2][2][67],
B_[3][0][67],
B_[3][1][67],
B_[3][2][67],
B_[4][0][67],
B_[4][1][67],
B_[4][2][67],
B_[5][0][67],
B_[5][1][67],
B_[5][2][67],
B_[6][0][67],
B_[6][1][67],
B_[6][2][67],
B_[7][0][67],
B_[7][1][67],
B_[7][2][67],
B_[8][0][67],
B_[8][1][67],
B_[8][2][67],
B_[9][0][67],
B_[9][1][67],
B_[9][2][67],
B_[10][0][67],
B_[10][1][67],
B_[10][2][67],
B_[11][0][67],
B_[11][1][67],
B_[11][2][67],
B_[12][0][67],
B_[12][1][67],
B_[12][2][67],
B_[13][0][67],
B_[13][1][67],
B_[13][2][67],
B_[14][0][67],
B_[14][1][67],
B_[14][2][67],
B_[15][0][67],
B_[15][1][67],
B_[15][2][67],
B_[0][0][68],
B_[0][1][68],
B_[0][2][68],
B_[1][0][68],
B_[1][1][68],
B_[1][2][68],
B_[2][0][68],
B_[2][1][68],
B_[2][2][68],
B_[3][0][68],
B_[3][1][68],
B_[3][2][68],
B_[4][0][68],
B_[4][1][68],
B_[4][2][68],
B_[5][0][68],
B_[5][1][68],
B_[5][2][68],
B_[6][0][68],
B_[6][1][68],
B_[6][2][68],
B_[7][0][68],
B_[7][1][68],
B_[7][2][68],
B_[8][0][68],
B_[8][1][68],
B_[8][2][68],
B_[9][0][68],
B_[9][1][68],
B_[9][2][68],
B_[10][0][68],
B_[10][1][68],
B_[10][2][68],
B_[11][0][68],
B_[11][1][68],
B_[11][2][68],
B_[12][0][68],
B_[12][1][68],
B_[12][2][68],
B_[13][0][68],
B_[13][1][68],
B_[13][2][68],
B_[14][0][68],
B_[14][1][68],
B_[14][2][68],
B_[15][0][68],
B_[15][1][68],
B_[15][2][68],
B_[0][0][69],
B_[0][1][69],
B_[0][2][69],
B_[1][0][69],
B_[1][1][69],
B_[1][2][69],
B_[2][0][69],
B_[2][1][69],
B_[2][2][69],
B_[3][0][69],
B_[3][1][69],
B_[3][2][69],
B_[4][0][69],
B_[4][1][69],
B_[4][2][69],
B_[5][0][69],
B_[5][1][69],
B_[5][2][69],
B_[6][0][69],
B_[6][1][69],
B_[6][2][69],
B_[7][0][69],
B_[7][1][69],
B_[7][2][69],
B_[8][0][69],
B_[8][1][69],
B_[8][2][69],
B_[9][0][69],
B_[9][1][69],
B_[9][2][69],
B_[10][0][69],
B_[10][1][69],
B_[10][2][69],
B_[11][0][69],
B_[11][1][69],
B_[11][2][69],
B_[12][0][69],
B_[12][1][69],
B_[12][2][69],
B_[13][0][69],
B_[13][1][69],
B_[13][2][69],
B_[14][0][69],
B_[14][1][69],
B_[14][2][69],
B_[15][0][69],
B_[15][1][69],
B_[15][2][69],
B_[0][0][70],
B_[0][1][70],
B_[0][2][70],
B_[1][0][70],
B_[1][1][70],
B_[1][2][70],
B_[2][0][70],
B_[2][1][70],
B_[2][2][70],
B_[3][0][70],
B_[3][1][70],
B_[3][2][70],
B_[4][0][70],
B_[4][1][70],
B_[4][2][70],
B_[5][0][70],
B_[5][1][70],
B_[5][2][70],
B_[6][0][70],
B_[6][1][70],
B_[6][2][70],
B_[7][0][70],
B_[7][1][70],
B_[7][2][70],
B_[8][0][70],
B_[8][1][70],
B_[8][2][70],
B_[9][0][70],
B_[9][1][70],
B_[9][2][70],
B_[10][0][70],
B_[10][1][70],
B_[10][2][70],
B_[11][0][70],
B_[11][1][70],
B_[11][2][70],
B_[12][0][70],
B_[12][1][70],
B_[12][2][70],
B_[13][0][70],
B_[13][1][70],
B_[13][2][70],
B_[14][0][70],
B_[14][1][70],
B_[14][2][70],
B_[15][0][70],
B_[15][1][70],
B_[15][2][70],
B_[0][0][71],
B_[0][1][71],
B_[0][2][71],
B_[1][0][71],
B_[1][1][71],
B_[1][2][71],
B_[2][0][71],
B_[2][1][71],
B_[2][2][71],
B_[3][0][71],
B_[3][1][71],
B_[3][2][71],
B_[4][0][71],
B_[4][1][71],
B_[4][2][71],
B_[5][0][71],
B_[5][1][71],
B_[5][2][71],
B_[6][0][71],
B_[6][1][71],
B_[6][2][71],
B_[7][0][71],
B_[7][1][71],
B_[7][2][71],
B_[8][0][71],
B_[8][1][71],
B_[8][2][71],
B_[9][0][71],
B_[9][1][71],
B_[9][2][71],
B_[10][0][71],
B_[10][1][71],
B_[10][2][71],
B_[11][0][71],
B_[11][1][71],
B_[11][2][71],
B_[12][0][71],
B_[12][1][71],
B_[12][2][71],
B_[13][0][71],
B_[13][1][71],
B_[13][2][71],
B_[14][0][71],
B_[14][1][71],
B_[14][2][71],
B_[15][0][71],
B_[15][1][71],
B_[15][2][71],
B_[0][0][72],
B_[0][1][72],
B_[0][2][72],
B_[1][0][72],
B_[1][1][72],
B_[1][2][72],
B_[2][0][72],
B_[2][1][72],
B_[2][2][72],
B_[3][0][72],
B_[3][1][72],
B_[3][2][72],
B_[4][0][72],
B_[4][1][72],
B_[4][2][72],
B_[5][0][72],
B_[5][1][72],
B_[5][2][72],
B_[6][0][72],
B_[6][1][72],
B_[6][2][72],
B_[7][0][72],
B_[7][1][72],
B_[7][2][72],
B_[8][0][72],
B_[8][1][72],
B_[8][2][72],
B_[9][0][72],
B_[9][1][72],
B_[9][2][72],
B_[10][0][72],
B_[10][1][72],
B_[10][2][72],
B_[11][0][72],
B_[11][1][72],
B_[11][2][72],
B_[12][0][72],
B_[12][1][72],
B_[12][2][72],
B_[13][0][72],
B_[13][1][72],
B_[13][2][72],
B_[14][0][72],
B_[14][1][72],
B_[14][2][72],
B_[15][0][72],
B_[15][1][72],
B_[15][2][72],
B_[0][0][73],
B_[0][1][73],
B_[0][2][73],
B_[1][0][73],
B_[1][1][73],
B_[1][2][73],
B_[2][0][73],
B_[2][1][73],
B_[2][2][73],
B_[3][0][73],
B_[3][1][73],
B_[3][2][73],
B_[4][0][73],
B_[4][1][73],
B_[4][2][73],
B_[5][0][73],
B_[5][1][73],
B_[5][2][73],
B_[6][0][73],
B_[6][1][73],
B_[6][2][73],
B_[7][0][73],
B_[7][1][73],
B_[7][2][73],
B_[8][0][73],
B_[8][1][73],
B_[8][2][73],
B_[9][0][73],
B_[9][1][73],
B_[9][2][73],
B_[10][0][73],
B_[10][1][73],
B_[10][2][73],
B_[11][0][73],
B_[11][1][73],
B_[11][2][73],
B_[12][0][73],
B_[12][1][73],
B_[12][2][73],
B_[13][0][73],
B_[13][1][73],
B_[13][2][73],
B_[14][0][73],
B_[14][1][73],
B_[14][2][73],
B_[15][0][73],
B_[15][1][73],
B_[15][2][73],
B_[0][0][74],
B_[0][1][74],
B_[0][2][74],
B_[1][0][74],
B_[1][1][74],
B_[1][2][74],
B_[2][0][74],
B_[2][1][74],
B_[2][2][74],
B_[3][0][74],
B_[3][1][74],
B_[3][2][74],
B_[4][0][74],
B_[4][1][74],
B_[4][2][74],
B_[5][0][74],
B_[5][1][74],
B_[5][2][74],
B_[6][0][74],
B_[6][1][74],
B_[6][2][74],
B_[7][0][74],
B_[7][1][74],
B_[7][2][74],
B_[8][0][74],
B_[8][1][74],
B_[8][2][74],
B_[9][0][74],
B_[9][1][74],
B_[9][2][74],
B_[10][0][74],
B_[10][1][74],
B_[10][2][74],
B_[11][0][74],
B_[11][1][74],
B_[11][2][74],
B_[12][0][74],
B_[12][1][74],
B_[12][2][74],
B_[13][0][74],
B_[13][1][74],
B_[13][2][74],
B_[14][0][74],
B_[14][1][74],
B_[14][2][74],
B_[15][0][74],
B_[15][1][74],
B_[15][2][74],
B_[0][0][75],
B_[0][1][75],
B_[0][2][75],
B_[1][0][75],
B_[1][1][75],
B_[1][2][75],
B_[2][0][75],
B_[2][1][75],
B_[2][2][75],
B_[3][0][75],
B_[3][1][75],
B_[3][2][75],
B_[4][0][75],
B_[4][1][75],
B_[4][2][75],
B_[5][0][75],
B_[5][1][75],
B_[5][2][75],
B_[6][0][75],
B_[6][1][75],
B_[6][2][75],
B_[7][0][75],
B_[7][1][75],
B_[7][2][75],
B_[8][0][75],
B_[8][1][75],
B_[8][2][75],
B_[9][0][75],
B_[9][1][75],
B_[9][2][75],
B_[10][0][75],
B_[10][1][75],
B_[10][2][75],
B_[11][0][75],
B_[11][1][75],
B_[11][2][75],
B_[12][0][75],
B_[12][1][75],
B_[12][2][75],
B_[13][0][75],
B_[13][1][75],
B_[13][2][75],
B_[14][0][75],
B_[14][1][75],
B_[14][2][75],
B_[15][0][75],
B_[15][1][75],
B_[15][2][75],
B_[0][0][76],
B_[0][1][76],
B_[0][2][76],
B_[1][0][76],
B_[1][1][76],
B_[1][2][76],
B_[2][0][76],
B_[2][1][76],
B_[2][2][76],
B_[3][0][76],
B_[3][1][76],
B_[3][2][76],
B_[4][0][76],
B_[4][1][76],
B_[4][2][76],
B_[5][0][76],
B_[5][1][76],
B_[5][2][76],
B_[6][0][76],
B_[6][1][76],
B_[6][2][76],
B_[7][0][76],
B_[7][1][76],
B_[7][2][76],
B_[8][0][76],
B_[8][1][76],
B_[8][2][76],
B_[9][0][76],
B_[9][1][76],
B_[9][2][76],
B_[10][0][76],
B_[10][1][76],
B_[10][2][76],
B_[11][0][76],
B_[11][1][76],
B_[11][2][76],
B_[12][0][76],
B_[12][1][76],
B_[12][2][76],
B_[13][0][76],
B_[13][1][76],
B_[13][2][76],
B_[14][0][76],
B_[14][1][76],
B_[14][2][76],
B_[15][0][76],
B_[15][1][76],
B_[15][2][76],
B_[0][0][77],
B_[0][1][77],
B_[0][2][77],
B_[1][0][77],
B_[1][1][77],
B_[1][2][77],
B_[2][0][77],
B_[2][1][77],
B_[2][2][77],
B_[3][0][77],
B_[3][1][77],
B_[3][2][77],
B_[4][0][77],
B_[4][1][77],
B_[4][2][77],
B_[5][0][77],
B_[5][1][77],
B_[5][2][77],
B_[6][0][77],
B_[6][1][77],
B_[6][2][77],
B_[7][0][77],
B_[7][1][77],
B_[7][2][77],
B_[8][0][77],
B_[8][1][77],
B_[8][2][77],
B_[9][0][77],
B_[9][1][77],
B_[9][2][77],
B_[10][0][77],
B_[10][1][77],
B_[10][2][77],
B_[11][0][77],
B_[11][1][77],
B_[11][2][77],
B_[12][0][77],
B_[12][1][77],
B_[12][2][77],
B_[13][0][77],
B_[13][1][77],
B_[13][2][77],
B_[14][0][77],
B_[14][1][77],
B_[14][2][77],
B_[15][0][77],
B_[15][1][77],
B_[15][2][77],
B_[0][0][78],
B_[0][1][78],
B_[0][2][78],
B_[1][0][78],
B_[1][1][78],
B_[1][2][78],
B_[2][0][78],
B_[2][1][78],
B_[2][2][78],
B_[3][0][78],
B_[3][1][78],
B_[3][2][78],
B_[4][0][78],
B_[4][1][78],
B_[4][2][78],
B_[5][0][78],
B_[5][1][78],
B_[5][2][78],
B_[6][0][78],
B_[6][1][78],
B_[6][2][78],
B_[7][0][78],
B_[7][1][78],
B_[7][2][78],
B_[8][0][78],
B_[8][1][78],
B_[8][2][78],
B_[9][0][78],
B_[9][1][78],
B_[9][2][78],
B_[10][0][78],
B_[10][1][78],
B_[10][2][78],
B_[11][0][78],
B_[11][1][78],
B_[11][2][78],
B_[12][0][78],
B_[12][1][78],
B_[12][2][78],
B_[13][0][78],
B_[13][1][78],
B_[13][2][78],
B_[14][0][78],
B_[14][1][78],
B_[14][2][78],
B_[15][0][78],
B_[15][1][78],
B_[15][2][78],
B_[0][0][79],
B_[0][1][79],
B_[0][2][79],
B_[1][0][79],
B_[1][1][79],
B_[1][2][79],
B_[2][0][79],
B_[2][1][79],
B_[2][2][79],
B_[3][0][79],
B_[3][1][79],
B_[3][2][79],
B_[4][0][79],
B_[4][1][79],
B_[4][2][79],
B_[5][0][79],
B_[5][1][79],
B_[5][2][79],
B_[6][0][79],
B_[6][1][79],
B_[6][2][79],
B_[7][0][79],
B_[7][1][79],
B_[7][2][79],
B_[8][0][79],
B_[8][1][79],
B_[8][2][79],
B_[9][0][79],
B_[9][1][79],
B_[9][2][79],
B_[10][0][79],
B_[10][1][79],
B_[10][2][79],
B_[11][0][79],
B_[11][1][79],
B_[11][2][79],
B_[12][0][79],
B_[12][1][79],
B_[12][2][79],
B_[13][0][79],
B_[13][1][79],
B_[13][2][79],
B_[14][0][79],
B_[14][1][79],
B_[14][2][79],
B_[15][0][79],
B_[15][1][79],
B_[15][2][79],
B_[0][0][80],
B_[0][1][80],
B_[0][2][80],
B_[1][0][80],
B_[1][1][80],
B_[1][2][80],
B_[2][0][80],
B_[2][1][80],
B_[2][2][80],
B_[3][0][80],
B_[3][1][80],
B_[3][2][80],
B_[4][0][80],
B_[4][1][80],
B_[4][2][80],
B_[5][0][80],
B_[5][1][80],
B_[5][2][80],
B_[6][0][80],
B_[6][1][80],
B_[6][2][80],
B_[7][0][80],
B_[7][1][80],
B_[7][2][80],
B_[8][0][80],
B_[8][1][80],
B_[8][2][80],
B_[9][0][80],
B_[9][1][80],
B_[9][2][80],
B_[10][0][80],
B_[10][1][80],
B_[10][2][80],
B_[11][0][80],
B_[11][1][80],
B_[11][2][80],
B_[12][0][80],
B_[12][1][80],
B_[12][2][80],
B_[13][0][80],
B_[13][1][80],
B_[13][2][80],
B_[14][0][80],
B_[14][1][80],
B_[14][2][80],
B_[15][0][80],
B_[15][1][80],
B_[15][2][80],
B_[0][0][81],
B_[0][1][81],
B_[0][2][81],
B_[1][0][81],
B_[1][1][81],
B_[1][2][81],
B_[2][0][81],
B_[2][1][81],
B_[2][2][81],
B_[3][0][81],
B_[3][1][81],
B_[3][2][81],
B_[4][0][81],
B_[4][1][81],
B_[4][2][81],
B_[5][0][81],
B_[5][1][81],
B_[5][2][81],
B_[6][0][81],
B_[6][1][81],
B_[6][2][81],
B_[7][0][81],
B_[7][1][81],
B_[7][2][81],
B_[8][0][81],
B_[8][1][81],
B_[8][2][81],
B_[9][0][81],
B_[9][1][81],
B_[9][2][81],
B_[10][0][81],
B_[10][1][81],
B_[10][2][81],
B_[11][0][81],
B_[11][1][81],
B_[11][2][81],
B_[12][0][81],
B_[12][1][81],
B_[12][2][81],
B_[13][0][81],
B_[13][1][81],
B_[13][2][81],
B_[14][0][81],
B_[14][1][81],
B_[14][2][81],
B_[15][0][81],
B_[15][1][81],
B_[15][2][81],
B_[0][0][82],
B_[0][1][82],
B_[0][2][82],
B_[1][0][82],
B_[1][1][82],
B_[1][2][82],
B_[2][0][82],
B_[2][1][82],
B_[2][2][82],
B_[3][0][82],
B_[3][1][82],
B_[3][2][82],
B_[4][0][82],
B_[4][1][82],
B_[4][2][82],
B_[5][0][82],
B_[5][1][82],
B_[5][2][82],
B_[6][0][82],
B_[6][1][82],
B_[6][2][82],
B_[7][0][82],
B_[7][1][82],
B_[7][2][82],
B_[8][0][82],
B_[8][1][82],
B_[8][2][82],
B_[9][0][82],
B_[9][1][82],
B_[9][2][82],
B_[10][0][82],
B_[10][1][82],
B_[10][2][82],
B_[11][0][82],
B_[11][1][82],
B_[11][2][82],
B_[12][0][82],
B_[12][1][82],
B_[12][2][82],
B_[13][0][82],
B_[13][1][82],
B_[13][2][82],
B_[14][0][82],
B_[14][1][82],
B_[14][2][82],
B_[15][0][82],
B_[15][1][82],
B_[15][2][82],
B_[0][0][83],
B_[0][1][83],
B_[0][2][83],
B_[1][0][83],
B_[1][1][83],
B_[1][2][83],
B_[2][0][83],
B_[2][1][83],
B_[2][2][83],
B_[3][0][83],
B_[3][1][83],
B_[3][2][83],
B_[4][0][83],
B_[4][1][83],
B_[4][2][83],
B_[5][0][83],
B_[5][1][83],
B_[5][2][83],
B_[6][0][83],
B_[6][1][83],
B_[6][2][83],
B_[7][0][83],
B_[7][1][83],
B_[7][2][83],
B_[8][0][83],
B_[8][1][83],
B_[8][2][83],
B_[9][0][83],
B_[9][1][83],
B_[9][2][83],
B_[10][0][83],
B_[10][1][83],
B_[10][2][83],
B_[11][0][83],
B_[11][1][83],
B_[11][2][83],
B_[12][0][83],
B_[12][1][83],
B_[12][2][83],
B_[13][0][83],
B_[13][1][83],
B_[13][2][83],
B_[14][0][83],
B_[14][1][83],
B_[14][2][83],
B_[15][0][83],
B_[15][1][83],
B_[15][2][83],
B_[0][0][84],
B_[0][1][84],
B_[0][2][84],
B_[1][0][84],
B_[1][1][84],
B_[1][2][84],
B_[2][0][84],
B_[2][1][84],
B_[2][2][84],
B_[3][0][84],
B_[3][1][84],
B_[3][2][84],
B_[4][0][84],
B_[4][1][84],
B_[4][2][84],
B_[5][0][84],
B_[5][1][84],
B_[5][2][84],
B_[6][0][84],
B_[6][1][84],
B_[6][2][84],
B_[7][0][84],
B_[7][1][84],
B_[7][2][84],
B_[8][0][84],
B_[8][1][84],
B_[8][2][84],
B_[9][0][84],
B_[9][1][84],
B_[9][2][84],
B_[10][0][84],
B_[10][1][84],
B_[10][2][84],
B_[11][0][84],
B_[11][1][84],
B_[11][2][84],
B_[12][0][84],
B_[12][1][84],
B_[12][2][84],
B_[13][0][84],
B_[13][1][84],
B_[13][2][84],
B_[14][0][84],
B_[14][1][84],
B_[14][2][84],
B_[15][0][84],
B_[15][1][84],
B_[15][2][84],
B_[0][0][85],
B_[0][1][85],
B_[0][2][85],
B_[1][0][85],
B_[1][1][85],
B_[1][2][85],
B_[2][0][85],
B_[2][1][85],
B_[2][2][85],
B_[3][0][85],
B_[3][1][85],
B_[3][2][85],
B_[4][0][85],
B_[4][1][85],
B_[4][2][85],
B_[5][0][85],
B_[5][1][85],
B_[5][2][85],
B_[6][0][85],
B_[6][1][85],
B_[6][2][85],
B_[7][0][85],
B_[7][1][85],
B_[7][2][85],
B_[8][0][85],
B_[8][1][85],
B_[8][2][85],
B_[9][0][85],
B_[9][1][85],
B_[9][2][85],
B_[10][0][85],
B_[10][1][85],
B_[10][2][85],
B_[11][0][85],
B_[11][1][85],
B_[11][2][85],
B_[12][0][85],
B_[12][1][85],
B_[12][2][85],
B_[13][0][85],
B_[13][1][85],
B_[13][2][85],
B_[14][0][85],
B_[14][1][85],
B_[14][2][85],
B_[15][0][85],
B_[15][1][85],
B_[15][2][85],
B_[0][0][86],
B_[0][1][86],
B_[0][2][86],
B_[1][0][86],
B_[1][1][86],
B_[1][2][86],
B_[2][0][86],
B_[2][1][86],
B_[2][2][86],
B_[3][0][86],
B_[3][1][86],
B_[3][2][86],
B_[4][0][86],
B_[4][1][86],
B_[4][2][86],
B_[5][0][86],
B_[5][1][86],
B_[5][2][86],
B_[6][0][86],
B_[6][1][86],
B_[6][2][86],
B_[7][0][86],
B_[7][1][86],
B_[7][2][86],
B_[8][0][86],
B_[8][1][86],
B_[8][2][86],
B_[9][0][86],
B_[9][1][86],
B_[9][2][86],
B_[10][0][86],
B_[10][1][86],
B_[10][2][86],
B_[11][0][86],
B_[11][1][86],
B_[11][2][86],
B_[12][0][86],
B_[12][1][86],
B_[12][2][86],
B_[13][0][86],
B_[13][1][86],
B_[13][2][86],
B_[14][0][86],
B_[14][1][86],
B_[14][2][86],
B_[15][0][86],
B_[15][1][86],
B_[15][2][86],
B_[0][0][87],
B_[0][1][87],
B_[0][2][87],
B_[1][0][87],
B_[1][1][87],
B_[1][2][87],
B_[2][0][87],
B_[2][1][87],
B_[2][2][87],
B_[3][0][87],
B_[3][1][87],
B_[3][2][87],
B_[4][0][87],
B_[4][1][87],
B_[4][2][87],
B_[5][0][87],
B_[5][1][87],
B_[5][2][87],
B_[6][0][87],
B_[6][1][87],
B_[6][2][87],
B_[7][0][87],
B_[7][1][87],
B_[7][2][87],
B_[8][0][87],
B_[8][1][87],
B_[8][2][87],
B_[9][0][87],
B_[9][1][87],
B_[9][2][87],
B_[10][0][87],
B_[10][1][87],
B_[10][2][87],
B_[11][0][87],
B_[11][1][87],
B_[11][2][87],
B_[12][0][87],
B_[12][1][87],
B_[12][2][87],
B_[13][0][87],
B_[13][1][87],
B_[13][2][87],
B_[14][0][87],
B_[14][1][87],
B_[14][2][87],
B_[15][0][87],
B_[15][1][87],
B_[15][2][87],
B_[0][0][88],
B_[0][1][88],
B_[0][2][88],
B_[1][0][88],
B_[1][1][88],
B_[1][2][88],
B_[2][0][88],
B_[2][1][88],
B_[2][2][88],
B_[3][0][88],
B_[3][1][88],
B_[3][2][88],
B_[4][0][88],
B_[4][1][88],
B_[4][2][88],
B_[5][0][88],
B_[5][1][88],
B_[5][2][88],
B_[6][0][88],
B_[6][1][88],
B_[6][2][88],
B_[7][0][88],
B_[7][1][88],
B_[7][2][88],
B_[8][0][88],
B_[8][1][88],
B_[8][2][88],
B_[9][0][88],
B_[9][1][88],
B_[9][2][88],
B_[10][0][88],
B_[10][1][88],
B_[10][2][88],
B_[11][0][88],
B_[11][1][88],
B_[11][2][88],
B_[12][0][88],
B_[12][1][88],
B_[12][2][88],
B_[13][0][88],
B_[13][1][88],
B_[13][2][88],
B_[14][0][88],
B_[14][1][88],
B_[14][2][88],
B_[15][0][88],
B_[15][1][88],
B_[15][2][88],
B_[0][0][89],
B_[0][1][89],
B_[0][2][89],
B_[1][0][89],
B_[1][1][89],
B_[1][2][89],
B_[2][0][89],
B_[2][1][89],
B_[2][2][89],
B_[3][0][89],
B_[3][1][89],
B_[3][2][89],
B_[4][0][89],
B_[4][1][89],
B_[4][2][89],
B_[5][0][89],
B_[5][1][89],
B_[5][2][89],
B_[6][0][89],
B_[6][1][89],
B_[6][2][89],
B_[7][0][89],
B_[7][1][89],
B_[7][2][89],
B_[8][0][89],
B_[8][1][89],
B_[8][2][89],
B_[9][0][89],
B_[9][1][89],
B_[9][2][89],
B_[10][0][89],
B_[10][1][89],
B_[10][2][89],
B_[11][0][89],
B_[11][1][89],
B_[11][2][89],
B_[12][0][89],
B_[12][1][89],
B_[12][2][89],
B_[13][0][89],
B_[13][1][89],
B_[13][2][89],
B_[14][0][89],
B_[14][1][89],
B_[14][2][89],
B_[15][0][89],
B_[15][1][89],
B_[15][2][89],
B_[0][0][90],
B_[0][1][90],
B_[0][2][90],
B_[1][0][90],
B_[1][1][90],
B_[1][2][90],
B_[2][0][90],
B_[2][1][90],
B_[2][2][90],
B_[3][0][90],
B_[3][1][90],
B_[3][2][90],
B_[4][0][90],
B_[4][1][90],
B_[4][2][90],
B_[5][0][90],
B_[5][1][90],
B_[5][2][90],
B_[6][0][90],
B_[6][1][90],
B_[6][2][90],
B_[7][0][90],
B_[7][1][90],
B_[7][2][90],
B_[8][0][90],
B_[8][1][90],
B_[8][2][90],
B_[9][0][90],
B_[9][1][90],
B_[9][2][90],
B_[10][0][90],
B_[10][1][90],
B_[10][2][90],
B_[11][0][90],
B_[11][1][90],
B_[11][2][90],
B_[12][0][90],
B_[12][1][90],
B_[12][2][90],
B_[13][0][90],
B_[13][1][90],
B_[13][2][90],
B_[14][0][90],
B_[14][1][90],
B_[14][2][90],
B_[15][0][90],
B_[15][1][90],
B_[15][2][90],
B_[0][0][91],
B_[0][1][91],
B_[0][2][91],
B_[1][0][91],
B_[1][1][91],
B_[1][2][91],
B_[2][0][91],
B_[2][1][91],
B_[2][2][91],
B_[3][0][91],
B_[3][1][91],
B_[3][2][91],
B_[4][0][91],
B_[4][1][91],
B_[4][2][91],
B_[5][0][91],
B_[5][1][91],
B_[5][2][91],
B_[6][0][91],
B_[6][1][91],
B_[6][2][91],
B_[7][0][91],
B_[7][1][91],
B_[7][2][91],
B_[8][0][91],
B_[8][1][91],
B_[8][2][91],
B_[9][0][91],
B_[9][1][91],
B_[9][2][91],
B_[10][0][91],
B_[10][1][91],
B_[10][2][91],
B_[11][0][91],
B_[11][1][91],
B_[11][2][91],
B_[12][0][91],
B_[12][1][91],
B_[12][2][91],
B_[13][0][91],
B_[13][1][91],
B_[13][2][91],
B_[14][0][91],
B_[14][1][91],
B_[14][2][91],
B_[15][0][91],
B_[15][1][91],
B_[15][2][91],
B_[0][0][92],
B_[0][1][92],
B_[0][2][92],
B_[1][0][92],
B_[1][1][92],
B_[1][2][92],
B_[2][0][92],
B_[2][1][92],
B_[2][2][92],
B_[3][0][92],
B_[3][1][92],
B_[3][2][92],
B_[4][0][92],
B_[4][1][92],
B_[4][2][92],
B_[5][0][92],
B_[5][1][92],
B_[5][2][92],
B_[6][0][92],
B_[6][1][92],
B_[6][2][92],
B_[7][0][92],
B_[7][1][92],
B_[7][2][92],
B_[8][0][92],
B_[8][1][92],
B_[8][2][92],
B_[9][0][92],
B_[9][1][92],
B_[9][2][92],
B_[10][0][92],
B_[10][1][92],
B_[10][2][92],
B_[11][0][92],
B_[11][1][92],
B_[11][2][92],
B_[12][0][92],
B_[12][1][92],
B_[12][2][92],
B_[13][0][92],
B_[13][1][92],
B_[13][2][92],
B_[14][0][92],
B_[14][1][92],
B_[14][2][92],
B_[15][0][92],
B_[15][1][92],
B_[15][2][92],
B_[0][0][93],
B_[0][1][93],
B_[0][2][93],
B_[1][0][93],
B_[1][1][93],
B_[1][2][93],
B_[2][0][93],
B_[2][1][93],
B_[2][2][93],
B_[3][0][93],
B_[3][1][93],
B_[3][2][93],
B_[4][0][93],
B_[4][1][93],
B_[4][2][93],
B_[5][0][93],
B_[5][1][93],
B_[5][2][93],
B_[6][0][93],
B_[6][1][93],
B_[6][2][93],
B_[7][0][93],
B_[7][1][93],
B_[7][2][93],
B_[8][0][93],
B_[8][1][93],
B_[8][2][93],
B_[9][0][93],
B_[9][1][93],
B_[9][2][93],
B_[10][0][93],
B_[10][1][93],
B_[10][2][93],
B_[11][0][93],
B_[11][1][93],
B_[11][2][93],
B_[12][0][93],
B_[12][1][93],
B_[12][2][93],
B_[13][0][93],
B_[13][1][93],
B_[13][2][93],
B_[14][0][93],
B_[14][1][93],
B_[14][2][93],
B_[15][0][93],
B_[15][1][93],
B_[15][2][93],
B_[0][0][94],
B_[0][1][94],
B_[0][2][94],
B_[1][0][94],
B_[1][1][94],
B_[1][2][94],
B_[2][0][94],
B_[2][1][94],
B_[2][2][94],
B_[3][0][94],
B_[3][1][94],
B_[3][2][94],
B_[4][0][94],
B_[4][1][94],
B_[4][2][94],
B_[5][0][94],
B_[5][1][94],
B_[5][2][94],
B_[6][0][94],
B_[6][1][94],
B_[6][2][94],
B_[7][0][94],
B_[7][1][94],
B_[7][2][94],
B_[8][0][94],
B_[8][1][94],
B_[8][2][94],
B_[9][0][94],
B_[9][1][94],
B_[9][2][94],
B_[10][0][94],
B_[10][1][94],
B_[10][2][94],
B_[11][0][94],
B_[11][1][94],
B_[11][2][94],
B_[12][0][94],
B_[12][1][94],
B_[12][2][94],
B_[13][0][94],
B_[13][1][94],
B_[13][2][94],
B_[14][0][94],
B_[14][1][94],
B_[14][2][94],
B_[15][0][94],
B_[15][1][94],
B_[15][2][94],
B_[0][0][95],
B_[0][1][95],
B_[0][2][95],
B_[1][0][95],
B_[1][1][95],
B_[1][2][95],
B_[2][0][95],
B_[2][1][95],
B_[2][2][95],
B_[3][0][95],
B_[3][1][95],
B_[3][2][95],
B_[4][0][95],
B_[4][1][95],
B_[4][2][95],
B_[5][0][95],
B_[5][1][95],
B_[5][2][95],
B_[6][0][95],
B_[6][1][95],
B_[6][2][95],
B_[7][0][95],
B_[7][1][95],
B_[7][2][95],
B_[8][0][95],
B_[8][1][95],
B_[8][2][95],
B_[9][0][95],
B_[9][1][95],
B_[9][2][95],
B_[10][0][95],
B_[10][1][95],
B_[10][2][95],
B_[11][0][95],
B_[11][1][95],
B_[11][2][95],
B_[12][0][95],
B_[12][1][95],
B_[12][2][95],
B_[13][0][95],
B_[13][1][95],
B_[13][2][95],
B_[14][0][95],
B_[14][1][95],
B_[14][2][95],
B_[15][0][95],
B_[15][1][95],
B_[15][2][95],
B_[0][0][96],
B_[0][1][96],
B_[0][2][96],
B_[1][0][96],
B_[1][1][96],
B_[1][2][96],
B_[2][0][96],
B_[2][1][96],
B_[2][2][96],
B_[3][0][96],
B_[3][1][96],
B_[3][2][96],
B_[4][0][96],
B_[4][1][96],
B_[4][2][96],
B_[5][0][96],
B_[5][1][96],
B_[5][2][96],
B_[6][0][96],
B_[6][1][96],
B_[6][2][96],
B_[7][0][96],
B_[7][1][96],
B_[7][2][96],
B_[8][0][96],
B_[8][1][96],
B_[8][2][96],
B_[9][0][96],
B_[9][1][96],
B_[9][2][96],
B_[10][0][96],
B_[10][1][96],
B_[10][2][96],
B_[11][0][96],
B_[11][1][96],
B_[11][2][96],
B_[12][0][96],
B_[12][1][96],
B_[12][2][96],
B_[13][0][96],
B_[13][1][96],
B_[13][2][96],
B_[14][0][96],
B_[14][1][96],
B_[14][2][96],
B_[15][0][96],
B_[15][1][96],
B_[15][2][96],
B_[0][0][97],
B_[0][1][97],
B_[0][2][97],
B_[1][0][97],
B_[1][1][97],
B_[1][2][97],
B_[2][0][97],
B_[2][1][97],
B_[2][2][97],
B_[3][0][97],
B_[3][1][97],
B_[3][2][97],
B_[4][0][97],
B_[4][1][97],
B_[4][2][97],
B_[5][0][97],
B_[5][1][97],
B_[5][2][97],
B_[6][0][97],
B_[6][1][97],
B_[6][2][97],
B_[7][0][97],
B_[7][1][97],
B_[7][2][97],
B_[8][0][97],
B_[8][1][97],
B_[8][2][97],
B_[9][0][97],
B_[9][1][97],
B_[9][2][97],
B_[10][0][97],
B_[10][1][97],
B_[10][2][97],
B_[11][0][97],
B_[11][1][97],
B_[11][2][97],
B_[12][0][97],
B_[12][1][97],
B_[12][2][97],
B_[13][0][97],
B_[13][1][97],
B_[13][2][97],
B_[14][0][97],
B_[14][1][97],
B_[14][2][97],
B_[15][0][97],
B_[15][1][97],
B_[15][2][97],
B_[0][0][98],
B_[0][1][98],
B_[0][2][98],
B_[1][0][98],
B_[1][1][98],
B_[1][2][98],
B_[2][0][98],
B_[2][1][98],
B_[2][2][98],
B_[3][0][98],
B_[3][1][98],
B_[3][2][98],
B_[4][0][98],
B_[4][1][98],
B_[4][2][98],
B_[5][0][98],
B_[5][1][98],
B_[5][2][98],
B_[6][0][98],
B_[6][1][98],
B_[6][2][98],
B_[7][0][98],
B_[7][1][98],
B_[7][2][98],
B_[8][0][98],
B_[8][1][98],
B_[8][2][98],
B_[9][0][98],
B_[9][1][98],
B_[9][2][98],
B_[10][0][98],
B_[10][1][98],
B_[10][2][98],
B_[11][0][98],
B_[11][1][98],
B_[11][2][98],
B_[12][0][98],
B_[12][1][98],
B_[12][2][98],
B_[13][0][98],
B_[13][1][98],
B_[13][2][98],
B_[14][0][98],
B_[14][1][98],
B_[14][2][98],
B_[15][0][98],
B_[15][1][98],
B_[15][2][98],
B_[0][0][99],
B_[0][1][99],
B_[0][2][99],
B_[1][0][99],
B_[1][1][99],
B_[1][2][99],
B_[2][0][99],
B_[2][1][99],
B_[2][2][99],
B_[3][0][99],
B_[3][1][99],
B_[3][2][99],
B_[4][0][99],
B_[4][1][99],
B_[4][2][99],
B_[5][0][99],
B_[5][1][99],
B_[5][2][99],
B_[6][0][99],
B_[6][1][99],
B_[6][2][99],
B_[7][0][99],
B_[7][1][99],
B_[7][2][99],
B_[8][0][99],
B_[8][1][99],
B_[8][2][99],
B_[9][0][99],
B_[9][1][99],
B_[9][2][99],
B_[10][0][99],
B_[10][1][99],
B_[10][2][99],
B_[11][0][99],
B_[11][1][99],
B_[11][2][99],
B_[12][0][99],
B_[12][1][99],
B_[12][2][99],
B_[13][0][99],
B_[13][1][99],
B_[13][2][99],
B_[14][0][99],
B_[14][1][99],
B_[14][2][99],
B_[15][0][99],
B_[15][1][99],
B_[15][2][99],
B_[0][0][100],
B_[0][1][100],
B_[0][2][100],
B_[1][0][100],
B_[1][1][100],
B_[1][2][100],
B_[2][0][100],
B_[2][1][100],
B_[2][2][100],
B_[3][0][100],
B_[3][1][100],
B_[3][2][100],
B_[4][0][100],
B_[4][1][100],
B_[4][2][100],
B_[5][0][100],
B_[5][1][100],
B_[5][2][100],
B_[6][0][100],
B_[6][1][100],
B_[6][2][100],
B_[7][0][100],
B_[7][1][100],
B_[7][2][100],
B_[8][0][100],
B_[8][1][100],
B_[8][2][100],
B_[9][0][100],
B_[9][1][100],
B_[9][2][100],
B_[10][0][100],
B_[10][1][100],
B_[10][2][100],
B_[11][0][100],
B_[11][1][100],
B_[11][2][100],
B_[12][0][100],
B_[12][1][100],
B_[12][2][100],
B_[13][0][100],
B_[13][1][100],
B_[13][2][100],
B_[14][0][100],
B_[14][1][100],
B_[14][2][100],
B_[15][0][100],
B_[15][1][100],
B_[15][2][100],
B_[0][0][101],
B_[0][1][101],
B_[0][2][101],
B_[1][0][101],
B_[1][1][101],
B_[1][2][101],
B_[2][0][101],
B_[2][1][101],
B_[2][2][101],
B_[3][0][101],
B_[3][1][101],
B_[3][2][101],
B_[4][0][101],
B_[4][1][101],
B_[4][2][101],
B_[5][0][101],
B_[5][1][101],
B_[5][2][101],
B_[6][0][101],
B_[6][1][101],
B_[6][2][101],
B_[7][0][101],
B_[7][1][101],
B_[7][2][101],
B_[8][0][101],
B_[8][1][101],
B_[8][2][101],
B_[9][0][101],
B_[9][1][101],
B_[9][2][101],
B_[10][0][101],
B_[10][1][101],
B_[10][2][101],
B_[11][0][101],
B_[11][1][101],
B_[11][2][101],
B_[12][0][101],
B_[12][1][101],
B_[12][2][101],
B_[13][0][101],
B_[13][1][101],
B_[13][2][101],
B_[14][0][101],
B_[14][1][101],
B_[14][2][101],
B_[15][0][101],
B_[15][1][101],
B_[15][2][101],
B_[0][0][102],
B_[0][1][102],
B_[0][2][102],
B_[1][0][102],
B_[1][1][102],
B_[1][2][102],
B_[2][0][102],
B_[2][1][102],
B_[2][2][102],
B_[3][0][102],
B_[3][1][102],
B_[3][2][102],
B_[4][0][102],
B_[4][1][102],
B_[4][2][102],
B_[5][0][102],
B_[5][1][102],
B_[5][2][102],
B_[6][0][102],
B_[6][1][102],
B_[6][2][102],
B_[7][0][102],
B_[7][1][102],
B_[7][2][102],
B_[8][0][102],
B_[8][1][102],
B_[8][2][102],
B_[9][0][102],
B_[9][1][102],
B_[9][2][102],
B_[10][0][102],
B_[10][1][102],
B_[10][2][102],
B_[11][0][102],
B_[11][1][102],
B_[11][2][102],
B_[12][0][102],
B_[12][1][102],
B_[12][2][102],
B_[13][0][102],
B_[13][1][102],
B_[13][2][102],
B_[14][0][102],
B_[14][1][102],
B_[14][2][102],
B_[15][0][102],
B_[15][1][102],
B_[15][2][102],
B_[0][0][103],
B_[0][1][103],
B_[0][2][103],
B_[1][0][103],
B_[1][1][103],
B_[1][2][103],
B_[2][0][103],
B_[2][1][103],
B_[2][2][103],
B_[3][0][103],
B_[3][1][103],
B_[3][2][103],
B_[4][0][103],
B_[4][1][103],
B_[4][2][103],
B_[5][0][103],
B_[5][1][103],
B_[5][2][103],
B_[6][0][103],
B_[6][1][103],
B_[6][2][103],
B_[7][0][103],
B_[7][1][103],
B_[7][2][103],
B_[8][0][103],
B_[8][1][103],
B_[8][2][103],
B_[9][0][103],
B_[9][1][103],
B_[9][2][103],
B_[10][0][103],
B_[10][1][103],
B_[10][2][103],
B_[11][0][103],
B_[11][1][103],
B_[11][2][103],
B_[12][0][103],
B_[12][1][103],
B_[12][2][103],
B_[13][0][103],
B_[13][1][103],
B_[13][2][103],
B_[14][0][103],
B_[14][1][103],
B_[14][2][103],
B_[15][0][103],
B_[15][1][103],
B_[15][2][103],
B_[0][0][104],
B_[0][1][104],
B_[0][2][104],
B_[1][0][104],
B_[1][1][104],
B_[1][2][104],
B_[2][0][104],
B_[2][1][104],
B_[2][2][104],
B_[3][0][104],
B_[3][1][104],
B_[3][2][104],
B_[4][0][104],
B_[4][1][104],
B_[4][2][104],
B_[5][0][104],
B_[5][1][104],
B_[5][2][104],
B_[6][0][104],
B_[6][1][104],
B_[6][2][104],
B_[7][0][104],
B_[7][1][104],
B_[7][2][104],
B_[8][0][104],
B_[8][1][104],
B_[8][2][104],
B_[9][0][104],
B_[9][1][104],
B_[9][2][104],
B_[10][0][104],
B_[10][1][104],
B_[10][2][104],
B_[11][0][104],
B_[11][1][104],
B_[11][2][104],
B_[12][0][104],
B_[12][1][104],
B_[12][2][104],
B_[13][0][104],
B_[13][1][104],
B_[13][2][104],
B_[14][0][104],
B_[14][1][104],
B_[14][2][104],
B_[15][0][104],
B_[15][1][104],
B_[15][2][104],
B_[0][0][105],
B_[0][1][105],
B_[0][2][105],
B_[1][0][105],
B_[1][1][105],
B_[1][2][105],
B_[2][0][105],
B_[2][1][105],
B_[2][2][105],
B_[3][0][105],
B_[3][1][105],
B_[3][2][105],
B_[4][0][105],
B_[4][1][105],
B_[4][2][105],
B_[5][0][105],
B_[5][1][105],
B_[5][2][105],
B_[6][0][105],
B_[6][1][105],
B_[6][2][105],
B_[7][0][105],
B_[7][1][105],
B_[7][2][105],
B_[8][0][105],
B_[8][1][105],
B_[8][2][105],
B_[9][0][105],
B_[9][1][105],
B_[9][2][105],
B_[10][0][105],
B_[10][1][105],
B_[10][2][105],
B_[11][0][105],
B_[11][1][105],
B_[11][2][105],
B_[12][0][105],
B_[12][1][105],
B_[12][2][105],
B_[13][0][105],
B_[13][1][105],
B_[13][2][105],
B_[14][0][105],
B_[14][1][105],
B_[14][2][105],
B_[15][0][105],
B_[15][1][105],
B_[15][2][105],
B_[0][0][106],
B_[0][1][106],
B_[0][2][106],
B_[1][0][106],
B_[1][1][106],
B_[1][2][106],
B_[2][0][106],
B_[2][1][106],
B_[2][2][106],
B_[3][0][106],
B_[3][1][106],
B_[3][2][106],
B_[4][0][106],
B_[4][1][106],
B_[4][2][106],
B_[5][0][106],
B_[5][1][106],
B_[5][2][106],
B_[6][0][106],
B_[6][1][106],
B_[6][2][106],
B_[7][0][106],
B_[7][1][106],
B_[7][2][106],
B_[8][0][106],
B_[8][1][106],
B_[8][2][106],
B_[9][0][106],
B_[9][1][106],
B_[9][2][106],
B_[10][0][106],
B_[10][1][106],
B_[10][2][106],
B_[11][0][106],
B_[11][1][106],
B_[11][2][106],
B_[12][0][106],
B_[12][1][106],
B_[12][2][106],
B_[13][0][106],
B_[13][1][106],
B_[13][2][106],
B_[14][0][106],
B_[14][1][106],
B_[14][2][106],
B_[15][0][106],
B_[15][1][106],
B_[15][2][106],
B_[0][0][107],
B_[0][1][107],
B_[0][2][107],
B_[1][0][107],
B_[1][1][107],
B_[1][2][107],
B_[2][0][107],
B_[2][1][107],
B_[2][2][107],
B_[3][0][107],
B_[3][1][107],
B_[3][2][107],
B_[4][0][107],
B_[4][1][107],
B_[4][2][107],
B_[5][0][107],
B_[5][1][107],
B_[5][2][107],
B_[6][0][107],
B_[6][1][107],
B_[6][2][107],
B_[7][0][107],
B_[7][1][107],
B_[7][2][107],
B_[8][0][107],
B_[8][1][107],
B_[8][2][107],
B_[9][0][107],
B_[9][1][107],
B_[9][2][107],
B_[10][0][107],
B_[10][1][107],
B_[10][2][107],
B_[11][0][107],
B_[11][1][107],
B_[11][2][107],
B_[12][0][107],
B_[12][1][107],
B_[12][2][107],
B_[13][0][107],
B_[13][1][107],
B_[13][2][107],
B_[14][0][107],
B_[14][1][107],
B_[14][2][107],
B_[15][0][107],
B_[15][1][107],
B_[15][2][107],
B_[0][0][108],
B_[0][1][108],
B_[0][2][108],
B_[1][0][108],
B_[1][1][108],
B_[1][2][108],
B_[2][0][108],
B_[2][1][108],
B_[2][2][108],
B_[3][0][108],
B_[3][1][108],
B_[3][2][108],
B_[4][0][108],
B_[4][1][108],
B_[4][2][108],
B_[5][0][108],
B_[5][1][108],
B_[5][2][108],
B_[6][0][108],
B_[6][1][108],
B_[6][2][108],
B_[7][0][108],
B_[7][1][108],
B_[7][2][108],
B_[8][0][108],
B_[8][1][108],
B_[8][2][108],
B_[9][0][108],
B_[9][1][108],
B_[9][2][108],
B_[10][0][108],
B_[10][1][108],
B_[10][2][108],
B_[11][0][108],
B_[11][1][108],
B_[11][2][108],
B_[12][0][108],
B_[12][1][108],
B_[12][2][108],
B_[13][0][108],
B_[13][1][108],
B_[13][2][108],
B_[14][0][108],
B_[14][1][108],
B_[14][2][108],
B_[15][0][108],
B_[15][1][108],
B_[15][2][108],
B_[0][0][109],
B_[0][1][109],
B_[0][2][109],
B_[1][0][109],
B_[1][1][109],
B_[1][2][109],
B_[2][0][109],
B_[2][1][109],
B_[2][2][109],
B_[3][0][109],
B_[3][1][109],
B_[3][2][109],
B_[4][0][109],
B_[4][1][109],
B_[4][2][109],
B_[5][0][109],
B_[5][1][109],
B_[5][2][109],
B_[6][0][109],
B_[6][1][109],
B_[6][2][109],
B_[7][0][109],
B_[7][1][109],
B_[7][2][109],
B_[8][0][109],
B_[8][1][109],
B_[8][2][109],
B_[9][0][109],
B_[9][1][109],
B_[9][2][109],
B_[10][0][109],
B_[10][1][109],
B_[10][2][109],
B_[11][0][109],
B_[11][1][109],
B_[11][2][109],
B_[12][0][109],
B_[12][1][109],
B_[12][2][109],
B_[13][0][109],
B_[13][1][109],
B_[13][2][109],
B_[14][0][109],
B_[14][1][109],
B_[14][2][109],
B_[15][0][109],
B_[15][1][109],
B_[15][2][109],
B_[0][0][110],
B_[0][1][110],
B_[0][2][110],
B_[1][0][110],
B_[1][1][110],
B_[1][2][110],
B_[2][0][110],
B_[2][1][110],
B_[2][2][110],
B_[3][0][110],
B_[3][1][110],
B_[3][2][110],
B_[4][0][110],
B_[4][1][110],
B_[4][2][110],
B_[5][0][110],
B_[5][1][110],
B_[5][2][110],
B_[6][0][110],
B_[6][1][110],
B_[6][2][110],
B_[7][0][110],
B_[7][1][110],
B_[7][2][110],
B_[8][0][110],
B_[8][1][110],
B_[8][2][110],
B_[9][0][110],
B_[9][1][110],
B_[9][2][110],
B_[10][0][110],
B_[10][1][110],
B_[10][2][110],
B_[11][0][110],
B_[11][1][110],
B_[11][2][110],
B_[12][0][110],
B_[12][1][110],
B_[12][2][110],
B_[13][0][110],
B_[13][1][110],
B_[13][2][110],
B_[14][0][110],
B_[14][1][110],
B_[14][2][110],
B_[15][0][110],
B_[15][1][110],
B_[15][2][110],
B_[0][0][111],
B_[0][1][111],
B_[0][2][111],
B_[1][0][111],
B_[1][1][111],
B_[1][2][111],
B_[2][0][111],
B_[2][1][111],
B_[2][2][111],
B_[3][0][111],
B_[3][1][111],
B_[3][2][111],
B_[4][0][111],
B_[4][1][111],
B_[4][2][111],
B_[5][0][111],
B_[5][1][111],
B_[5][2][111],
B_[6][0][111],
B_[6][1][111],
B_[6][2][111],
B_[7][0][111],
B_[7][1][111],
B_[7][2][111],
B_[8][0][111],
B_[8][1][111],
B_[8][2][111],
B_[9][0][111],
B_[9][1][111],
B_[9][2][111],
B_[10][0][111],
B_[10][1][111],
B_[10][2][111],
B_[11][0][111],
B_[11][1][111],
B_[11][2][111],
B_[12][0][111],
B_[12][1][111],
B_[12][2][111],
B_[13][0][111],
B_[13][1][111],
B_[13][2][111],
B_[14][0][111],
B_[14][1][111],
B_[14][2][111],
B_[15][0][111],
B_[15][1][111],
B_[15][2][111],
B_[0][0][112],
B_[0][1][112],
B_[0][2][112],
B_[1][0][112],
B_[1][1][112],
B_[1][2][112],
B_[2][0][112],
B_[2][1][112],
B_[2][2][112],
B_[3][0][112],
B_[3][1][112],
B_[3][2][112],
B_[4][0][112],
B_[4][1][112],
B_[4][2][112],
B_[5][0][112],
B_[5][1][112],
B_[5][2][112],
B_[6][0][112],
B_[6][1][112],
B_[6][2][112],
B_[7][0][112],
B_[7][1][112],
B_[7][2][112],
B_[8][0][112],
B_[8][1][112],
B_[8][2][112],
B_[9][0][112],
B_[9][1][112],
B_[9][2][112],
B_[10][0][112],
B_[10][1][112],
B_[10][2][112],
B_[11][0][112],
B_[11][1][112],
B_[11][2][112],
B_[12][0][112],
B_[12][1][112],
B_[12][2][112],
B_[13][0][112],
B_[13][1][112],
B_[13][2][112],
B_[14][0][112],
B_[14][1][112],
B_[14][2][112],
B_[15][0][112],
B_[15][1][112],
B_[15][2][112],
B_[0][0][113],
B_[0][1][113],
B_[0][2][113],
B_[1][0][113],
B_[1][1][113],
B_[1][2][113],
B_[2][0][113],
B_[2][1][113],
B_[2][2][113],
B_[3][0][113],
B_[3][1][113],
B_[3][2][113],
B_[4][0][113],
B_[4][1][113],
B_[4][2][113],
B_[5][0][113],
B_[5][1][113],
B_[5][2][113],
B_[6][0][113],
B_[6][1][113],
B_[6][2][113],
B_[7][0][113],
B_[7][1][113],
B_[7][2][113],
B_[8][0][113],
B_[8][1][113],
B_[8][2][113],
B_[9][0][113],
B_[9][1][113],
B_[9][2][113],
B_[10][0][113],
B_[10][1][113],
B_[10][2][113],
B_[11][0][113],
B_[11][1][113],
B_[11][2][113],
B_[12][0][113],
B_[12][1][113],
B_[12][2][113],
B_[13][0][113],
B_[13][1][113],
B_[13][2][113],
B_[14][0][113],
B_[14][1][113],
B_[14][2][113],
B_[15][0][113],
B_[15][1][113],
B_[15][2][113],
B_[0][0][114],
B_[0][1][114],
B_[0][2][114],
B_[1][0][114],
B_[1][1][114],
B_[1][2][114],
B_[2][0][114],
B_[2][1][114],
B_[2][2][114],
B_[3][0][114],
B_[3][1][114],
B_[3][2][114],
B_[4][0][114],
B_[4][1][114],
B_[4][2][114],
B_[5][0][114],
B_[5][1][114],
B_[5][2][114],
B_[6][0][114],
B_[6][1][114],
B_[6][2][114],
B_[7][0][114],
B_[7][1][114],
B_[7][2][114],
B_[8][0][114],
B_[8][1][114],
B_[8][2][114],
B_[9][0][114],
B_[9][1][114],
B_[9][2][114],
B_[10][0][114],
B_[10][1][114],
B_[10][2][114],
B_[11][0][114],
B_[11][1][114],
B_[11][2][114],
B_[12][0][114],
B_[12][1][114],
B_[12][2][114],
B_[13][0][114],
B_[13][1][114],
B_[13][2][114],
B_[14][0][114],
B_[14][1][114],
B_[14][2][114],
B_[15][0][114],
B_[15][1][114],
B_[15][2][114],
B_[0][0][115],
B_[0][1][115],
B_[0][2][115],
B_[1][0][115],
B_[1][1][115],
B_[1][2][115],
B_[2][0][115],
B_[2][1][115],
B_[2][2][115],
B_[3][0][115],
B_[3][1][115],
B_[3][2][115],
B_[4][0][115],
B_[4][1][115],
B_[4][2][115],
B_[5][0][115],
B_[5][1][115],
B_[5][2][115],
B_[6][0][115],
B_[6][1][115],
B_[6][2][115],
B_[7][0][115],
B_[7][1][115],
B_[7][2][115],
B_[8][0][115],
B_[8][1][115],
B_[8][2][115],
B_[9][0][115],
B_[9][1][115],
B_[9][2][115],
B_[10][0][115],
B_[10][1][115],
B_[10][2][115],
B_[11][0][115],
B_[11][1][115],
B_[11][2][115],
B_[12][0][115],
B_[12][1][115],
B_[12][2][115],
B_[13][0][115],
B_[13][1][115],
B_[13][2][115],
B_[14][0][115],
B_[14][1][115],
B_[14][2][115],
B_[15][0][115],
B_[15][1][115],
B_[15][2][115],
B_[0][0][116],
B_[0][1][116],
B_[0][2][116],
B_[1][0][116],
B_[1][1][116],
B_[1][2][116],
B_[2][0][116],
B_[2][1][116],
B_[2][2][116],
B_[3][0][116],
B_[3][1][116],
B_[3][2][116],
B_[4][0][116],
B_[4][1][116],
B_[4][2][116],
B_[5][0][116],
B_[5][1][116],
B_[5][2][116],
B_[6][0][116],
B_[6][1][116],
B_[6][2][116],
B_[7][0][116],
B_[7][1][116],
B_[7][2][116],
B_[8][0][116],
B_[8][1][116],
B_[8][2][116],
B_[9][0][116],
B_[9][1][116],
B_[9][2][116],
B_[10][0][116],
B_[10][1][116],
B_[10][2][116],
B_[11][0][116],
B_[11][1][116],
B_[11][2][116],
B_[12][0][116],
B_[12][1][116],
B_[12][2][116],
B_[13][0][116],
B_[13][1][116],
B_[13][2][116],
B_[14][0][116],
B_[14][1][116],
B_[14][2][116],
B_[15][0][116],
B_[15][1][116],
B_[15][2][116],
B_[0][0][117],
B_[0][1][117],
B_[0][2][117],
B_[1][0][117],
B_[1][1][117],
B_[1][2][117],
B_[2][0][117],
B_[2][1][117],
B_[2][2][117],
B_[3][0][117],
B_[3][1][117],
B_[3][2][117],
B_[4][0][117],
B_[4][1][117],
B_[4][2][117],
B_[5][0][117],
B_[5][1][117],
B_[5][2][117],
B_[6][0][117],
B_[6][1][117],
B_[6][2][117],
B_[7][0][117],
B_[7][1][117],
B_[7][2][117],
B_[8][0][117],
B_[8][1][117],
B_[8][2][117],
B_[9][0][117],
B_[9][1][117],
B_[9][2][117],
B_[10][0][117],
B_[10][1][117],
B_[10][2][117],
B_[11][0][117],
B_[11][1][117],
B_[11][2][117],
B_[12][0][117],
B_[12][1][117],
B_[12][2][117],
B_[13][0][117],
B_[13][1][117],
B_[13][2][117],
B_[14][0][117],
B_[14][1][117],
B_[14][2][117],
B_[15][0][117],
B_[15][1][117],
B_[15][2][117],
B_[0][0][118],
B_[0][1][118],
B_[0][2][118],
B_[1][0][118],
B_[1][1][118],
B_[1][2][118],
B_[2][0][118],
B_[2][1][118],
B_[2][2][118],
B_[3][0][118],
B_[3][1][118],
B_[3][2][118],
B_[4][0][118],
B_[4][1][118],
B_[4][2][118],
B_[5][0][118],
B_[5][1][118],
B_[5][2][118],
B_[6][0][118],
B_[6][1][118],
B_[6][2][118],
B_[7][0][118],
B_[7][1][118],
B_[7][2][118],
B_[8][0][118],
B_[8][1][118],
B_[8][2][118],
B_[9][0][118],
B_[9][1][118],
B_[9][2][118],
B_[10][0][118],
B_[10][1][118],
B_[10][2][118],
B_[11][0][118],
B_[11][1][118],
B_[11][2][118],
B_[12][0][118],
B_[12][1][118],
B_[12][2][118],
B_[13][0][118],
B_[13][1][118],
B_[13][2][118],
B_[14][0][118],
B_[14][1][118],
B_[14][2][118],
B_[15][0][118],
B_[15][1][118],
B_[15][2][118],
B_[0][0][119],
B_[0][1][119],
B_[0][2][119],
B_[1][0][119],
B_[1][1][119],
B_[1][2][119],
B_[2][0][119],
B_[2][1][119],
B_[2][2][119],
B_[3][0][119],
B_[3][1][119],
B_[3][2][119],
B_[4][0][119],
B_[4][1][119],
B_[4][2][119],
B_[5][0][119],
B_[5][1][119],
B_[5][2][119],
B_[6][0][119],
B_[6][1][119],
B_[6][2][119],
B_[7][0][119],
B_[7][1][119],
B_[7][2][119],
B_[8][0][119],
B_[8][1][119],
B_[8][2][119],
B_[9][0][119],
B_[9][1][119],
B_[9][2][119],
B_[10][0][119],
B_[10][1][119],
B_[10][2][119],
B_[11][0][119],
B_[11][1][119],
B_[11][2][119],
B_[12][0][119],
B_[12][1][119],
B_[12][2][119],
B_[13][0][119],
B_[13][1][119],
B_[13][2][119],
B_[14][0][119],
B_[14][1][119],
B_[14][2][119],
B_[15][0][119],
B_[15][1][119],
B_[15][2][119],
B_[0][0][120],
B_[0][1][120],
B_[0][2][120],
B_[1][0][120],
B_[1][1][120],
B_[1][2][120],
B_[2][0][120],
B_[2][1][120],
B_[2][2][120],
B_[3][0][120],
B_[3][1][120],
B_[3][2][120],
B_[4][0][120],
B_[4][1][120],
B_[4][2][120],
B_[5][0][120],
B_[5][1][120],
B_[5][2][120],
B_[6][0][120],
B_[6][1][120],
B_[6][2][120],
B_[7][0][120],
B_[7][1][120],
B_[7][2][120],
B_[8][0][120],
B_[8][1][120],
B_[8][2][120],
B_[9][0][120],
B_[9][1][120],
B_[9][2][120],
B_[10][0][120],
B_[10][1][120],
B_[10][2][120],
B_[11][0][120],
B_[11][1][120],
B_[11][2][120],
B_[12][0][120],
B_[12][1][120],
B_[12][2][120],
B_[13][0][120],
B_[13][1][120],
B_[13][2][120],
B_[14][0][120],
B_[14][1][120],
B_[14][2][120],
B_[15][0][120],
B_[15][1][120],
B_[15][2][120],
B_[0][0][121],
B_[0][1][121],
B_[0][2][121],
B_[1][0][121],
B_[1][1][121],
B_[1][2][121],
B_[2][0][121],
B_[2][1][121],
B_[2][2][121],
B_[3][0][121],
B_[3][1][121],
B_[3][2][121],
B_[4][0][121],
B_[4][1][121],
B_[4][2][121],
B_[5][0][121],
B_[5][1][121],
B_[5][2][121],
B_[6][0][121],
B_[6][1][121],
B_[6][2][121],
B_[7][0][121],
B_[7][1][121],
B_[7][2][121],
B_[8][0][121],
B_[8][1][121],
B_[8][2][121],
B_[9][0][121],
B_[9][1][121],
B_[9][2][121],
B_[10][0][121],
B_[10][1][121],
B_[10][2][121],
B_[11][0][121],
B_[11][1][121],
B_[11][2][121],
B_[12][0][121],
B_[12][1][121],
B_[12][2][121],
B_[13][0][121],
B_[13][1][121],
B_[13][2][121],
B_[14][0][121],
B_[14][1][121],
B_[14][2][121],
B_[15][0][121],
B_[15][1][121],
B_[15][2][121],
B_[0][0][122],
B_[0][1][122],
B_[0][2][122],
B_[1][0][122],
B_[1][1][122],
B_[1][2][122],
B_[2][0][122],
B_[2][1][122],
B_[2][2][122],
B_[3][0][122],
B_[3][1][122],
B_[3][2][122],
B_[4][0][122],
B_[4][1][122],
B_[4][2][122],
B_[5][0][122],
B_[5][1][122],
B_[5][2][122],
B_[6][0][122],
B_[6][1][122],
B_[6][2][122],
B_[7][0][122],
B_[7][1][122],
B_[7][2][122],
B_[8][0][122],
B_[8][1][122],
B_[8][2][122],
B_[9][0][122],
B_[9][1][122],
B_[9][2][122],
B_[10][0][122],
B_[10][1][122],
B_[10][2][122],
B_[11][0][122],
B_[11][1][122],
B_[11][2][122],
B_[12][0][122],
B_[12][1][122],
B_[12][2][122],
B_[13][0][122],
B_[13][1][122],
B_[13][2][122],
B_[14][0][122],
B_[14][1][122],
B_[14][2][122],
B_[15][0][122],
B_[15][1][122],
B_[15][2][122],
B_[0][0][123],
B_[0][1][123],
B_[0][2][123],
B_[1][0][123],
B_[1][1][123],
B_[1][2][123],
B_[2][0][123],
B_[2][1][123],
B_[2][2][123],
B_[3][0][123],
B_[3][1][123],
B_[3][2][123],
B_[4][0][123],
B_[4][1][123],
B_[4][2][123],
B_[5][0][123],
B_[5][1][123],
B_[5][2][123],
B_[6][0][123],
B_[6][1][123],
B_[6][2][123],
B_[7][0][123],
B_[7][1][123],
B_[7][2][123],
B_[8][0][123],
B_[8][1][123],
B_[8][2][123],
B_[9][0][123],
B_[9][1][123],
B_[9][2][123],
B_[10][0][123],
B_[10][1][123],
B_[10][2][123],
B_[11][0][123],
B_[11][1][123],
B_[11][2][123],
B_[12][0][123],
B_[12][1][123],
B_[12][2][123],
B_[13][0][123],
B_[13][1][123],
B_[13][2][123],
B_[14][0][123],
B_[14][1][123],
B_[14][2][123],
B_[15][0][123],
B_[15][1][123],
B_[15][2][123],
B_[0][0][124],
B_[0][1][124],
B_[0][2][124],
B_[1][0][124],
B_[1][1][124],
B_[1][2][124],
B_[2][0][124],
B_[2][1][124],
B_[2][2][124],
B_[3][0][124],
B_[3][1][124],
B_[3][2][124],
B_[4][0][124],
B_[4][1][124],
B_[4][2][124],
B_[5][0][124],
B_[5][1][124],
B_[5][2][124],
B_[6][0][124],
B_[6][1][124],
B_[6][2][124],
B_[7][0][124],
B_[7][1][124],
B_[7][2][124],
B_[8][0][124],
B_[8][1][124],
B_[8][2][124],
B_[9][0][124],
B_[9][1][124],
B_[9][2][124],
B_[10][0][124],
B_[10][1][124],
B_[10][2][124],
B_[11][0][124],
B_[11][1][124],
B_[11][2][124],
B_[12][0][124],
B_[12][1][124],
B_[12][2][124],
B_[13][0][124],
B_[13][1][124],
B_[13][2][124],
B_[14][0][124],
B_[14][1][124],
B_[14][2][124],
B_[15][0][124],
B_[15][1][124],
B_[15][2][124],
B_[0][0][125],
B_[0][1][125],
B_[0][2][125],
B_[1][0][125],
B_[1][1][125],
B_[1][2][125],
B_[2][0][125],
B_[2][1][125],
B_[2][2][125],
B_[3][0][125],
B_[3][1][125],
B_[3][2][125],
B_[4][0][125],
B_[4][1][125],
B_[4][2][125],
B_[5][0][125],
B_[5][1][125],
B_[5][2][125],
B_[6][0][125],
B_[6][1][125],
B_[6][2][125],
B_[7][0][125],
B_[7][1][125],
B_[7][2][125],
B_[8][0][125],
B_[8][1][125],
B_[8][2][125],
B_[9][0][125],
B_[9][1][125],
B_[9][2][125],
B_[10][0][125],
B_[10][1][125],
B_[10][2][125],
B_[11][0][125],
B_[11][1][125],
B_[11][2][125],
B_[12][0][125],
B_[12][1][125],
B_[12][2][125],
B_[13][0][125],
B_[13][1][125],
B_[13][2][125],
B_[14][0][125],
B_[14][1][125],
B_[14][2][125],
B_[15][0][125],
B_[15][1][125],
B_[15][2][125],
B_[0][0][126],
B_[0][1][126],
B_[0][2][126],
B_[1][0][126],
B_[1][1][126],
B_[1][2][126],
B_[2][0][126],
B_[2][1][126],
B_[2][2][126],
B_[3][0][126],
B_[3][1][126],
B_[3][2][126],
B_[4][0][126],
B_[4][1][126],
B_[4][2][126],
B_[5][0][126],
B_[5][1][126],
B_[5][2][126],
B_[6][0][126],
B_[6][1][126],
B_[6][2][126],
B_[7][0][126],
B_[7][1][126],
B_[7][2][126],
B_[8][0][126],
B_[8][1][126],
B_[8][2][126],
B_[9][0][126],
B_[9][1][126],
B_[9][2][126],
B_[10][0][126],
B_[10][1][126],
B_[10][2][126],
B_[11][0][126],
B_[11][1][126],
B_[11][2][126],
B_[12][0][126],
B_[12][1][126],
B_[12][2][126],
B_[13][0][126],
B_[13][1][126],
B_[13][2][126],
B_[14][0][126],
B_[14][1][126],
B_[14][2][126],
B_[15][0][126],
B_[15][1][126],
B_[15][2][126],
B_[0][0][127],
B_[0][1][127],
B_[0][2][127],
B_[1][0][127],
B_[1][1][127],
B_[1][2][127],
B_[2][0][127],
B_[2][1][127],
B_[2][2][127],
B_[3][0][127],
B_[3][1][127],
B_[3][2][127],
B_[4][0][127],
B_[4][1][127],
B_[4][2][127],
B_[5][0][127],
B_[5][1][127],
B_[5][2][127],
B_[6][0][127],
B_[6][1][127],
B_[6][2][127],
B_[7][0][127],
B_[7][1][127],
B_[7][2][127],
B_[8][0][127],
B_[8][1][127],
B_[8][2][127],
B_[9][0][127],
B_[9][1][127],
B_[9][2][127],
B_[10][0][127],
B_[10][1][127],
B_[10][2][127],
B_[11][0][127],
B_[11][1][127],
B_[11][2][127],
B_[12][0][127],
B_[12][1][127],
B_[12][2][127],
B_[13][0][127],
B_[13][1][127],
B_[13][2][127],
B_[14][0][127],
B_[14][1][127],
B_[14][2][127],
B_[15][0][127],
B_[15][1][127],
B_[15][2][127],
B_[0][0][128],
B_[0][1][128],
B_[0][2][128],
B_[1][0][128],
B_[1][1][128],
B_[1][2][128],
B_[2][0][128],
B_[2][1][128],
B_[2][2][128],
B_[3][0][128],
B_[3][1][128],
B_[3][2][128],
B_[4][0][128],
B_[4][1][128],
B_[4][2][128],
B_[5][0][128],
B_[5][1][128],
B_[5][2][128],
B_[6][0][128],
B_[6][1][128],
B_[6][2][128],
B_[7][0][128],
B_[7][1][128],
B_[7][2][128],
B_[8][0][128],
B_[8][1][128],
B_[8][2][128],
B_[9][0][128],
B_[9][1][128],
B_[9][2][128],
B_[10][0][128],
B_[10][1][128],
B_[10][2][128],
B_[11][0][128],
B_[11][1][128],
B_[11][2][128],
B_[12][0][128],
B_[12][1][128],
B_[12][2][128],
B_[13][0][128],
B_[13][1][128],
B_[13][2][128],
B_[14][0][128],
B_[14][1][128],
B_[14][2][128],
B_[15][0][128],
B_[15][1][128],
B_[15][2][128],
B_[0][0][129],
B_[0][1][129],
B_[0][2][129],
B_[1][0][129],
B_[1][1][129],
B_[1][2][129],
B_[2][0][129],
B_[2][1][129],
B_[2][2][129],
B_[3][0][129],
B_[3][1][129],
B_[3][2][129],
B_[4][0][129],
B_[4][1][129],
B_[4][2][129],
B_[5][0][129],
B_[5][1][129],
B_[5][2][129],
B_[6][0][129],
B_[6][1][129],
B_[6][2][129],
B_[7][0][129],
B_[7][1][129],
B_[7][2][129],
B_[8][0][129],
B_[8][1][129],
B_[8][2][129],
B_[9][0][129],
B_[9][1][129],
B_[9][2][129],
B_[10][0][129],
B_[10][1][129],
B_[10][2][129],
B_[11][0][129],
B_[11][1][129],
B_[11][2][129],
B_[12][0][129],
B_[12][1][129],
B_[12][2][129],
B_[13][0][129],
B_[13][1][129],
B_[13][2][129],
B_[14][0][129],
B_[14][1][129],
B_[14][2][129],
B_[15][0][129],
B_[15][1][129],
B_[15][2][129],
B_[0][0][130],
B_[0][1][130],
B_[0][2][130],
B_[1][0][130],
B_[1][1][130],
B_[1][2][130],
B_[2][0][130],
B_[2][1][130],
B_[2][2][130],
B_[3][0][130],
B_[3][1][130],
B_[3][2][130],
B_[4][0][130],
B_[4][1][130],
B_[4][2][130],
B_[5][0][130],
B_[5][1][130],
B_[5][2][130],
B_[6][0][130],
B_[6][1][130],
B_[6][2][130],
B_[7][0][130],
B_[7][1][130],
B_[7][2][130],
B_[8][0][130],
B_[8][1][130],
B_[8][2][130],
B_[9][0][130],
B_[9][1][130],
B_[9][2][130],
B_[10][0][130],
B_[10][1][130],
B_[10][2][130],
B_[11][0][130],
B_[11][1][130],
B_[11][2][130],
B_[12][0][130],
B_[12][1][130],
B_[12][2][130],
B_[13][0][130],
B_[13][1][130],
B_[13][2][130],
B_[14][0][130],
B_[14][1][130],
B_[14][2][130],
B_[15][0][130],
B_[15][1][130],
B_[15][2][130],
B_[0][0][131],
B_[0][1][131],
B_[0][2][131],
B_[1][0][131],
B_[1][1][131],
B_[1][2][131],
B_[2][0][131],
B_[2][1][131],
B_[2][2][131],
B_[3][0][131],
B_[3][1][131],
B_[3][2][131],
B_[4][0][131],
B_[4][1][131],
B_[4][2][131],
B_[5][0][131],
B_[5][1][131],
B_[5][2][131],
B_[6][0][131],
B_[6][1][131],
B_[6][2][131],
B_[7][0][131],
B_[7][1][131],
B_[7][2][131],
B_[8][0][131],
B_[8][1][131],
B_[8][2][131],
B_[9][0][131],
B_[9][1][131],
B_[9][2][131],
B_[10][0][131],
B_[10][1][131],
B_[10][2][131],
B_[11][0][131],
B_[11][1][131],
B_[11][2][131],
B_[12][0][131],
B_[12][1][131],
B_[12][2][131],
B_[13][0][131],
B_[13][1][131],
B_[13][2][131],
B_[14][0][131],
B_[14][1][131],
B_[14][2][131],
B_[15][0][131],
B_[15][1][131],
B_[15][2][131],
B_[0][0][132],
B_[0][1][132],
B_[0][2][132],
B_[1][0][132],
B_[1][1][132],
B_[1][2][132],
B_[2][0][132],
B_[2][1][132],
B_[2][2][132],
B_[3][0][132],
B_[3][1][132],
B_[3][2][132],
B_[4][0][132],
B_[4][1][132],
B_[4][2][132],
B_[5][0][132],
B_[5][1][132],
B_[5][2][132],
B_[6][0][132],
B_[6][1][132],
B_[6][2][132],
B_[7][0][132],
B_[7][1][132],
B_[7][2][132],
B_[8][0][132],
B_[8][1][132],
B_[8][2][132],
B_[9][0][132],
B_[9][1][132],
B_[9][2][132],
B_[10][0][132],
B_[10][1][132],
B_[10][2][132],
B_[11][0][132],
B_[11][1][132],
B_[11][2][132],
B_[12][0][132],
B_[12][1][132],
B_[12][2][132],
B_[13][0][132],
B_[13][1][132],
B_[13][2][132],
B_[14][0][132],
B_[14][1][132],
B_[14][2][132],
B_[15][0][132],
B_[15][1][132],
B_[15][2][132],
B_[0][0][133],
B_[0][1][133],
B_[0][2][133],
B_[1][0][133],
B_[1][1][133],
B_[1][2][133],
B_[2][0][133],
B_[2][1][133],
B_[2][2][133],
B_[3][0][133],
B_[3][1][133],
B_[3][2][133],
B_[4][0][133],
B_[4][1][133],
B_[4][2][133],
B_[5][0][133],
B_[5][1][133],
B_[5][2][133],
B_[6][0][133],
B_[6][1][133],
B_[6][2][133],
B_[7][0][133],
B_[7][1][133],
B_[7][2][133],
B_[8][0][133],
B_[8][1][133],
B_[8][2][133],
B_[9][0][133],
B_[9][1][133],
B_[9][2][133],
B_[10][0][133],
B_[10][1][133],
B_[10][2][133],
B_[11][0][133],
B_[11][1][133],
B_[11][2][133],
B_[12][0][133],
B_[12][1][133],
B_[12][2][133],
B_[13][0][133],
B_[13][1][133],
B_[13][2][133],
B_[14][0][133],
B_[14][1][133],
B_[14][2][133],
B_[15][0][133],
B_[15][1][133],
B_[15][2][133],
B_[0][0][134],
B_[0][1][134],
B_[0][2][134],
B_[1][0][134],
B_[1][1][134],
B_[1][2][134],
B_[2][0][134],
B_[2][1][134],
B_[2][2][134],
B_[3][0][134],
B_[3][1][134],
B_[3][2][134],
B_[4][0][134],
B_[4][1][134],
B_[4][2][134],
B_[5][0][134],
B_[5][1][134],
B_[5][2][134],
B_[6][0][134],
B_[6][1][134],
B_[6][2][134],
B_[7][0][134],
B_[7][1][134],
B_[7][2][134],
B_[8][0][134],
B_[8][1][134],
B_[8][2][134],
B_[9][0][134],
B_[9][1][134],
B_[9][2][134],
B_[10][0][134],
B_[10][1][134],
B_[10][2][134],
B_[11][0][134],
B_[11][1][134],
B_[11][2][134],
B_[12][0][134],
B_[12][1][134],
B_[12][2][134],
B_[13][0][134],
B_[13][1][134],
B_[13][2][134],
B_[14][0][134],
B_[14][1][134],
B_[14][2][134],
B_[15][0][134],
B_[15][1][134],
B_[15][2][134],
B_[0][0][135],
B_[0][1][135],
B_[0][2][135],
B_[1][0][135],
B_[1][1][135],
B_[1][2][135],
B_[2][0][135],
B_[2][1][135],
B_[2][2][135],
B_[3][0][135],
B_[3][1][135],
B_[3][2][135],
B_[4][0][135],
B_[4][1][135],
B_[4][2][135],
B_[5][0][135],
B_[5][1][135],
B_[5][2][135],
B_[6][0][135],
B_[6][1][135],
B_[6][2][135],
B_[7][0][135],
B_[7][1][135],
B_[7][2][135],
B_[8][0][135],
B_[8][1][135],
B_[8][2][135],
B_[9][0][135],
B_[9][1][135],
B_[9][2][135],
B_[10][0][135],
B_[10][1][135],
B_[10][2][135],
B_[11][0][135],
B_[11][1][135],
B_[11][2][135],
B_[12][0][135],
B_[12][1][135],
B_[12][2][135],
B_[13][0][135],
B_[13][1][135],
B_[13][2][135],
B_[14][0][135],
B_[14][1][135],
B_[14][2][135],
B_[15][0][135],
B_[15][1][135],
B_[15][2][135],
B_[0][0][136],
B_[0][1][136],
B_[0][2][136],
B_[1][0][136],
B_[1][1][136],
B_[1][2][136],
B_[2][0][136],
B_[2][1][136],
B_[2][2][136],
B_[3][0][136],
B_[3][1][136],
B_[3][2][136],
B_[4][0][136],
B_[4][1][136],
B_[4][2][136],
B_[5][0][136],
B_[5][1][136],
B_[5][2][136],
B_[6][0][136],
B_[6][1][136],
B_[6][2][136],
B_[7][0][136],
B_[7][1][136],
B_[7][2][136],
B_[8][0][136],
B_[8][1][136],
B_[8][2][136],
B_[9][0][136],
B_[9][1][136],
B_[9][2][136],
B_[10][0][136],
B_[10][1][136],
B_[10][2][136],
B_[11][0][136],
B_[11][1][136],
B_[11][2][136],
B_[12][0][136],
B_[12][1][136],
B_[12][2][136],
B_[13][0][136],
B_[13][1][136],
B_[13][2][136],
B_[14][0][136],
B_[14][1][136],
B_[14][2][136],
B_[15][0][136],
B_[15][1][136],
B_[15][2][136],
B_[0][0][137],
B_[0][1][137],
B_[0][2][137],
B_[1][0][137],
B_[1][1][137],
B_[1][2][137],
B_[2][0][137],
B_[2][1][137],
B_[2][2][137],
B_[3][0][137],
B_[3][1][137],
B_[3][2][137],
B_[4][0][137],
B_[4][1][137],
B_[4][2][137],
B_[5][0][137],
B_[5][1][137],
B_[5][2][137],
B_[6][0][137],
B_[6][1][137],
B_[6][2][137],
B_[7][0][137],
B_[7][1][137],
B_[7][2][137],
B_[8][0][137],
B_[8][1][137],
B_[8][2][137],
B_[9][0][137],
B_[9][1][137],
B_[9][2][137],
B_[10][0][137],
B_[10][1][137],
B_[10][2][137],
B_[11][0][137],
B_[11][1][137],
B_[11][2][137],
B_[12][0][137],
B_[12][1][137],
B_[12][2][137],
B_[13][0][137],
B_[13][1][137],
B_[13][2][137],
B_[14][0][137],
B_[14][1][137],
B_[14][2][137],
B_[15][0][137],
B_[15][1][137],
B_[15][2][137],
B_[0][0][138],
B_[0][1][138],
B_[0][2][138],
B_[1][0][138],
B_[1][1][138],
B_[1][2][138],
B_[2][0][138],
B_[2][1][138],
B_[2][2][138],
B_[3][0][138],
B_[3][1][138],
B_[3][2][138],
B_[4][0][138],
B_[4][1][138],
B_[4][2][138],
B_[5][0][138],
B_[5][1][138],
B_[5][2][138],
B_[6][0][138],
B_[6][1][138],
B_[6][2][138],
B_[7][0][138],
B_[7][1][138],
B_[7][2][138],
B_[8][0][138],
B_[8][1][138],
B_[8][2][138],
B_[9][0][138],
B_[9][1][138],
B_[9][2][138],
B_[10][0][138],
B_[10][1][138],
B_[10][2][138],
B_[11][0][138],
B_[11][1][138],
B_[11][2][138],
B_[12][0][138],
B_[12][1][138],
B_[12][2][138],
B_[13][0][138],
B_[13][1][138],
B_[13][2][138],
B_[14][0][138],
B_[14][1][138],
B_[14][2][138],
B_[15][0][138],
B_[15][1][138],
B_[15][2][138],
B_[0][0][139],
B_[0][1][139],
B_[0][2][139],
B_[1][0][139],
B_[1][1][139],
B_[1][2][139],
B_[2][0][139],
B_[2][1][139],
B_[2][2][139],
B_[3][0][139],
B_[3][1][139],
B_[3][2][139],
B_[4][0][139],
B_[4][1][139],
B_[4][2][139],
B_[5][0][139],
B_[5][1][139],
B_[5][2][139],
B_[6][0][139],
B_[6][1][139],
B_[6][2][139],
B_[7][0][139],
B_[7][1][139],
B_[7][2][139],
B_[8][0][139],
B_[8][1][139],
B_[8][2][139],
B_[9][0][139],
B_[9][1][139],
B_[9][2][139],
B_[10][0][139],
B_[10][1][139],
B_[10][2][139],
B_[11][0][139],
B_[11][1][139],
B_[11][2][139],
B_[12][0][139],
B_[12][1][139],
B_[12][2][139],
B_[13][0][139],
B_[13][1][139],
B_[13][2][139],
B_[14][0][139],
B_[14][1][139],
B_[14][2][139],
B_[15][0][139],
B_[15][1][139],
B_[15][2][139],
B_[0][0][140],
B_[0][1][140],
B_[0][2][140],
B_[1][0][140],
B_[1][1][140],
B_[1][2][140],
B_[2][0][140],
B_[2][1][140],
B_[2][2][140],
B_[3][0][140],
B_[3][1][140],
B_[3][2][140],
B_[4][0][140],
B_[4][1][140],
B_[4][2][140],
B_[5][0][140],
B_[5][1][140],
B_[5][2][140],
B_[6][0][140],
B_[6][1][140],
B_[6][2][140],
B_[7][0][140],
B_[7][1][140],
B_[7][2][140],
B_[8][0][140],
B_[8][1][140],
B_[8][2][140],
B_[9][0][140],
B_[9][1][140],
B_[9][2][140],
B_[10][0][140],
B_[10][1][140],
B_[10][2][140],
B_[11][0][140],
B_[11][1][140],
B_[11][2][140],
B_[12][0][140],
B_[12][1][140],
B_[12][2][140],
B_[13][0][140],
B_[13][1][140],
B_[13][2][140],
B_[14][0][140],
B_[14][1][140],
B_[14][2][140],
B_[15][0][140],
B_[15][1][140],
B_[15][2][140],
B_[0][0][141],
B_[0][1][141],
B_[0][2][141],
B_[1][0][141],
B_[1][1][141],
B_[1][2][141],
B_[2][0][141],
B_[2][1][141],
B_[2][2][141],
B_[3][0][141],
B_[3][1][141],
B_[3][2][141],
B_[4][0][141],
B_[4][1][141],
B_[4][2][141],
B_[5][0][141],
B_[5][1][141],
B_[5][2][141],
B_[6][0][141],
B_[6][1][141],
B_[6][2][141],
B_[7][0][141],
B_[7][1][141],
B_[7][2][141],
B_[8][0][141],
B_[8][1][141],
B_[8][2][141],
B_[9][0][141],
B_[9][1][141],
B_[9][2][141],
B_[10][0][141],
B_[10][1][141],
B_[10][2][141],
B_[11][0][141],
B_[11][1][141],
B_[11][2][141],
B_[12][0][141],
B_[12][1][141],
B_[12][2][141],
B_[13][0][141],
B_[13][1][141],
B_[13][2][141],
B_[14][0][141],
B_[14][1][141],
B_[14][2][141],
B_[15][0][141],
B_[15][1][141],
B_[15][2][141],
B_[0][0][142],
B_[0][1][142],
B_[0][2][142],
B_[1][0][142],
B_[1][1][142],
B_[1][2][142],
B_[2][0][142],
B_[2][1][142],
B_[2][2][142],
B_[3][0][142],
B_[3][1][142],
B_[3][2][142],
B_[4][0][142],
B_[4][1][142],
B_[4][2][142],
B_[5][0][142],
B_[5][1][142],
B_[5][2][142],
B_[6][0][142],
B_[6][1][142],
B_[6][2][142],
B_[7][0][142],
B_[7][1][142],
B_[7][2][142],
B_[8][0][142],
B_[8][1][142],
B_[8][2][142],
B_[9][0][142],
B_[9][1][142],
B_[9][2][142],
B_[10][0][142],
B_[10][1][142],
B_[10][2][142],
B_[11][0][142],
B_[11][1][142],
B_[11][2][142],
B_[12][0][142],
B_[12][1][142],
B_[12][2][142],
B_[13][0][142],
B_[13][1][142],
B_[13][2][142],
B_[14][0][142],
B_[14][1][142],
B_[14][2][142],
B_[15][0][142],
B_[15][1][142],
B_[15][2][142],
B_[0][0][143],
B_[0][1][143],
B_[0][2][143],
B_[1][0][143],
B_[1][1][143],
B_[1][2][143],
B_[2][0][143],
B_[2][1][143],
B_[2][2][143],
B_[3][0][143],
B_[3][1][143],
B_[3][2][143],
B_[4][0][143],
B_[4][1][143],
B_[4][2][143],
B_[5][0][143],
B_[5][1][143],
B_[5][2][143],
B_[6][0][143],
B_[6][1][143],
B_[6][2][143],
B_[7][0][143],
B_[7][1][143],
B_[7][2][143],
B_[8][0][143],
B_[8][1][143],
B_[8][2][143],
B_[9][0][143],
B_[9][1][143],
B_[9][2][143],
B_[10][0][143],
B_[10][1][143],
B_[10][2][143],
B_[11][0][143],
B_[11][1][143],
B_[11][2][143],
B_[12][0][143],
B_[12][1][143],
B_[12][2][143],
B_[13][0][143],
B_[13][1][143],
B_[13][2][143],
B_[14][0][143],
B_[14][1][143],
B_[14][2][143],
B_[15][0][143],
B_[15][1][143],
B_[15][2][143],
B_[0][0][144],
B_[0][1][144],
B_[0][2][144],
B_[1][0][144],
B_[1][1][144],
B_[1][2][144],
B_[2][0][144],
B_[2][1][144],
B_[2][2][144],
B_[3][0][144],
B_[3][1][144],
B_[3][2][144],
B_[4][0][144],
B_[4][1][144],
B_[4][2][144],
B_[5][0][144],
B_[5][1][144],
B_[5][2][144],
B_[6][0][144],
B_[6][1][144],
B_[6][2][144],
B_[7][0][144],
B_[7][1][144],
B_[7][2][144],
B_[8][0][144],
B_[8][1][144],
B_[8][2][144],
B_[9][0][144],
B_[9][1][144],
B_[9][2][144],
B_[10][0][144],
B_[10][1][144],
B_[10][2][144],
B_[11][0][144],
B_[11][1][144],
B_[11][2][144],
B_[12][0][144],
B_[12][1][144],
B_[12][2][144],
B_[13][0][144],
B_[13][1][144],
B_[13][2][144],
B_[14][0][144],
B_[14][1][144],
B_[14][2][144],
B_[15][0][144],
B_[15][1][144],
B_[15][2][144],
B_[0][0][145],
B_[0][1][145],
B_[0][2][145],
B_[1][0][145],
B_[1][1][145],
B_[1][2][145],
B_[2][0][145],
B_[2][1][145],
B_[2][2][145],
B_[3][0][145],
B_[3][1][145],
B_[3][2][145],
B_[4][0][145],
B_[4][1][145],
B_[4][2][145],
B_[5][0][145],
B_[5][1][145],
B_[5][2][145],
B_[6][0][145],
B_[6][1][145],
B_[6][2][145],
B_[7][0][145],
B_[7][1][145],
B_[7][2][145],
B_[8][0][145],
B_[8][1][145],
B_[8][2][145],
B_[9][0][145],
B_[9][1][145],
B_[9][2][145],
B_[10][0][145],
B_[10][1][145],
B_[10][2][145],
B_[11][0][145],
B_[11][1][145],
B_[11][2][145],
B_[12][0][145],
B_[12][1][145],
B_[12][2][145],
B_[13][0][145],
B_[13][1][145],
B_[13][2][145],
B_[14][0][145],
B_[14][1][145],
B_[14][2][145],
B_[15][0][145],
B_[15][1][145],
B_[15][2][145],
B_[0][0][146],
B_[0][1][146],
B_[0][2][146],
B_[1][0][146],
B_[1][1][146],
B_[1][2][146],
B_[2][0][146],
B_[2][1][146],
B_[2][2][146],
B_[3][0][146],
B_[3][1][146],
B_[3][2][146],
B_[4][0][146],
B_[4][1][146],
B_[4][2][146],
B_[5][0][146],
B_[5][1][146],
B_[5][2][146],
B_[6][0][146],
B_[6][1][146],
B_[6][2][146],
B_[7][0][146],
B_[7][1][146],
B_[7][2][146],
B_[8][0][146],
B_[8][1][146],
B_[8][2][146],
B_[9][0][146],
B_[9][1][146],
B_[9][2][146],
B_[10][0][146],
B_[10][1][146],
B_[10][2][146],
B_[11][0][146],
B_[11][1][146],
B_[11][2][146],
B_[12][0][146],
B_[12][1][146],
B_[12][2][146],
B_[13][0][146],
B_[13][1][146],
B_[13][2][146],
B_[14][0][146],
B_[14][1][146],
B_[14][2][146],
B_[15][0][146],
B_[15][1][146],
B_[15][2][146],
B_[0][0][147],
B_[0][1][147],
B_[0][2][147],
B_[1][0][147],
B_[1][1][147],
B_[1][2][147],
B_[2][0][147],
B_[2][1][147],
B_[2][2][147],
B_[3][0][147],
B_[3][1][147],
B_[3][2][147],
B_[4][0][147],
B_[4][1][147],
B_[4][2][147],
B_[5][0][147],
B_[5][1][147],
B_[5][2][147],
B_[6][0][147],
B_[6][1][147],
B_[6][2][147],
B_[7][0][147],
B_[7][1][147],
B_[7][2][147],
B_[8][0][147],
B_[8][1][147],
B_[8][2][147],
B_[9][0][147],
B_[9][1][147],
B_[9][2][147],
B_[10][0][147],
B_[10][1][147],
B_[10][2][147],
B_[11][0][147],
B_[11][1][147],
B_[11][2][147],
B_[12][0][147],
B_[12][1][147],
B_[12][2][147],
B_[13][0][147],
B_[13][1][147],
B_[13][2][147],
B_[14][0][147],
B_[14][1][147],
B_[14][2][147],
B_[15][0][147],
B_[15][1][147],
B_[15][2][147],
B_[0][0][148],
B_[0][1][148],
B_[0][2][148],
B_[1][0][148],
B_[1][1][148],
B_[1][2][148],
B_[2][0][148],
B_[2][1][148],
B_[2][2][148],
B_[3][0][148],
B_[3][1][148],
B_[3][2][148],
B_[4][0][148],
B_[4][1][148],
B_[4][2][148],
B_[5][0][148],
B_[5][1][148],
B_[5][2][148],
B_[6][0][148],
B_[6][1][148],
B_[6][2][148],
B_[7][0][148],
B_[7][1][148],
B_[7][2][148],
B_[8][0][148],
B_[8][1][148],
B_[8][2][148],
B_[9][0][148],
B_[9][1][148],
B_[9][2][148],
B_[10][0][148],
B_[10][1][148],
B_[10][2][148],
B_[11][0][148],
B_[11][1][148],
B_[11][2][148],
B_[12][0][148],
B_[12][1][148],
B_[12][2][148],
B_[13][0][148],
B_[13][1][148],
B_[13][2][148],
B_[14][0][148],
B_[14][1][148],
B_[14][2][148],
B_[15][0][148],
B_[15][1][148],
B_[15][2][148],
B_[0][0][149],
B_[0][1][149],
B_[0][2][149],
B_[1][0][149],
B_[1][1][149],
B_[1][2][149],
B_[2][0][149],
B_[2][1][149],
B_[2][2][149],
B_[3][0][149],
B_[3][1][149],
B_[3][2][149],
B_[4][0][149],
B_[4][1][149],
B_[4][2][149],
B_[5][0][149],
B_[5][1][149],
B_[5][2][149],
B_[6][0][149],
B_[6][1][149],
B_[6][2][149],
B_[7][0][149],
B_[7][1][149],
B_[7][2][149],
B_[8][0][149],
B_[8][1][149],
B_[8][2][149],
B_[9][0][149],
B_[9][1][149],
B_[9][2][149],
B_[10][0][149],
B_[10][1][149],
B_[10][2][149],
B_[11][0][149],
B_[11][1][149],
B_[11][2][149],
B_[12][0][149],
B_[12][1][149],
B_[12][2][149],
B_[13][0][149],
B_[13][1][149],
B_[13][2][149],
B_[14][0][149],
B_[14][1][149],
B_[14][2][149],
B_[15][0][149],
B_[15][1][149],
B_[15][2][149],
B_[0][0][150],
B_[0][1][150],
B_[0][2][150],
B_[1][0][150],
B_[1][1][150],
B_[1][2][150],
B_[2][0][150],
B_[2][1][150],
B_[2][2][150],
B_[3][0][150],
B_[3][1][150],
B_[3][2][150],
B_[4][0][150],
B_[4][1][150],
B_[4][2][150],
B_[5][0][150],
B_[5][1][150],
B_[5][2][150],
B_[6][0][150],
B_[6][1][150],
B_[6][2][150],
B_[7][0][150],
B_[7][1][150],
B_[7][2][150],
B_[8][0][150],
B_[8][1][150],
B_[8][2][150],
B_[9][0][150],
B_[9][1][150],
B_[9][2][150],
B_[10][0][150],
B_[10][1][150],
B_[10][2][150],
B_[11][0][150],
B_[11][1][150],
B_[11][2][150],
B_[12][0][150],
B_[12][1][150],
B_[12][2][150],
B_[13][0][150],
B_[13][1][150],
B_[13][2][150],
B_[14][0][150],
B_[14][1][150],
B_[14][2][150],
B_[15][0][150],
B_[15][1][150],
B_[15][2][150],
B_[0][0][151],
B_[0][1][151],
B_[0][2][151],
B_[1][0][151],
B_[1][1][151],
B_[1][2][151],
B_[2][0][151],
B_[2][1][151],
B_[2][2][151],
B_[3][0][151],
B_[3][1][151],
B_[3][2][151],
B_[4][0][151],
B_[4][1][151],
B_[4][2][151],
B_[5][0][151],
B_[5][1][151],
B_[5][2][151],
B_[6][0][151],
B_[6][1][151],
B_[6][2][151],
B_[7][0][151],
B_[7][1][151],
B_[7][2][151],
B_[8][0][151],
B_[8][1][151],
B_[8][2][151],
B_[9][0][151],
B_[9][1][151],
B_[9][2][151],
B_[10][0][151],
B_[10][1][151],
B_[10][2][151],
B_[11][0][151],
B_[11][1][151],
B_[11][2][151],
B_[12][0][151],
B_[12][1][151],
B_[12][2][151],
B_[13][0][151],
B_[13][1][151],
B_[13][2][151],
B_[14][0][151],
B_[14][1][151],
B_[14][2][151],
B_[15][0][151],
B_[15][1][151],
B_[15][2][151],
B_[0][0][152],
B_[0][1][152],
B_[0][2][152],
B_[1][0][152],
B_[1][1][152],
B_[1][2][152],
B_[2][0][152],
B_[2][1][152],
B_[2][2][152],
B_[3][0][152],
B_[3][1][152],
B_[3][2][152],
B_[4][0][152],
B_[4][1][152],
B_[4][2][152],
B_[5][0][152],
B_[5][1][152],
B_[5][2][152],
B_[6][0][152],
B_[6][1][152],
B_[6][2][152],
B_[7][0][152],
B_[7][1][152],
B_[7][2][152],
B_[8][0][152],
B_[8][1][152],
B_[8][2][152],
B_[9][0][152],
B_[9][1][152],
B_[9][2][152],
B_[10][0][152],
B_[10][1][152],
B_[10][2][152],
B_[11][0][152],
B_[11][1][152],
B_[11][2][152],
B_[12][0][152],
B_[12][1][152],
B_[12][2][152],
B_[13][0][152],
B_[13][1][152],
B_[13][2][152],
B_[14][0][152],
B_[14][1][152],
B_[14][2][152],
B_[15][0][152],
B_[15][1][152],
B_[15][2][152],
B_[0][0][153],
B_[0][1][153],
B_[0][2][153],
B_[1][0][153],
B_[1][1][153],
B_[1][2][153],
B_[2][0][153],
B_[2][1][153],
B_[2][2][153],
B_[3][0][153],
B_[3][1][153],
B_[3][2][153],
B_[4][0][153],
B_[4][1][153],
B_[4][2][153],
B_[5][0][153],
B_[5][1][153],
B_[5][2][153],
B_[6][0][153],
B_[6][1][153],
B_[6][2][153],
B_[7][0][153],
B_[7][1][153],
B_[7][2][153],
B_[8][0][153],
B_[8][1][153],
B_[8][2][153],
B_[9][0][153],
B_[9][1][153],
B_[9][2][153],
B_[10][0][153],
B_[10][1][153],
B_[10][2][153],
B_[11][0][153],
B_[11][1][153],
B_[11][2][153],
B_[12][0][153],
B_[12][1][153],
B_[12][2][153],
B_[13][0][153],
B_[13][1][153],
B_[13][2][153],
B_[14][0][153],
B_[14][1][153],
B_[14][2][153],
B_[15][0][153],
B_[15][1][153],
B_[15][2][153],
B_[0][0][154],
B_[0][1][154],
B_[0][2][154],
B_[1][0][154],
B_[1][1][154],
B_[1][2][154],
B_[2][0][154],
B_[2][1][154],
B_[2][2][154],
B_[3][0][154],
B_[3][1][154],
B_[3][2][154],
B_[4][0][154],
B_[4][1][154],
B_[4][2][154],
B_[5][0][154],
B_[5][1][154],
B_[5][2][154],
B_[6][0][154],
B_[6][1][154],
B_[6][2][154],
B_[7][0][154],
B_[7][1][154],
B_[7][2][154],
B_[8][0][154],
B_[8][1][154],
B_[8][2][154],
B_[9][0][154],
B_[9][1][154],
B_[9][2][154],
B_[10][0][154],
B_[10][1][154],
B_[10][2][154],
B_[11][0][154],
B_[11][1][154],
B_[11][2][154],
B_[12][0][154],
B_[12][1][154],
B_[12][2][154],
B_[13][0][154],
B_[13][1][154],
B_[13][2][154],
B_[14][0][154],
B_[14][1][154],
B_[14][2][154],
B_[15][0][154],
B_[15][1][154],
B_[15][2][154],
B_[0][0][155],
B_[0][1][155],
B_[0][2][155],
B_[1][0][155],
B_[1][1][155],
B_[1][2][155],
B_[2][0][155],
B_[2][1][155],
B_[2][2][155],
B_[3][0][155],
B_[3][1][155],
B_[3][2][155],
B_[4][0][155],
B_[4][1][155],
B_[4][2][155],
B_[5][0][155],
B_[5][1][155],
B_[5][2][155],
B_[6][0][155],
B_[6][1][155],
B_[6][2][155],
B_[7][0][155],
B_[7][1][155],
B_[7][2][155],
B_[8][0][155],
B_[8][1][155],
B_[8][2][155],
B_[9][0][155],
B_[9][1][155],
B_[9][2][155],
B_[10][0][155],
B_[10][1][155],
B_[10][2][155],
B_[11][0][155],
B_[11][1][155],
B_[11][2][155],
B_[12][0][155],
B_[12][1][155],
B_[12][2][155],
B_[13][0][155],
B_[13][1][155],
B_[13][2][155],
B_[14][0][155],
B_[14][1][155],
B_[14][2][155],
B_[15][0][155],
B_[15][1][155],
B_[15][2][155],
B_[0][0][156],
B_[0][1][156],
B_[0][2][156],
B_[1][0][156],
B_[1][1][156],
B_[1][2][156],
B_[2][0][156],
B_[2][1][156],
B_[2][2][156],
B_[3][0][156],
B_[3][1][156],
B_[3][2][156],
B_[4][0][156],
B_[4][1][156],
B_[4][2][156],
B_[5][0][156],
B_[5][1][156],
B_[5][2][156],
B_[6][0][156],
B_[6][1][156],
B_[6][2][156],
B_[7][0][156],
B_[7][1][156],
B_[7][2][156],
B_[8][0][156],
B_[8][1][156],
B_[8][2][156],
B_[9][0][156],
B_[9][1][156],
B_[9][2][156],
B_[10][0][156],
B_[10][1][156],
B_[10][2][156],
B_[11][0][156],
B_[11][1][156],
B_[11][2][156],
B_[12][0][156],
B_[12][1][156],
B_[12][2][156],
B_[13][0][156],
B_[13][1][156],
B_[13][2][156],
B_[14][0][156],
B_[14][1][156],
B_[14][2][156],
B_[15][0][156],
B_[15][1][156],
B_[15][2][156],
B_[0][0][157],
B_[0][1][157],
B_[0][2][157],
B_[1][0][157],
B_[1][1][157],
B_[1][2][157],
B_[2][0][157],
B_[2][1][157],
B_[2][2][157],
B_[3][0][157],
B_[3][1][157],
B_[3][2][157],
B_[4][0][157],
B_[4][1][157],
B_[4][2][157],
B_[5][0][157],
B_[5][1][157],
B_[5][2][157],
B_[6][0][157],
B_[6][1][157],
B_[6][2][157],
B_[7][0][157],
B_[7][1][157],
B_[7][2][157],
B_[8][0][157],
B_[8][1][157],
B_[8][2][157],
B_[9][0][157],
B_[9][1][157],
B_[9][2][157],
B_[10][0][157],
B_[10][1][157],
B_[10][2][157],
B_[11][0][157],
B_[11][1][157],
B_[11][2][157],
B_[12][0][157],
B_[12][1][157],
B_[12][2][157],
B_[13][0][157],
B_[13][1][157],
B_[13][2][157],
B_[14][0][157],
B_[14][1][157],
B_[14][2][157],
B_[15][0][157],
B_[15][1][157],
B_[15][2][157],
B_[0][0][158],
B_[0][1][158],
B_[0][2][158],
B_[1][0][158],
B_[1][1][158],
B_[1][2][158],
B_[2][0][158],
B_[2][1][158],
B_[2][2][158],
B_[3][0][158],
B_[3][1][158],
B_[3][2][158],
B_[4][0][158],
B_[4][1][158],
B_[4][2][158],
B_[5][0][158],
B_[5][1][158],
B_[5][2][158],
B_[6][0][158],
B_[6][1][158],
B_[6][2][158],
B_[7][0][158],
B_[7][1][158],
B_[7][2][158],
B_[8][0][158],
B_[8][1][158],
B_[8][2][158],
B_[9][0][158],
B_[9][1][158],
B_[9][2][158],
B_[10][0][158],
B_[10][1][158],
B_[10][2][158],
B_[11][0][158],
B_[11][1][158],
B_[11][2][158],
B_[12][0][158],
B_[12][1][158],
B_[12][2][158],
B_[13][0][158],
B_[13][1][158],
B_[13][2][158],
B_[14][0][158],
B_[14][1][158],
B_[14][2][158],
B_[15][0][158],
B_[15][1][158],
B_[15][2][158],
B_[0][0][159],
B_[0][1][159],
B_[0][2][159],
B_[1][0][159],
B_[1][1][159],
B_[1][2][159],
B_[2][0][159],
B_[2][1][159],
B_[2][2][159],
B_[3][0][159],
B_[3][1][159],
B_[3][2][159],
B_[4][0][159],
B_[4][1][159],
B_[4][2][159],
B_[5][0][159],
B_[5][1][159],
B_[5][2][159],
B_[6][0][159],
B_[6][1][159],
B_[6][2][159],
B_[7][0][159],
B_[7][1][159],
B_[7][2][159],
B_[8][0][159],
B_[8][1][159],
B_[8][2][159],
B_[9][0][159],
B_[9][1][159],
B_[9][2][159],
B_[10][0][159],
B_[10][1][159],
B_[10][2][159],
B_[11][0][159],
B_[11][1][159],
B_[11][2][159],
B_[12][0][159],
B_[12][1][159],
B_[12][2][159],
B_[13][0][159],
B_[13][1][159],
B_[13][2][159],
B_[14][0][159],
B_[14][1][159],
B_[14][2][159],
B_[15][0][159],
B_[15][1][159],
B_[15][2][159],
B_[0][0][160],
B_[0][1][160],
B_[0][2][160],
B_[1][0][160],
B_[1][1][160],
B_[1][2][160],
B_[2][0][160],
B_[2][1][160],
B_[2][2][160],
B_[3][0][160],
B_[3][1][160],
B_[3][2][160],
B_[4][0][160],
B_[4][1][160],
B_[4][2][160],
B_[5][0][160],
B_[5][1][160],
B_[5][2][160],
B_[6][0][160],
B_[6][1][160],
B_[6][2][160],
B_[7][0][160],
B_[7][1][160],
B_[7][2][160],
B_[8][0][160],
B_[8][1][160],
B_[8][2][160],
B_[9][0][160],
B_[9][1][160],
B_[9][2][160],
B_[10][0][160],
B_[10][1][160],
B_[10][2][160],
B_[11][0][160],
B_[11][1][160],
B_[11][2][160],
B_[12][0][160],
B_[12][1][160],
B_[12][2][160],
B_[13][0][160],
B_[13][1][160],
B_[13][2][160],
B_[14][0][160],
B_[14][1][160],
B_[14][2][160],
B_[15][0][160],
B_[15][1][160],
B_[15][2][160],
B_[0][0][161],
B_[0][1][161],
B_[0][2][161],
B_[1][0][161],
B_[1][1][161],
B_[1][2][161],
B_[2][0][161],
B_[2][1][161],
B_[2][2][161],
B_[3][0][161],
B_[3][1][161],
B_[3][2][161],
B_[4][0][161],
B_[4][1][161],
B_[4][2][161],
B_[5][0][161],
B_[5][1][161],
B_[5][2][161],
B_[6][0][161],
B_[6][1][161],
B_[6][2][161],
B_[7][0][161],
B_[7][1][161],
B_[7][2][161],
B_[8][0][161],
B_[8][1][161],
B_[8][2][161],
B_[9][0][161],
B_[9][1][161],
B_[9][2][161],
B_[10][0][161],
B_[10][1][161],
B_[10][2][161],
B_[11][0][161],
B_[11][1][161],
B_[11][2][161],
B_[12][0][161],
B_[12][1][161],
B_[12][2][161],
B_[13][0][161],
B_[13][1][161],
B_[13][2][161],
B_[14][0][161],
B_[14][1][161],
B_[14][2][161],
B_[15][0][161],
B_[15][1][161],
B_[15][2][161],
B_[0][0][162],
B_[0][1][162],
B_[0][2][162],
B_[1][0][162],
B_[1][1][162],
B_[1][2][162],
B_[2][0][162],
B_[2][1][162],
B_[2][2][162],
B_[3][0][162],
B_[3][1][162],
B_[3][2][162],
B_[4][0][162],
B_[4][1][162],
B_[4][2][162],
B_[5][0][162],
B_[5][1][162],
B_[5][2][162],
B_[6][0][162],
B_[6][1][162],
B_[6][2][162],
B_[7][0][162],
B_[7][1][162],
B_[7][2][162],
B_[8][0][162],
B_[8][1][162],
B_[8][2][162],
B_[9][0][162],
B_[9][1][162],
B_[9][2][162],
B_[10][0][162],
B_[10][1][162],
B_[10][2][162],
B_[11][0][162],
B_[11][1][162],
B_[11][2][162],
B_[12][0][162],
B_[12][1][162],
B_[12][2][162],
B_[13][0][162],
B_[13][1][162],
B_[13][2][162],
B_[14][0][162],
B_[14][1][162],
B_[14][2][162],
B_[15][0][162],
B_[15][1][162],
B_[15][2][162],
B_[0][0][163],
B_[0][1][163],
B_[0][2][163],
B_[1][0][163],
B_[1][1][163],
B_[1][2][163],
B_[2][0][163],
B_[2][1][163],
B_[2][2][163],
B_[3][0][163],
B_[3][1][163],
B_[3][2][163],
B_[4][0][163],
B_[4][1][163],
B_[4][2][163],
B_[5][0][163],
B_[5][1][163],
B_[5][2][163],
B_[6][0][163],
B_[6][1][163],
B_[6][2][163],
B_[7][0][163],
B_[7][1][163],
B_[7][2][163],
B_[8][0][163],
B_[8][1][163],
B_[8][2][163],
B_[9][0][163],
B_[9][1][163],
B_[9][2][163],
B_[10][0][163],
B_[10][1][163],
B_[10][2][163],
B_[11][0][163],
B_[11][1][163],
B_[11][2][163],
B_[12][0][163],
B_[12][1][163],
B_[12][2][163],
B_[13][0][163],
B_[13][1][163],
B_[13][2][163],
B_[14][0][163],
B_[14][1][163],
B_[14][2][163],
B_[15][0][163],
B_[15][1][163],
B_[15][2][163],
B_[0][0][164],
B_[0][1][164],
B_[0][2][164],
B_[1][0][164],
B_[1][1][164],
B_[1][2][164],
B_[2][0][164],
B_[2][1][164],
B_[2][2][164],
B_[3][0][164],
B_[3][1][164],
B_[3][2][164],
B_[4][0][164],
B_[4][1][164],
B_[4][2][164],
B_[5][0][164],
B_[5][1][164],
B_[5][2][164],
B_[6][0][164],
B_[6][1][164],
B_[6][2][164],
B_[7][0][164],
B_[7][1][164],
B_[7][2][164],
B_[8][0][164],
B_[8][1][164],
B_[8][2][164],
B_[9][0][164],
B_[9][1][164],
B_[9][2][164],
B_[10][0][164],
B_[10][1][164],
B_[10][2][164],
B_[11][0][164],
B_[11][1][164],
B_[11][2][164],
B_[12][0][164],
B_[12][1][164],
B_[12][2][164],
B_[13][0][164],
B_[13][1][164],
B_[13][2][164],
B_[14][0][164],
B_[14][1][164],
B_[14][2][164],
B_[15][0][164],
B_[15][1][164],
B_[15][2][164],
B_[0][0][165],
B_[0][1][165],
B_[0][2][165],
B_[1][0][165],
B_[1][1][165],
B_[1][2][165],
B_[2][0][165],
B_[2][1][165],
B_[2][2][165],
B_[3][0][165],
B_[3][1][165],
B_[3][2][165],
B_[4][0][165],
B_[4][1][165],
B_[4][2][165],
B_[5][0][165],
B_[5][1][165],
B_[5][2][165],
B_[6][0][165],
B_[6][1][165],
B_[6][2][165],
B_[7][0][165],
B_[7][1][165],
B_[7][2][165],
B_[8][0][165],
B_[8][1][165],
B_[8][2][165],
B_[9][0][165],
B_[9][1][165],
B_[9][2][165],
B_[10][0][165],
B_[10][1][165],
B_[10][2][165],
B_[11][0][165],
B_[11][1][165],
B_[11][2][165],
B_[12][0][165],
B_[12][1][165],
B_[12][2][165],
B_[13][0][165],
B_[13][1][165],
B_[13][2][165],
B_[14][0][165],
B_[14][1][165],
B_[14][2][165],
B_[15][0][165],
B_[15][1][165],
B_[15][2][165],
B_[0][0][166],
B_[0][1][166],
B_[0][2][166],
B_[1][0][166],
B_[1][1][166],
B_[1][2][166],
B_[2][0][166],
B_[2][1][166],
B_[2][2][166],
B_[3][0][166],
B_[3][1][166],
B_[3][2][166],
B_[4][0][166],
B_[4][1][166],
B_[4][2][166],
B_[5][0][166],
B_[5][1][166],
B_[5][2][166],
B_[6][0][166],
B_[6][1][166],
B_[6][2][166],
B_[7][0][166],
B_[7][1][166],
B_[7][2][166],
B_[8][0][166],
B_[8][1][166],
B_[8][2][166],
B_[9][0][166],
B_[9][1][166],
B_[9][2][166],
B_[10][0][166],
B_[10][1][166],
B_[10][2][166],
B_[11][0][166],
B_[11][1][166],
B_[11][2][166],
B_[12][0][166],
B_[12][1][166],
B_[12][2][166],
B_[13][0][166],
B_[13][1][166],
B_[13][2][166],
B_[14][0][166],
B_[14][1][166],
B_[14][2][166],
B_[15][0][166],
B_[15][1][166],
B_[15][2][166],
B_[0][0][167],
B_[0][1][167],
B_[0][2][167],
B_[1][0][167],
B_[1][1][167],
B_[1][2][167],
B_[2][0][167],
B_[2][1][167],
B_[2][2][167],
B_[3][0][167],
B_[3][1][167],
B_[3][2][167],
B_[4][0][167],
B_[4][1][167],
B_[4][2][167],
B_[5][0][167],
B_[5][1][167],
B_[5][2][167],
B_[6][0][167],
B_[6][1][167],
B_[6][2][167],
B_[7][0][167],
B_[7][1][167],
B_[7][2][167],
B_[8][0][167],
B_[8][1][167],
B_[8][2][167],
B_[9][0][167],
B_[9][1][167],
B_[9][2][167],
B_[10][0][167],
B_[10][1][167],
B_[10][2][167],
B_[11][0][167],
B_[11][1][167],
B_[11][2][167],
B_[12][0][167],
B_[12][1][167],
B_[12][2][167],
B_[13][0][167],
B_[13][1][167],
B_[13][2][167],
B_[14][0][167],
B_[14][1][167],
B_[14][2][167],
B_[15][0][167],
B_[15][1][167],
B_[15][2][167],
B_[0][0][168],
B_[0][1][168],
B_[0][2][168],
B_[1][0][168],
B_[1][1][168],
B_[1][2][168],
B_[2][0][168],
B_[2][1][168],
B_[2][2][168],
B_[3][0][168],
B_[3][1][168],
B_[3][2][168],
B_[4][0][168],
B_[4][1][168],
B_[4][2][168],
B_[5][0][168],
B_[5][1][168],
B_[5][2][168],
B_[6][0][168],
B_[6][1][168],
B_[6][2][168],
B_[7][0][168],
B_[7][1][168],
B_[7][2][168],
B_[8][0][168],
B_[8][1][168],
B_[8][2][168],
B_[9][0][168],
B_[9][1][168],
B_[9][2][168],
B_[10][0][168],
B_[10][1][168],
B_[10][2][168],
B_[11][0][168],
B_[11][1][168],
B_[11][2][168],
B_[12][0][168],
B_[12][1][168],
B_[12][2][168],
B_[13][0][168],
B_[13][1][168],
B_[13][2][168],
B_[14][0][168],
B_[14][1][168],
B_[14][2][168],
B_[15][0][168],
B_[15][1][168],
B_[15][2][168],
B_[0][0][169],
B_[0][1][169],
B_[0][2][169],
B_[1][0][169],
B_[1][1][169],
B_[1][2][169],
B_[2][0][169],
B_[2][1][169],
B_[2][2][169],
B_[3][0][169],
B_[3][1][169],
B_[3][2][169],
B_[4][0][169],
B_[4][1][169],
B_[4][2][169],
B_[5][0][169],
B_[5][1][169],
B_[5][2][169],
B_[6][0][169],
B_[6][1][169],
B_[6][2][169],
B_[7][0][169],
B_[7][1][169],
B_[7][2][169],
B_[8][0][169],
B_[8][1][169],
B_[8][2][169],
B_[9][0][169],
B_[9][1][169],
B_[9][2][169],
B_[10][0][169],
B_[10][1][169],
B_[10][2][169],
B_[11][0][169],
B_[11][1][169],
B_[11][2][169],
B_[12][0][169],
B_[12][1][169],
B_[12][2][169],
B_[13][0][169],
B_[13][1][169],
B_[13][2][169],
B_[14][0][169],
B_[14][1][169],
B_[14][2][169],
B_[15][0][169],
B_[15][1][169],
B_[15][2][169],
B_[0][0][170],
B_[0][1][170],
B_[0][2][170],
B_[1][0][170],
B_[1][1][170],
B_[1][2][170],
B_[2][0][170],
B_[2][1][170],
B_[2][2][170],
B_[3][0][170],
B_[3][1][170],
B_[3][2][170],
B_[4][0][170],
B_[4][1][170],
B_[4][2][170],
B_[5][0][170],
B_[5][1][170],
B_[5][2][170],
B_[6][0][170],
B_[6][1][170],
B_[6][2][170],
B_[7][0][170],
B_[7][1][170],
B_[7][2][170],
B_[8][0][170],
B_[8][1][170],
B_[8][2][170],
B_[9][0][170],
B_[9][1][170],
B_[9][2][170],
B_[10][0][170],
B_[10][1][170],
B_[10][2][170],
B_[11][0][170],
B_[11][1][170],
B_[11][2][170],
B_[12][0][170],
B_[12][1][170],
B_[12][2][170],
B_[13][0][170],
B_[13][1][170],
B_[13][2][170],
B_[14][0][170],
B_[14][1][170],
B_[14][2][170],
B_[15][0][170],
B_[15][1][170],
B_[15][2][170],
B_[0][0][171],
B_[0][1][171],
B_[0][2][171],
B_[1][0][171],
B_[1][1][171],
B_[1][2][171],
B_[2][0][171],
B_[2][1][171],
B_[2][2][171],
B_[3][0][171],
B_[3][1][171],
B_[3][2][171],
B_[4][0][171],
B_[4][1][171],
B_[4][2][171],
B_[5][0][171],
B_[5][1][171],
B_[5][2][171],
B_[6][0][171],
B_[6][1][171],
B_[6][2][171],
B_[7][0][171],
B_[7][1][171],
B_[7][2][171],
B_[8][0][171],
B_[8][1][171],
B_[8][2][171],
B_[9][0][171],
B_[9][1][171],
B_[9][2][171],
B_[10][0][171],
B_[10][1][171],
B_[10][2][171],
B_[11][0][171],
B_[11][1][171],
B_[11][2][171],
B_[12][0][171],
B_[12][1][171],
B_[12][2][171],
B_[13][0][171],
B_[13][1][171],
B_[13][2][171],
B_[14][0][171],
B_[14][1][171],
B_[14][2][171],
B_[15][0][171],
B_[15][1][171],
B_[15][2][171],
B_[0][0][172],
B_[0][1][172],
B_[0][2][172],
B_[1][0][172],
B_[1][1][172],
B_[1][2][172],
B_[2][0][172],
B_[2][1][172],
B_[2][2][172],
B_[3][0][172],
B_[3][1][172],
B_[3][2][172],
B_[4][0][172],
B_[4][1][172],
B_[4][2][172],
B_[5][0][172],
B_[5][1][172],
B_[5][2][172],
B_[6][0][172],
B_[6][1][172],
B_[6][2][172],
B_[7][0][172],
B_[7][1][172],
B_[7][2][172],
B_[8][0][172],
B_[8][1][172],
B_[8][2][172],
B_[9][0][172],
B_[9][1][172],
B_[9][2][172],
B_[10][0][172],
B_[10][1][172],
B_[10][2][172],
B_[11][0][172],
B_[11][1][172],
B_[11][2][172],
B_[12][0][172],
B_[12][1][172],
B_[12][2][172],
B_[13][0][172],
B_[13][1][172],
B_[13][2][172],
B_[14][0][172],
B_[14][1][172],
B_[14][2][172],
B_[15][0][172],
B_[15][1][172],
B_[15][2][172],
B_[0][0][173],
B_[0][1][173],
B_[0][2][173],
B_[1][0][173],
B_[1][1][173],
B_[1][2][173],
B_[2][0][173],
B_[2][1][173],
B_[2][2][173],
B_[3][0][173],
B_[3][1][173],
B_[3][2][173],
B_[4][0][173],
B_[4][1][173],
B_[4][2][173],
B_[5][0][173],
B_[5][1][173],
B_[5][2][173],
B_[6][0][173],
B_[6][1][173],
B_[6][2][173],
B_[7][0][173],
B_[7][1][173],
B_[7][2][173],
B_[8][0][173],
B_[8][1][173],
B_[8][2][173],
B_[9][0][173],
B_[9][1][173],
B_[9][2][173],
B_[10][0][173],
B_[10][1][173],
B_[10][2][173],
B_[11][0][173],
B_[11][1][173],
B_[11][2][173],
B_[12][0][173],
B_[12][1][173],
B_[12][2][173],
B_[13][0][173],
B_[13][1][173],
B_[13][2][173],
B_[14][0][173],
B_[14][1][173],
B_[14][2][173],
B_[15][0][173],
B_[15][1][173],
B_[15][2][173],
B_[0][0][174],
B_[0][1][174],
B_[0][2][174],
B_[1][0][174],
B_[1][1][174],
B_[1][2][174],
B_[2][0][174],
B_[2][1][174],
B_[2][2][174],
B_[3][0][174],
B_[3][1][174],
B_[3][2][174],
B_[4][0][174],
B_[4][1][174],
B_[4][2][174],
B_[5][0][174],
B_[5][1][174],
B_[5][2][174],
B_[6][0][174],
B_[6][1][174],
B_[6][2][174],
B_[7][0][174],
B_[7][1][174],
B_[7][2][174],
B_[8][0][174],
B_[8][1][174],
B_[8][2][174],
B_[9][0][174],
B_[9][1][174],
B_[9][2][174],
B_[10][0][174],
B_[10][1][174],
B_[10][2][174],
B_[11][0][174],
B_[11][1][174],
B_[11][2][174],
B_[12][0][174],
B_[12][1][174],
B_[12][2][174],
B_[13][0][174],
B_[13][1][174],
B_[13][2][174],
B_[14][0][174],
B_[14][1][174],
B_[14][2][174],
B_[15][0][174],
B_[15][1][174],
B_[15][2][174],
B_[0][0][175],
B_[0][1][175],
B_[0][2][175],
B_[1][0][175],
B_[1][1][175],
B_[1][2][175],
B_[2][0][175],
B_[2][1][175],
B_[2][2][175],
B_[3][0][175],
B_[3][1][175],
B_[3][2][175],
B_[4][0][175],
B_[4][1][175],
B_[4][2][175],
B_[5][0][175],
B_[5][1][175],
B_[5][2][175],
B_[6][0][175],
B_[6][1][175],
B_[6][2][175],
B_[7][0][175],
B_[7][1][175],
B_[7][2][175],
B_[8][0][175],
B_[8][1][175],
B_[8][2][175],
B_[9][0][175],
B_[9][1][175],
B_[9][2][175],
B_[10][0][175],
B_[10][1][175],
B_[10][2][175],
B_[11][0][175],
B_[11][1][175],
B_[11][2][175],
B_[12][0][175],
B_[12][1][175],
B_[12][2][175],
B_[13][0][175],
B_[13][1][175],
B_[13][2][175],
B_[14][0][175],
B_[14][1][175],
B_[14][2][175],
B_[15][0][175],
B_[15][1][175],
B_[15][2][175],
B_[0][0][176],
B_[0][1][176],
B_[0][2][176],
B_[1][0][176],
B_[1][1][176],
B_[1][2][176],
B_[2][0][176],
B_[2][1][176],
B_[2][2][176],
B_[3][0][176],
B_[3][1][176],
B_[3][2][176],
B_[4][0][176],
B_[4][1][176],
B_[4][2][176],
B_[5][0][176],
B_[5][1][176],
B_[5][2][176],
B_[6][0][176],
B_[6][1][176],
B_[6][2][176],
B_[7][0][176],
B_[7][1][176],
B_[7][2][176],
B_[8][0][176],
B_[8][1][176],
B_[8][2][176],
B_[9][0][176],
B_[9][1][176],
B_[9][2][176],
B_[10][0][176],
B_[10][1][176],
B_[10][2][176],
B_[11][0][176],
B_[11][1][176],
B_[11][2][176],
B_[12][0][176],
B_[12][1][176],
B_[12][2][176],
B_[13][0][176],
B_[13][1][176],
B_[13][2][176],
B_[14][0][176],
B_[14][1][176],
B_[14][2][176],
B_[15][0][176],
B_[15][1][176],
B_[15][2][176],
B_[0][0][177],
B_[0][1][177],
B_[0][2][177],
B_[1][0][177],
B_[1][1][177],
B_[1][2][177],
B_[2][0][177],
B_[2][1][177],
B_[2][2][177],
B_[3][0][177],
B_[3][1][177],
B_[3][2][177],
B_[4][0][177],
B_[4][1][177],
B_[4][2][177],
B_[5][0][177],
B_[5][1][177],
B_[5][2][177],
B_[6][0][177],
B_[6][1][177],
B_[6][2][177],
B_[7][0][177],
B_[7][1][177],
B_[7][2][177],
B_[8][0][177],
B_[8][1][177],
B_[8][2][177],
B_[9][0][177],
B_[9][1][177],
B_[9][2][177],
B_[10][0][177],
B_[10][1][177],
B_[10][2][177],
B_[11][0][177],
B_[11][1][177],
B_[11][2][177],
B_[12][0][177],
B_[12][1][177],
B_[12][2][177],
B_[13][0][177],
B_[13][1][177],
B_[13][2][177],
B_[14][0][177],
B_[14][1][177],
B_[14][2][177],
B_[15][0][177],
B_[15][1][177],
B_[15][2][177],
B_[0][0][178],
B_[0][1][178],
B_[0][2][178],
B_[1][0][178],
B_[1][1][178],
B_[1][2][178],
B_[2][0][178],
B_[2][1][178],
B_[2][2][178],
B_[3][0][178],
B_[3][1][178],
B_[3][2][178],
B_[4][0][178],
B_[4][1][178],
B_[4][2][178],
B_[5][0][178],
B_[5][1][178],
B_[5][2][178],
B_[6][0][178],
B_[6][1][178],
B_[6][2][178],
B_[7][0][178],
B_[7][1][178],
B_[7][2][178],
B_[8][0][178],
B_[8][1][178],
B_[8][2][178],
B_[9][0][178],
B_[9][1][178],
B_[9][2][178],
B_[10][0][178],
B_[10][1][178],
B_[10][2][178],
B_[11][0][178],
B_[11][1][178],
B_[11][2][178],
B_[12][0][178],
B_[12][1][178],
B_[12][2][178],
B_[13][0][178],
B_[13][1][178],
B_[13][2][178],
B_[14][0][178],
B_[14][1][178],
B_[14][2][178],
B_[15][0][178],
B_[15][1][178],
B_[15][2][178],
B_[0][0][179],
B_[0][1][179],
B_[0][2][179],
B_[1][0][179],
B_[1][1][179],
B_[1][2][179],
B_[2][0][179],
B_[2][1][179],
B_[2][2][179],
B_[3][0][179],
B_[3][1][179],
B_[3][2][179],
B_[4][0][179],
B_[4][1][179],
B_[4][2][179],
B_[5][0][179],
B_[5][1][179],
B_[5][2][179],
B_[6][0][179],
B_[6][1][179],
B_[6][2][179],
B_[7][0][179],
B_[7][1][179],
B_[7][2][179],
B_[8][0][179],
B_[8][1][179],
B_[8][2][179],
B_[9][0][179],
B_[9][1][179],
B_[9][2][179],
B_[10][0][179],
B_[10][1][179],
B_[10][2][179],
B_[11][0][179],
B_[11][1][179],
B_[11][2][179],
B_[12][0][179],
B_[12][1][179],
B_[12][2][179],
B_[13][0][179],
B_[13][1][179],
B_[13][2][179],
B_[14][0][179],
B_[14][1][179],
B_[14][2][179],
B_[15][0][179],
B_[15][1][179],
B_[15][2][179],
B_[0][0][180],
B_[0][1][180],
B_[0][2][180],
B_[1][0][180],
B_[1][1][180],
B_[1][2][180],
B_[2][0][180],
B_[2][1][180],
B_[2][2][180],
B_[3][0][180],
B_[3][1][180],
B_[3][2][180],
B_[4][0][180],
B_[4][1][180],
B_[4][2][180],
B_[5][0][180],
B_[5][1][180],
B_[5][2][180],
B_[6][0][180],
B_[6][1][180],
B_[6][2][180],
B_[7][0][180],
B_[7][1][180],
B_[7][2][180],
B_[8][0][180],
B_[8][1][180],
B_[8][2][180],
B_[9][0][180],
B_[9][1][180],
B_[9][2][180],
B_[10][0][180],
B_[10][1][180],
B_[10][2][180],
B_[11][0][180],
B_[11][1][180],
B_[11][2][180],
B_[12][0][180],
B_[12][1][180],
B_[12][2][180],
B_[13][0][180],
B_[13][1][180],
B_[13][2][180],
B_[14][0][180],
B_[14][1][180],
B_[14][2][180],
B_[15][0][180],
B_[15][1][180],
B_[15][2][180],
B_[0][0][181],
B_[0][1][181],
B_[0][2][181],
B_[1][0][181],
B_[1][1][181],
B_[1][2][181],
B_[2][0][181],
B_[2][1][181],
B_[2][2][181],
B_[3][0][181],
B_[3][1][181],
B_[3][2][181],
B_[4][0][181],
B_[4][1][181],
B_[4][2][181],
B_[5][0][181],
B_[5][1][181],
B_[5][2][181],
B_[6][0][181],
B_[6][1][181],
B_[6][2][181],
B_[7][0][181],
B_[7][1][181],
B_[7][2][181],
B_[8][0][181],
B_[8][1][181],
B_[8][2][181],
B_[9][0][181],
B_[9][1][181],
B_[9][2][181],
B_[10][0][181],
B_[10][1][181],
B_[10][2][181],
B_[11][0][181],
B_[11][1][181],
B_[11][2][181],
B_[12][0][181],
B_[12][1][181],
B_[12][2][181],
B_[13][0][181],
B_[13][1][181],
B_[13][2][181],
B_[14][0][181],
B_[14][1][181],
B_[14][2][181],
B_[15][0][181],
B_[15][1][181],
B_[15][2][181],
B_[0][0][182],
B_[0][1][182],
B_[0][2][182],
B_[1][0][182],
B_[1][1][182],
B_[1][2][182],
B_[2][0][182],
B_[2][1][182],
B_[2][2][182],
B_[3][0][182],
B_[3][1][182],
B_[3][2][182],
B_[4][0][182],
B_[4][1][182],
B_[4][2][182],
B_[5][0][182],
B_[5][1][182],
B_[5][2][182],
B_[6][0][182],
B_[6][1][182],
B_[6][2][182],
B_[7][0][182],
B_[7][1][182],
B_[7][2][182],
B_[8][0][182],
B_[8][1][182],
B_[8][2][182],
B_[9][0][182],
B_[9][1][182],
B_[9][2][182],
B_[10][0][182],
B_[10][1][182],
B_[10][2][182],
B_[11][0][182],
B_[11][1][182],
B_[11][2][182],
B_[12][0][182],
B_[12][1][182],
B_[12][2][182],
B_[13][0][182],
B_[13][1][182],
B_[13][2][182],
B_[14][0][182],
B_[14][1][182],
B_[14][2][182],
B_[15][0][182],
B_[15][1][182],
B_[15][2][182],
B_[0][0][183],
B_[0][1][183],
B_[0][2][183],
B_[1][0][183],
B_[1][1][183],
B_[1][2][183],
B_[2][0][183],
B_[2][1][183],
B_[2][2][183],
B_[3][0][183],
B_[3][1][183],
B_[3][2][183],
B_[4][0][183],
B_[4][1][183],
B_[4][2][183],
B_[5][0][183],
B_[5][1][183],
B_[5][2][183],
B_[6][0][183],
B_[6][1][183],
B_[6][2][183],
B_[7][0][183],
B_[7][1][183],
B_[7][2][183],
B_[8][0][183],
B_[8][1][183],
B_[8][2][183],
B_[9][0][183],
B_[9][1][183],
B_[9][2][183],
B_[10][0][183],
B_[10][1][183],
B_[10][2][183],
B_[11][0][183],
B_[11][1][183],
B_[11][2][183],
B_[12][0][183],
B_[12][1][183],
B_[12][2][183],
B_[13][0][183],
B_[13][1][183],
B_[13][2][183],
B_[14][0][183],
B_[14][1][183],
B_[14][2][183],
B_[15][0][183],
B_[15][1][183],
B_[15][2][183],
B_[0][0][184],
B_[0][1][184],
B_[0][2][184],
B_[1][0][184],
B_[1][1][184],
B_[1][2][184],
B_[2][0][184],
B_[2][1][184],
B_[2][2][184],
B_[3][0][184],
B_[3][1][184],
B_[3][2][184],
B_[4][0][184],
B_[4][1][184],
B_[4][2][184],
B_[5][0][184],
B_[5][1][184],
B_[5][2][184],
B_[6][0][184],
B_[6][1][184],
B_[6][2][184],
B_[7][0][184],
B_[7][1][184],
B_[7][2][184],
B_[8][0][184],
B_[8][1][184],
B_[8][2][184],
B_[9][0][184],
B_[9][1][184],
B_[9][2][184],
B_[10][0][184],
B_[10][1][184],
B_[10][2][184],
B_[11][0][184],
B_[11][1][184],
B_[11][2][184],
B_[12][0][184],
B_[12][1][184],
B_[12][2][184],
B_[13][0][184],
B_[13][1][184],
B_[13][2][184],
B_[14][0][184],
B_[14][1][184],
B_[14][2][184],
B_[15][0][184],
B_[15][1][184],
B_[15][2][184],
B_[0][0][185],
B_[0][1][185],
B_[0][2][185],
B_[1][0][185],
B_[1][1][185],
B_[1][2][185],
B_[2][0][185],
B_[2][1][185],
B_[2][2][185],
B_[3][0][185],
B_[3][1][185],
B_[3][2][185],
B_[4][0][185],
B_[4][1][185],
B_[4][2][185],
B_[5][0][185],
B_[5][1][185],
B_[5][2][185],
B_[6][0][185],
B_[6][1][185],
B_[6][2][185],
B_[7][0][185],
B_[7][1][185],
B_[7][2][185],
B_[8][0][185],
B_[8][1][185],
B_[8][2][185],
B_[9][0][185],
B_[9][1][185],
B_[9][2][185],
B_[10][0][185],
B_[10][1][185],
B_[10][2][185],
B_[11][0][185],
B_[11][1][185],
B_[11][2][185],
B_[12][0][185],
B_[12][1][185],
B_[12][2][185],
B_[13][0][185],
B_[13][1][185],
B_[13][2][185],
B_[14][0][185],
B_[14][1][185],
B_[14][2][185],
B_[15][0][185],
B_[15][1][185],
B_[15][2][185],
B_[0][0][186],
B_[0][1][186],
B_[0][2][186],
B_[1][0][186],
B_[1][1][186],
B_[1][2][186],
B_[2][0][186],
B_[2][1][186],
B_[2][2][186],
B_[3][0][186],
B_[3][1][186],
B_[3][2][186],
B_[4][0][186],
B_[4][1][186],
B_[4][2][186],
B_[5][0][186],
B_[5][1][186],
B_[5][2][186],
B_[6][0][186],
B_[6][1][186],
B_[6][2][186],
B_[7][0][186],
B_[7][1][186],
B_[7][2][186],
B_[8][0][186],
B_[8][1][186],
B_[8][2][186],
B_[9][0][186],
B_[9][1][186],
B_[9][2][186],
B_[10][0][186],
B_[10][1][186],
B_[10][2][186],
B_[11][0][186],
B_[11][1][186],
B_[11][2][186],
B_[12][0][186],
B_[12][1][186],
B_[12][2][186],
B_[13][0][186],
B_[13][1][186],
B_[13][2][186],
B_[14][0][186],
B_[14][1][186],
B_[14][2][186],
B_[15][0][186],
B_[15][1][186],
B_[15][2][186],
B_[0][0][187],
B_[0][1][187],
B_[0][2][187],
B_[1][0][187],
B_[1][1][187],
B_[1][2][187],
B_[2][0][187],
B_[2][1][187],
B_[2][2][187],
B_[3][0][187],
B_[3][1][187],
B_[3][2][187],
B_[4][0][187],
B_[4][1][187],
B_[4][2][187],
B_[5][0][187],
B_[5][1][187],
B_[5][2][187],
B_[6][0][187],
B_[6][1][187],
B_[6][2][187],
B_[7][0][187],
B_[7][1][187],
B_[7][2][187],
B_[8][0][187],
B_[8][1][187],
B_[8][2][187],
B_[9][0][187],
B_[9][1][187],
B_[9][2][187],
B_[10][0][187],
B_[10][1][187],
B_[10][2][187],
B_[11][0][187],
B_[11][1][187],
B_[11][2][187],
B_[12][0][187],
B_[12][1][187],
B_[12][2][187],
B_[13][0][187],
B_[13][1][187],
B_[13][2][187],
B_[14][0][187],
B_[14][1][187],
B_[14][2][187],
B_[15][0][187],
B_[15][1][187],
B_[15][2][187],
B_[0][0][188],
B_[0][1][188],
B_[0][2][188],
B_[1][0][188],
B_[1][1][188],
B_[1][2][188],
B_[2][0][188],
B_[2][1][188],
B_[2][2][188],
B_[3][0][188],
B_[3][1][188],
B_[3][2][188],
B_[4][0][188],
B_[4][1][188],
B_[4][2][188],
B_[5][0][188],
B_[5][1][188],
B_[5][2][188],
B_[6][0][188],
B_[6][1][188],
B_[6][2][188],
B_[7][0][188],
B_[7][1][188],
B_[7][2][188],
B_[8][0][188],
B_[8][1][188],
B_[8][2][188],
B_[9][0][188],
B_[9][1][188],
B_[9][2][188],
B_[10][0][188],
B_[10][1][188],
B_[10][2][188],
B_[11][0][188],
B_[11][1][188],
B_[11][2][188],
B_[12][0][188],
B_[12][1][188],
B_[12][2][188],
B_[13][0][188],
B_[13][1][188],
B_[13][2][188],
B_[14][0][188],
B_[14][1][188],
B_[14][2][188],
B_[15][0][188],
B_[15][1][188],
B_[15][2][188],
B_[0][0][189],
B_[0][1][189],
B_[0][2][189],
B_[1][0][189],
B_[1][1][189],
B_[1][2][189],
B_[2][0][189],
B_[2][1][189],
B_[2][2][189],
B_[3][0][189],
B_[3][1][189],
B_[3][2][189],
B_[4][0][189],
B_[4][1][189],
B_[4][2][189],
B_[5][0][189],
B_[5][1][189],
B_[5][2][189],
B_[6][0][189],
B_[6][1][189],
B_[6][2][189],
B_[7][0][189],
B_[7][1][189],
B_[7][2][189],
B_[8][0][189],
B_[8][1][189],
B_[8][2][189],
B_[9][0][189],
B_[9][1][189],
B_[9][2][189],
B_[10][0][189],
B_[10][1][189],
B_[10][2][189],
B_[11][0][189],
B_[11][1][189],
B_[11][2][189],
B_[12][0][189],
B_[12][1][189],
B_[12][2][189],
B_[13][0][189],
B_[13][1][189],
B_[13][2][189],
B_[14][0][189],
B_[14][1][189],
B_[14][2][189],
B_[15][0][189],
B_[15][1][189],
B_[15][2][189],
B_[0][0][190],
B_[0][1][190],
B_[0][2][190],
B_[1][0][190],
B_[1][1][190],
B_[1][2][190],
B_[2][0][190],
B_[2][1][190],
B_[2][2][190],
B_[3][0][190],
B_[3][1][190],
B_[3][2][190],
B_[4][0][190],
B_[4][1][190],
B_[4][2][190],
B_[5][0][190],
B_[5][1][190],
B_[5][2][190],
B_[6][0][190],
B_[6][1][190],
B_[6][2][190],
B_[7][0][190],
B_[7][1][190],
B_[7][2][190],
B_[8][0][190],
B_[8][1][190],
B_[8][2][190],
B_[9][0][190],
B_[9][1][190],
B_[9][2][190],
B_[10][0][190],
B_[10][1][190],
B_[10][2][190],
B_[11][0][190],
B_[11][1][190],
B_[11][2][190],
B_[12][0][190],
B_[12][1][190],
B_[12][2][190],
B_[13][0][190],
B_[13][1][190],
B_[13][2][190],
B_[14][0][190],
B_[14][1][190],
B_[14][2][190],
B_[15][0][190],
B_[15][1][190],
B_[15][2][190],
B_[0][0][191],
B_[0][1][191],
B_[0][2][191],
B_[1][0][191],
B_[1][1][191],
B_[1][2][191],
B_[2][0][191],
B_[2][1][191],
B_[2][2][191],
B_[3][0][191],
B_[3][1][191],
B_[3][2][191],
B_[4][0][191],
B_[4][1][191],
B_[4][2][191],
B_[5][0][191],
B_[5][1][191],
B_[5][2][191],
B_[6][0][191],
B_[6][1][191],
B_[6][2][191],
B_[7][0][191],
B_[7][1][191],
B_[7][2][191],
B_[8][0][191],
B_[8][1][191],
B_[8][2][191],
B_[9][0][191],
B_[9][1][191],
B_[9][2][191],
B_[10][0][191],
B_[10][1][191],
B_[10][2][191],
B_[11][0][191],
B_[11][1][191],
B_[11][2][191],
B_[12][0][191],
B_[12][1][191],
B_[12][2][191],
B_[13][0][191],
B_[13][1][191],
B_[13][2][191],
B_[14][0][191],
B_[14][1][191],
B_[14][2][191],
B_[15][0][191],
B_[15][1][191],
B_[15][2][191],
B_[0][0][192],
B_[0][1][192],
B_[0][2][192],
B_[1][0][192],
B_[1][1][192],
B_[1][2][192],
B_[2][0][192],
B_[2][1][192],
B_[2][2][192],
B_[3][0][192],
B_[3][1][192],
B_[3][2][192],
B_[4][0][192],
B_[4][1][192],
B_[4][2][192],
B_[5][0][192],
B_[5][1][192],
B_[5][2][192],
B_[6][0][192],
B_[6][1][192],
B_[6][2][192],
B_[7][0][192],
B_[7][1][192],
B_[7][2][192],
B_[8][0][192],
B_[8][1][192],
B_[8][2][192],
B_[9][0][192],
B_[9][1][192],
B_[9][2][192],
B_[10][0][192],
B_[10][1][192],
B_[10][2][192],
B_[11][0][192],
B_[11][1][192],
B_[11][2][192],
B_[12][0][192],
B_[12][1][192],
B_[12][2][192],
B_[13][0][192],
B_[13][1][192],
B_[13][2][192],
B_[14][0][192],
B_[14][1][192],
B_[14][2][192],
B_[15][0][192],
B_[15][1][192],
B_[15][2][192],
B_[0][0][193],
B_[0][1][193],
B_[0][2][193],
B_[1][0][193],
B_[1][1][193],
B_[1][2][193],
B_[2][0][193],
B_[2][1][193],
B_[2][2][193],
B_[3][0][193],
B_[3][1][193],
B_[3][2][193],
B_[4][0][193],
B_[4][1][193],
B_[4][2][193],
B_[5][0][193],
B_[5][1][193],
B_[5][2][193],
B_[6][0][193],
B_[6][1][193],
B_[6][2][193],
B_[7][0][193],
B_[7][1][193],
B_[7][2][193],
B_[8][0][193],
B_[8][1][193],
B_[8][2][193],
B_[9][0][193],
B_[9][1][193],
B_[9][2][193],
B_[10][0][193],
B_[10][1][193],
B_[10][2][193],
B_[11][0][193],
B_[11][1][193],
B_[11][2][193],
B_[12][0][193],
B_[12][1][193],
B_[12][2][193],
B_[13][0][193],
B_[13][1][193],
B_[13][2][193],
B_[14][0][193],
B_[14][1][193],
B_[14][2][193],
B_[15][0][193],
B_[15][1][193],
B_[15][2][193],
B_[0][0][194],
B_[0][1][194],
B_[0][2][194],
B_[1][0][194],
B_[1][1][194],
B_[1][2][194],
B_[2][0][194],
B_[2][1][194],
B_[2][2][194],
B_[3][0][194],
B_[3][1][194],
B_[3][2][194],
B_[4][0][194],
B_[4][1][194],
B_[4][2][194],
B_[5][0][194],
B_[5][1][194],
B_[5][2][194],
B_[6][0][194],
B_[6][1][194],
B_[6][2][194],
B_[7][0][194],
B_[7][1][194],
B_[7][2][194],
B_[8][0][194],
B_[8][1][194],
B_[8][2][194],
B_[9][0][194],
B_[9][1][194],
B_[9][2][194],
B_[10][0][194],
B_[10][1][194],
B_[10][2][194],
B_[11][0][194],
B_[11][1][194],
B_[11][2][194],
B_[12][0][194],
B_[12][1][194],
B_[12][2][194],
B_[13][0][194],
B_[13][1][194],
B_[13][2][194],
B_[14][0][194],
B_[14][1][194],
B_[14][2][194],
B_[15][0][194],
B_[15][1][194],
B_[15][2][194],
B_[0][0][195],
B_[0][1][195],
B_[0][2][195],
B_[1][0][195],
B_[1][1][195],
B_[1][2][195],
B_[2][0][195],
B_[2][1][195],
B_[2][2][195],
B_[3][0][195],
B_[3][1][195],
B_[3][2][195],
B_[4][0][195],
B_[4][1][195],
B_[4][2][195],
B_[5][0][195],
B_[5][1][195],
B_[5][2][195],
B_[6][0][195],
B_[6][1][195],
B_[6][2][195],
B_[7][0][195],
B_[7][1][195],
B_[7][2][195],
B_[8][0][195],
B_[8][1][195],
B_[8][2][195],
B_[9][0][195],
B_[9][1][195],
B_[9][2][195],
B_[10][0][195],
B_[10][1][195],
B_[10][2][195],
B_[11][0][195],
B_[11][1][195],
B_[11][2][195],
B_[12][0][195],
B_[12][1][195],
B_[12][2][195],
B_[13][0][195],
B_[13][1][195],
B_[13][2][195],
B_[14][0][195],
B_[14][1][195],
B_[14][2][195],
B_[15][0][195],
B_[15][1][195],
B_[15][2][195],
B_[0][0][196],
B_[0][1][196],
B_[0][2][196],
B_[1][0][196],
B_[1][1][196],
B_[1][2][196],
B_[2][0][196],
B_[2][1][196],
B_[2][2][196],
B_[3][0][196],
B_[3][1][196],
B_[3][2][196],
B_[4][0][196],
B_[4][1][196],
B_[4][2][196],
B_[5][0][196],
B_[5][1][196],
B_[5][2][196],
B_[6][0][196],
B_[6][1][196],
B_[6][2][196],
B_[7][0][196],
B_[7][1][196],
B_[7][2][196],
B_[8][0][196],
B_[8][1][196],
B_[8][2][196],
B_[9][0][196],
B_[9][1][196],
B_[9][2][196],
B_[10][0][196],
B_[10][1][196],
B_[10][2][196],
B_[11][0][196],
B_[11][1][196],
B_[11][2][196],
B_[12][0][196],
B_[12][1][196],
B_[12][2][196],
B_[13][0][196],
B_[13][1][196],
B_[13][2][196],
B_[14][0][196],
B_[14][1][196],
B_[14][2][196],
B_[15][0][196],
B_[15][1][196],
B_[15][2][196],
B_[0][0][197],
B_[0][1][197],
B_[0][2][197],
B_[1][0][197],
B_[1][1][197],
B_[1][2][197],
B_[2][0][197],
B_[2][1][197],
B_[2][2][197],
B_[3][0][197],
B_[3][1][197],
B_[3][2][197],
B_[4][0][197],
B_[4][1][197],
B_[4][2][197],
B_[5][0][197],
B_[5][1][197],
B_[5][2][197],
B_[6][0][197],
B_[6][1][197],
B_[6][2][197],
B_[7][0][197],
B_[7][1][197],
B_[7][2][197],
B_[8][0][197],
B_[8][1][197],
B_[8][2][197],
B_[9][0][197],
B_[9][1][197],
B_[9][2][197],
B_[10][0][197],
B_[10][1][197],
B_[10][2][197],
B_[11][0][197],
B_[11][1][197],
B_[11][2][197],
B_[12][0][197],
B_[12][1][197],
B_[12][2][197],
B_[13][0][197],
B_[13][1][197],
B_[13][2][197],
B_[14][0][197],
B_[14][1][197],
B_[14][2][197],
B_[15][0][197],
B_[15][1][197],
B_[15][2][197],
B_[0][0][198],
B_[0][1][198],
B_[0][2][198],
B_[1][0][198],
B_[1][1][198],
B_[1][2][198],
B_[2][0][198],
B_[2][1][198],
B_[2][2][198],
B_[3][0][198],
B_[3][1][198],
B_[3][2][198],
B_[4][0][198],
B_[4][1][198],
B_[4][2][198],
B_[5][0][198],
B_[5][1][198],
B_[5][2][198],
B_[6][0][198],
B_[6][1][198],
B_[6][2][198],
B_[7][0][198],
B_[7][1][198],
B_[7][2][198],
B_[8][0][198],
B_[8][1][198],
B_[8][2][198],
B_[9][0][198],
B_[9][1][198],
B_[9][2][198],
B_[10][0][198],
B_[10][1][198],
B_[10][2][198],
B_[11][0][198],
B_[11][1][198],
B_[11][2][198],
B_[12][0][198],
B_[12][1][198],
B_[12][2][198],
B_[13][0][198],
B_[13][1][198],
B_[13][2][198],
B_[14][0][198],
B_[14][1][198],
B_[14][2][198],
B_[15][0][198],
B_[15][1][198],
B_[15][2][198],
B_[0][0][199],
B_[0][1][199],
B_[0][2][199],
B_[1][0][199],
B_[1][1][199],
B_[1][2][199],
B_[2][0][199],
B_[2][1][199],
B_[2][2][199],
B_[3][0][199],
B_[3][1][199],
B_[3][2][199],
B_[4][0][199],
B_[4][1][199],
B_[4][2][199],
B_[5][0][199],
B_[5][1][199],
B_[5][2][199],
B_[6][0][199],
B_[6][1][199],
B_[6][2][199],
B_[7][0][199],
B_[7][1][199],
B_[7][2][199],
B_[8][0][199],
B_[8][1][199],
B_[8][2][199],
B_[9][0][199],
B_[9][1][199],
B_[9][2][199],
B_[10][0][199],
B_[10][1][199],
B_[10][2][199],
B_[11][0][199],
B_[11][1][199],
B_[11][2][199],
B_[12][0][199],
B_[12][1][199],
B_[12][2][199],
B_[13][0][199],
B_[13][1][199],
B_[13][2][199],
B_[14][0][199],
B_[14][1][199],
B_[14][2][199],
B_[15][0][199],
B_[15][1][199],
B_[15][2][199],
B_[0][0][200],
B_[0][1][200],
B_[0][2][200],
B_[1][0][200],
B_[1][1][200],
B_[1][2][200],
B_[2][0][200],
B_[2][1][200],
B_[2][2][200],
B_[3][0][200],
B_[3][1][200],
B_[3][2][200],
B_[4][0][200],
B_[4][1][200],
B_[4][2][200],
B_[5][0][200],
B_[5][1][200],
B_[5][2][200],
B_[6][0][200],
B_[6][1][200],
B_[6][2][200],
B_[7][0][200],
B_[7][1][200],
B_[7][2][200],
B_[8][0][200],
B_[8][1][200],
B_[8][2][200],
B_[9][0][200],
B_[9][1][200],
B_[9][2][200],
B_[10][0][200],
B_[10][1][200],
B_[10][2][200],
B_[11][0][200],
B_[11][1][200],
B_[11][2][200],
B_[12][0][200],
B_[12][1][200],
B_[12][2][200],
B_[13][0][200],
B_[13][1][200],
B_[13][2][200],
B_[14][0][200],
B_[14][1][200],
B_[14][2][200],
B_[15][0][200],
B_[15][1][200],
B_[15][2][200],
B_[0][0][201],
B_[0][1][201],
B_[0][2][201],
B_[1][0][201],
B_[1][1][201],
B_[1][2][201],
B_[2][0][201],
B_[2][1][201],
B_[2][2][201],
B_[3][0][201],
B_[3][1][201],
B_[3][2][201],
B_[4][0][201],
B_[4][1][201],
B_[4][2][201],
B_[5][0][201],
B_[5][1][201],
B_[5][2][201],
B_[6][0][201],
B_[6][1][201],
B_[6][2][201],
B_[7][0][201],
B_[7][1][201],
B_[7][2][201],
B_[8][0][201],
B_[8][1][201],
B_[8][2][201],
B_[9][0][201],
B_[9][1][201],
B_[9][2][201],
B_[10][0][201],
B_[10][1][201],
B_[10][2][201],
B_[11][0][201],
B_[11][1][201],
B_[11][2][201],
B_[12][0][201],
B_[12][1][201],
B_[12][2][201],
B_[13][0][201],
B_[13][1][201],
B_[13][2][201],
B_[14][0][201],
B_[14][1][201],
B_[14][2][201],
B_[15][0][201],
B_[15][1][201],
B_[15][2][201],
B_[0][0][202],
B_[0][1][202],
B_[0][2][202],
B_[1][0][202],
B_[1][1][202],
B_[1][2][202],
B_[2][0][202],
B_[2][1][202],
B_[2][2][202],
B_[3][0][202],
B_[3][1][202],
B_[3][2][202],
B_[4][0][202],
B_[4][1][202],
B_[4][2][202],
B_[5][0][202],
B_[5][1][202],
B_[5][2][202],
B_[6][0][202],
B_[6][1][202],
B_[6][2][202],
B_[7][0][202],
B_[7][1][202],
B_[7][2][202],
B_[8][0][202],
B_[8][1][202],
B_[8][2][202],
B_[9][0][202],
B_[9][1][202],
B_[9][2][202],
B_[10][0][202],
B_[10][1][202],
B_[10][2][202],
B_[11][0][202],
B_[11][1][202],
B_[11][2][202],
B_[12][0][202],
B_[12][1][202],
B_[12][2][202],
B_[13][0][202],
B_[13][1][202],
B_[13][2][202],
B_[14][0][202],
B_[14][1][202],
B_[14][2][202],
B_[15][0][202],
B_[15][1][202],
B_[15][2][202],
B_[0][0][203],
B_[0][1][203],
B_[0][2][203],
B_[1][0][203],
B_[1][1][203],
B_[1][2][203],
B_[2][0][203],
B_[2][1][203],
B_[2][2][203],
B_[3][0][203],
B_[3][1][203],
B_[3][2][203],
B_[4][0][203],
B_[4][1][203],
B_[4][2][203],
B_[5][0][203],
B_[5][1][203],
B_[5][2][203],
B_[6][0][203],
B_[6][1][203],
B_[6][2][203],
B_[7][0][203],
B_[7][1][203],
B_[7][2][203],
B_[8][0][203],
B_[8][1][203],
B_[8][2][203],
B_[9][0][203],
B_[9][1][203],
B_[9][2][203],
B_[10][0][203],
B_[10][1][203],
B_[10][2][203],
B_[11][0][203],
B_[11][1][203],
B_[11][2][203],
B_[12][0][203],
B_[12][1][203],
B_[12][2][203],
B_[13][0][203],
B_[13][1][203],
B_[13][2][203],
B_[14][0][203],
B_[14][1][203],
B_[14][2][203],
B_[15][0][203],
B_[15][1][203],
B_[15][2][203],
B_[0][0][204],
B_[0][1][204],
B_[0][2][204],
B_[1][0][204],
B_[1][1][204],
B_[1][2][204],
B_[2][0][204],
B_[2][1][204],
B_[2][2][204],
B_[3][0][204],
B_[3][1][204],
B_[3][2][204],
B_[4][0][204],
B_[4][1][204],
B_[4][2][204],
B_[5][0][204],
B_[5][1][204],
B_[5][2][204],
B_[6][0][204],
B_[6][1][204],
B_[6][2][204],
B_[7][0][204],
B_[7][1][204],
B_[7][2][204],
B_[8][0][204],
B_[8][1][204],
B_[8][2][204],
B_[9][0][204],
B_[9][1][204],
B_[9][2][204],
B_[10][0][204],
B_[10][1][204],
B_[10][2][204],
B_[11][0][204],
B_[11][1][204],
B_[11][2][204],
B_[12][0][204],
B_[12][1][204],
B_[12][2][204],
B_[13][0][204],
B_[13][1][204],
B_[13][2][204],
B_[14][0][204],
B_[14][1][204],
B_[14][2][204],
B_[15][0][204],
B_[15][1][204],
B_[15][2][204],
B_[0][0][205],
B_[0][1][205],
B_[0][2][205],
B_[1][0][205],
B_[1][1][205],
B_[1][2][205],
B_[2][0][205],
B_[2][1][205],
B_[2][2][205],
B_[3][0][205],
B_[3][1][205],
B_[3][2][205],
B_[4][0][205],
B_[4][1][205],
B_[4][2][205],
B_[5][0][205],
B_[5][1][205],
B_[5][2][205],
B_[6][0][205],
B_[6][1][205],
B_[6][2][205],
B_[7][0][205],
B_[7][1][205],
B_[7][2][205],
B_[8][0][205],
B_[8][1][205],
B_[8][2][205],
B_[9][0][205],
B_[9][1][205],
B_[9][2][205],
B_[10][0][205],
B_[10][1][205],
B_[10][2][205],
B_[11][0][205],
B_[11][1][205],
B_[11][2][205],
B_[12][0][205],
B_[12][1][205],
B_[12][2][205],
B_[13][0][205],
B_[13][1][205],
B_[13][2][205],
B_[14][0][205],
B_[14][1][205],
B_[14][2][205],
B_[15][0][205],
B_[15][1][205],
B_[15][2][205],
B_[0][0][206],
B_[0][1][206],
B_[0][2][206],
B_[1][0][206],
B_[1][1][206],
B_[1][2][206],
B_[2][0][206],
B_[2][1][206],
B_[2][2][206],
B_[3][0][206],
B_[3][1][206],
B_[3][2][206],
B_[4][0][206],
B_[4][1][206],
B_[4][2][206],
B_[5][0][206],
B_[5][1][206],
B_[5][2][206],
B_[6][0][206],
B_[6][1][206],
B_[6][2][206],
B_[7][0][206],
B_[7][1][206],
B_[7][2][206],
B_[8][0][206],
B_[8][1][206],
B_[8][2][206],
B_[9][0][206],
B_[9][1][206],
B_[9][2][206],
B_[10][0][206],
B_[10][1][206],
B_[10][2][206],
B_[11][0][206],
B_[11][1][206],
B_[11][2][206],
B_[12][0][206],
B_[12][1][206],
B_[12][2][206],
B_[13][0][206],
B_[13][1][206],
B_[13][2][206],
B_[14][0][206],
B_[14][1][206],
B_[14][2][206],
B_[15][0][206],
B_[15][1][206],
B_[15][2][206],
B_[0][0][207],
B_[0][1][207],
B_[0][2][207],
B_[1][0][207],
B_[1][1][207],
B_[1][2][207],
B_[2][0][207],
B_[2][1][207],
B_[2][2][207],
B_[3][0][207],
B_[3][1][207],
B_[3][2][207],
B_[4][0][207],
B_[4][1][207],
B_[4][2][207],
B_[5][0][207],
B_[5][1][207],
B_[5][2][207],
B_[6][0][207],
B_[6][1][207],
B_[6][2][207],
B_[7][0][207],
B_[7][1][207],
B_[7][2][207],
B_[8][0][207],
B_[8][1][207],
B_[8][2][207],
B_[9][0][207],
B_[9][1][207],
B_[9][2][207],
B_[10][0][207],
B_[10][1][207],
B_[10][2][207],
B_[11][0][207],
B_[11][1][207],
B_[11][2][207],
B_[12][0][207],
B_[12][1][207],
B_[12][2][207],
B_[13][0][207],
B_[13][1][207],
B_[13][2][207],
B_[14][0][207],
B_[14][1][207],
B_[14][2][207],
B_[15][0][207],
B_[15][1][207],
B_[15][2][207],
B_[0][0][208],
B_[0][1][208],
B_[0][2][208],
B_[1][0][208],
B_[1][1][208],
B_[1][2][208],
B_[2][0][208],
B_[2][1][208],
B_[2][2][208],
B_[3][0][208],
B_[3][1][208],
B_[3][2][208],
B_[4][0][208],
B_[4][1][208],
B_[4][2][208],
B_[5][0][208],
B_[5][1][208],
B_[5][2][208],
B_[6][0][208],
B_[6][1][208],
B_[6][2][208],
B_[7][0][208],
B_[7][1][208],
B_[7][2][208],
B_[8][0][208],
B_[8][1][208],
B_[8][2][208],
B_[9][0][208],
B_[9][1][208],
B_[9][2][208],
B_[10][0][208],
B_[10][1][208],
B_[10][2][208],
B_[11][0][208],
B_[11][1][208],
B_[11][2][208],
B_[12][0][208],
B_[12][1][208],
B_[12][2][208],
B_[13][0][208],
B_[13][1][208],
B_[13][2][208],
B_[14][0][208],
B_[14][1][208],
B_[14][2][208],
B_[15][0][208],
B_[15][1][208],
B_[15][2][208],
B_[0][0][209],
B_[0][1][209],
B_[0][2][209],
B_[1][0][209],
B_[1][1][209],
B_[1][2][209],
B_[2][0][209],
B_[2][1][209],
B_[2][2][209],
B_[3][0][209],
B_[3][1][209],
B_[3][2][209],
B_[4][0][209],
B_[4][1][209],
B_[4][2][209],
B_[5][0][209],
B_[5][1][209],
B_[5][2][209],
B_[6][0][209],
B_[6][1][209],
B_[6][2][209],
B_[7][0][209],
B_[7][1][209],
B_[7][2][209],
B_[8][0][209],
B_[8][1][209],
B_[8][2][209],
B_[9][0][209],
B_[9][1][209],
B_[9][2][209],
B_[10][0][209],
B_[10][1][209],
B_[10][2][209],
B_[11][0][209],
B_[11][1][209],
B_[11][2][209],
B_[12][0][209],
B_[12][1][209],
B_[12][2][209],
B_[13][0][209],
B_[13][1][209],
B_[13][2][209],
B_[14][0][209],
B_[14][1][209],
B_[14][2][209],
B_[15][0][209],
B_[15][1][209],
B_[15][2][209],
B_[0][0][210],
B_[0][1][210],
B_[0][2][210],
B_[1][0][210],
B_[1][1][210],
B_[1][2][210],
B_[2][0][210],
B_[2][1][210],
B_[2][2][210],
B_[3][0][210],
B_[3][1][210],
B_[3][2][210],
B_[4][0][210],
B_[4][1][210],
B_[4][2][210],
B_[5][0][210],
B_[5][1][210],
B_[5][2][210],
B_[6][0][210],
B_[6][1][210],
B_[6][2][210],
B_[7][0][210],
B_[7][1][210],
B_[7][2][210],
B_[8][0][210],
B_[8][1][210],
B_[8][2][210],
B_[9][0][210],
B_[9][1][210],
B_[9][2][210],
B_[10][0][210],
B_[10][1][210],
B_[10][2][210],
B_[11][0][210],
B_[11][1][210],
B_[11][2][210],
B_[12][0][210],
B_[12][1][210],
B_[12][2][210],
B_[13][0][210],
B_[13][1][210],
B_[13][2][210],
B_[14][0][210],
B_[14][1][210],
B_[14][2][210],
B_[15][0][210],
B_[15][1][210],
B_[15][2][210],
B_[0][0][211],
B_[0][1][211],
B_[0][2][211],
B_[1][0][211],
B_[1][1][211],
B_[1][2][211],
B_[2][0][211],
B_[2][1][211],
B_[2][2][211],
B_[3][0][211],
B_[3][1][211],
B_[3][2][211],
B_[4][0][211],
B_[4][1][211],
B_[4][2][211],
B_[5][0][211],
B_[5][1][211],
B_[5][2][211],
B_[6][0][211],
B_[6][1][211],
B_[6][2][211],
B_[7][0][211],
B_[7][1][211],
B_[7][2][211],
B_[8][0][211],
B_[8][1][211],
B_[8][2][211],
B_[9][0][211],
B_[9][1][211],
B_[9][2][211],
B_[10][0][211],
B_[10][1][211],
B_[10][2][211],
B_[11][0][211],
B_[11][1][211],
B_[11][2][211],
B_[12][0][211],
B_[12][1][211],
B_[12][2][211],
B_[13][0][211],
B_[13][1][211],
B_[13][2][211],
B_[14][0][211],
B_[14][1][211],
B_[14][2][211],
B_[15][0][211],
B_[15][1][211],
B_[15][2][211],
B_[0][0][212],
B_[0][1][212],
B_[0][2][212],
B_[1][0][212],
B_[1][1][212],
B_[1][2][212],
B_[2][0][212],
B_[2][1][212],
B_[2][2][212],
B_[3][0][212],
B_[3][1][212],
B_[3][2][212],
B_[4][0][212],
B_[4][1][212],
B_[4][2][212],
B_[5][0][212],
B_[5][1][212],
B_[5][2][212],
B_[6][0][212],
B_[6][1][212],
B_[6][2][212],
B_[7][0][212],
B_[7][1][212],
B_[7][2][212],
B_[8][0][212],
B_[8][1][212],
B_[8][2][212],
B_[9][0][212],
B_[9][1][212],
B_[9][2][212],
B_[10][0][212],
B_[10][1][212],
B_[10][2][212],
B_[11][0][212],
B_[11][1][212],
B_[11][2][212],
B_[12][0][212],
B_[12][1][212],
B_[12][2][212],
B_[13][0][212],
B_[13][1][212],
B_[13][2][212],
B_[14][0][212],
B_[14][1][212],
B_[14][2][212],
B_[15][0][212],
B_[15][1][212],
B_[15][2][212],
B_[0][0][213],
B_[0][1][213],
B_[0][2][213],
B_[1][0][213],
B_[1][1][213],
B_[1][2][213],
B_[2][0][213],
B_[2][1][213],
B_[2][2][213],
B_[3][0][213],
B_[3][1][213],
B_[3][2][213],
B_[4][0][213],
B_[4][1][213],
B_[4][2][213],
B_[5][0][213],
B_[5][1][213],
B_[5][2][213],
B_[6][0][213],
B_[6][1][213],
B_[6][2][213],
B_[7][0][213],
B_[7][1][213],
B_[7][2][213],
B_[8][0][213],
B_[8][1][213],
B_[8][2][213],
B_[9][0][213],
B_[9][1][213],
B_[9][2][213],
B_[10][0][213],
B_[10][1][213],
B_[10][2][213],
B_[11][0][213],
B_[11][1][213],
B_[11][2][213],
B_[12][0][213],
B_[12][1][213],
B_[12][2][213],
B_[13][0][213],
B_[13][1][213],
B_[13][2][213],
B_[14][0][213],
B_[14][1][213],
B_[14][2][213],
B_[15][0][213],
B_[15][1][213],
B_[15][2][213],
B_[0][0][214],
B_[0][1][214],
B_[0][2][214],
B_[1][0][214],
B_[1][1][214],
B_[1][2][214],
B_[2][0][214],
B_[2][1][214],
B_[2][2][214],
B_[3][0][214],
B_[3][1][214],
B_[3][2][214],
B_[4][0][214],
B_[4][1][214],
B_[4][2][214],
B_[5][0][214],
B_[5][1][214],
B_[5][2][214],
B_[6][0][214],
B_[6][1][214],
B_[6][2][214],
B_[7][0][214],
B_[7][1][214],
B_[7][2][214],
B_[8][0][214],
B_[8][1][214],
B_[8][2][214],
B_[9][0][214],
B_[9][1][214],
B_[9][2][214],
B_[10][0][214],
B_[10][1][214],
B_[10][2][214],
B_[11][0][214],
B_[11][1][214],
B_[11][2][214],
B_[12][0][214],
B_[12][1][214],
B_[12][2][214],
B_[13][0][214],
B_[13][1][214],
B_[13][2][214],
B_[14][0][214],
B_[14][1][214],
B_[14][2][214],
B_[15][0][214],
B_[15][1][214],
B_[15][2][214],
B_[0][0][215],
B_[0][1][215],
B_[0][2][215],
B_[1][0][215],
B_[1][1][215],
B_[1][2][215],
B_[2][0][215],
B_[2][1][215],
B_[2][2][215],
B_[3][0][215],
B_[3][1][215],
B_[3][2][215],
B_[4][0][215],
B_[4][1][215],
B_[4][2][215],
B_[5][0][215],
B_[5][1][215],
B_[5][2][215],
B_[6][0][215],
B_[6][1][215],
B_[6][2][215],
B_[7][0][215],
B_[7][1][215],
B_[7][2][215],
B_[8][0][215],
B_[8][1][215],
B_[8][2][215],
B_[9][0][215],
B_[9][1][215],
B_[9][2][215],
B_[10][0][215],
B_[10][1][215],
B_[10][2][215],
B_[11][0][215],
B_[11][1][215],
B_[11][2][215],
B_[12][0][215],
B_[12][1][215],
B_[12][2][215],
B_[13][0][215],
B_[13][1][215],
B_[13][2][215],
B_[14][0][215],
B_[14][1][215],
B_[14][2][215],
B_[15][0][215],
B_[15][1][215],
B_[15][2][215],
B_[0][0][216],
B_[0][1][216],
B_[0][2][216],
B_[1][0][216],
B_[1][1][216],
B_[1][2][216],
B_[2][0][216],
B_[2][1][216],
B_[2][2][216],
B_[3][0][216],
B_[3][1][216],
B_[3][2][216],
B_[4][0][216],
B_[4][1][216],
B_[4][2][216],
B_[5][0][216],
B_[5][1][216],
B_[5][2][216],
B_[6][0][216],
B_[6][1][216],
B_[6][2][216],
B_[7][0][216],
B_[7][1][216],
B_[7][2][216],
B_[8][0][216],
B_[8][1][216],
B_[8][2][216],
B_[9][0][216],
B_[9][1][216],
B_[9][2][216],
B_[10][0][216],
B_[10][1][216],
B_[10][2][216],
B_[11][0][216],
B_[11][1][216],
B_[11][2][216],
B_[12][0][216],
B_[12][1][216],
B_[12][2][216],
B_[13][0][216],
B_[13][1][216],
B_[13][2][216],
B_[14][0][216],
B_[14][1][216],
B_[14][2][216],
B_[15][0][216],
B_[15][1][216],
B_[15][2][216],
B_[0][0][217],
B_[0][1][217],
B_[0][2][217],
B_[1][0][217],
B_[1][1][217],
B_[1][2][217],
B_[2][0][217],
B_[2][1][217],
B_[2][2][217],
B_[3][0][217],
B_[3][1][217],
B_[3][2][217],
B_[4][0][217],
B_[4][1][217],
B_[4][2][217],
B_[5][0][217],
B_[5][1][217],
B_[5][2][217],
B_[6][0][217],
B_[6][1][217],
B_[6][2][217],
B_[7][0][217],
B_[7][1][217],
B_[7][2][217],
B_[8][0][217],
B_[8][1][217],
B_[8][2][217],
B_[9][0][217],
B_[9][1][217],
B_[9][2][217],
B_[10][0][217],
B_[10][1][217],
B_[10][2][217],
B_[11][0][217],
B_[11][1][217],
B_[11][2][217],
B_[12][0][217],
B_[12][1][217],
B_[12][2][217],
B_[13][0][217],
B_[13][1][217],
B_[13][2][217],
B_[14][0][217],
B_[14][1][217],
B_[14][2][217],
B_[15][0][217],
B_[15][1][217],
B_[15][2][217],
B_[0][0][218],
B_[0][1][218],
B_[0][2][218],
B_[1][0][218],
B_[1][1][218],
B_[1][2][218],
B_[2][0][218],
B_[2][1][218],
B_[2][2][218],
B_[3][0][218],
B_[3][1][218],
B_[3][2][218],
B_[4][0][218],
B_[4][1][218],
B_[4][2][218],
B_[5][0][218],
B_[5][1][218],
B_[5][2][218],
B_[6][0][218],
B_[6][1][218],
B_[6][2][218],
B_[7][0][218],
B_[7][1][218],
B_[7][2][218],
B_[8][0][218],
B_[8][1][218],
B_[8][2][218],
B_[9][0][218],
B_[9][1][218],
B_[9][2][218],
B_[10][0][218],
B_[10][1][218],
B_[10][2][218],
B_[11][0][218],
B_[11][1][218],
B_[11][2][218],
B_[12][0][218],
B_[12][1][218],
B_[12][2][218],
B_[13][0][218],
B_[13][1][218],
B_[13][2][218],
B_[14][0][218],
B_[14][1][218],
B_[14][2][218],
B_[15][0][218],
B_[15][1][218],
B_[15][2][218],
B_[0][0][219],
B_[0][1][219],
B_[0][2][219],
B_[1][0][219],
B_[1][1][219],
B_[1][2][219],
B_[2][0][219],
B_[2][1][219],
B_[2][2][219],
B_[3][0][219],
B_[3][1][219],
B_[3][2][219],
B_[4][0][219],
B_[4][1][219],
B_[4][2][219],
B_[5][0][219],
B_[5][1][219],
B_[5][2][219],
B_[6][0][219],
B_[6][1][219],
B_[6][2][219],
B_[7][0][219],
B_[7][1][219],
B_[7][2][219],
B_[8][0][219],
B_[8][1][219],
B_[8][2][219],
B_[9][0][219],
B_[9][1][219],
B_[9][2][219],
B_[10][0][219],
B_[10][1][219],
B_[10][2][219],
B_[11][0][219],
B_[11][1][219],
B_[11][2][219],
B_[12][0][219],
B_[12][1][219],
B_[12][2][219],
B_[13][0][219],
B_[13][1][219],
B_[13][2][219],
B_[14][0][219],
B_[14][1][219],
B_[14][2][219],
B_[15][0][219],
B_[15][1][219],
B_[15][2][219],
B_[0][0][220],
B_[0][1][220],
B_[0][2][220],
B_[1][0][220],
B_[1][1][220],
B_[1][2][220],
B_[2][0][220],
B_[2][1][220],
B_[2][2][220],
B_[3][0][220],
B_[3][1][220],
B_[3][2][220],
B_[4][0][220],
B_[4][1][220],
B_[4][2][220],
B_[5][0][220],
B_[5][1][220],
B_[5][2][220],
B_[6][0][220],
B_[6][1][220],
B_[6][2][220],
B_[7][0][220],
B_[7][1][220],
B_[7][2][220],
B_[8][0][220],
B_[8][1][220],
B_[8][2][220],
B_[9][0][220],
B_[9][1][220],
B_[9][2][220],
B_[10][0][220],
B_[10][1][220],
B_[10][2][220],
B_[11][0][220],
B_[11][1][220],
B_[11][2][220],
B_[12][0][220],
B_[12][1][220],
B_[12][2][220],
B_[13][0][220],
B_[13][1][220],
B_[13][2][220],
B_[14][0][220],
B_[14][1][220],
B_[14][2][220],
B_[15][0][220],
B_[15][1][220],
B_[15][2][220],
B_[0][0][221],
B_[0][1][221],
B_[0][2][221],
B_[1][0][221],
B_[1][1][221],
B_[1][2][221],
B_[2][0][221],
B_[2][1][221],
B_[2][2][221],
B_[3][0][221],
B_[3][1][221],
B_[3][2][221],
B_[4][0][221],
B_[4][1][221],
B_[4][2][221],
B_[5][0][221],
B_[5][1][221],
B_[5][2][221],
B_[6][0][221],
B_[6][1][221],
B_[6][2][221],
B_[7][0][221],
B_[7][1][221],
B_[7][2][221],
B_[8][0][221],
B_[8][1][221],
B_[8][2][221],
B_[9][0][221],
B_[9][1][221],
B_[9][2][221],
B_[10][0][221],
B_[10][1][221],
B_[10][2][221],
B_[11][0][221],
B_[11][1][221],
B_[11][2][221],
B_[12][0][221],
B_[12][1][221],
B_[12][2][221],
B_[13][0][221],
B_[13][1][221],
B_[13][2][221],
B_[14][0][221],
B_[14][1][221],
B_[14][2][221],
B_[15][0][221],
B_[15][1][221],
B_[15][2][221],
B_[0][0][222],
B_[0][1][222],
B_[0][2][222],
B_[1][0][222],
B_[1][1][222],
B_[1][2][222],
B_[2][0][222],
B_[2][1][222],
B_[2][2][222],
B_[3][0][222],
B_[3][1][222],
B_[3][2][222],
B_[4][0][222],
B_[4][1][222],
B_[4][2][222],
B_[5][0][222],
B_[5][1][222],
B_[5][2][222],
B_[6][0][222],
B_[6][1][222],
B_[6][2][222],
B_[7][0][222],
B_[7][1][222],
B_[7][2][222],
B_[8][0][222],
B_[8][1][222],
B_[8][2][222],
B_[9][0][222],
B_[9][1][222],
B_[9][2][222],
B_[10][0][222],
B_[10][1][222],
B_[10][2][222],
B_[11][0][222],
B_[11][1][222],
B_[11][2][222],
B_[12][0][222],
B_[12][1][222],
B_[12][2][222],
B_[13][0][222],
B_[13][1][222],
B_[13][2][222],
B_[14][0][222],
B_[14][1][222],
B_[14][2][222],
B_[15][0][222],
B_[15][1][222],
B_[15][2][222],
B_[0][0][223],
B_[0][1][223],
B_[0][2][223],
B_[1][0][223],
B_[1][1][223],
B_[1][2][223],
B_[2][0][223],
B_[2][1][223],
B_[2][2][223],
B_[3][0][223],
B_[3][1][223],
B_[3][2][223],
B_[4][0][223],
B_[4][1][223],
B_[4][2][223],
B_[5][0][223],
B_[5][1][223],
B_[5][2][223],
B_[6][0][223],
B_[6][1][223],
B_[6][2][223],
B_[7][0][223],
B_[7][1][223],
B_[7][2][223],
B_[8][0][223],
B_[8][1][223],
B_[8][2][223],
B_[9][0][223],
B_[9][1][223],
B_[9][2][223],
B_[10][0][223],
B_[10][1][223],
B_[10][2][223],
B_[11][0][223],
B_[11][1][223],
B_[11][2][223],
B_[12][0][223],
B_[12][1][223],
B_[12][2][223],
B_[13][0][223],
B_[13][1][223],
B_[13][2][223],
B_[14][0][223],
B_[14][1][223],
B_[14][2][223],
B_[15][0][223],
B_[15][1][223],
B_[15][2][223],
B_[0][0][224],
B_[0][1][224],
B_[0][2][224],
B_[1][0][224],
B_[1][1][224],
B_[1][2][224],
B_[2][0][224],
B_[2][1][224],
B_[2][2][224],
B_[3][0][224],
B_[3][1][224],
B_[3][2][224],
B_[4][0][224],
B_[4][1][224],
B_[4][2][224],
B_[5][0][224],
B_[5][1][224],
B_[5][2][224],
B_[6][0][224],
B_[6][1][224],
B_[6][2][224],
B_[7][0][224],
B_[7][1][224],
B_[7][2][224],
B_[8][0][224],
B_[8][1][224],
B_[8][2][224],
B_[9][0][224],
B_[9][1][224],
B_[9][2][224],
B_[10][0][224],
B_[10][1][224],
B_[10][2][224],
B_[11][0][224],
B_[11][1][224],
B_[11][2][224],
B_[12][0][224],
B_[12][1][224],
B_[12][2][224],
B_[13][0][224],
B_[13][1][224],
B_[13][2][224],
B_[14][0][224],
B_[14][1][224],
B_[14][2][224],
B_[15][0][224],
B_[15][1][224],
B_[15][2][224],
B_[0][0][225],
B_[0][1][225],
B_[0][2][225],
B_[1][0][225],
B_[1][1][225],
B_[1][2][225],
B_[2][0][225],
B_[2][1][225],
B_[2][2][225],
B_[3][0][225],
B_[3][1][225],
B_[3][2][225],
B_[4][0][225],
B_[4][1][225],
B_[4][2][225],
B_[5][0][225],
B_[5][1][225],
B_[5][2][225],
B_[6][0][225],
B_[6][1][225],
B_[6][2][225],
B_[7][0][225],
B_[7][1][225],
B_[7][2][225],
B_[8][0][225],
B_[8][1][225],
B_[8][2][225],
B_[9][0][225],
B_[9][1][225],
B_[9][2][225],
B_[10][0][225],
B_[10][1][225],
B_[10][2][225],
B_[11][0][225],
B_[11][1][225],
B_[11][2][225],
B_[12][0][225],
B_[12][1][225],
B_[12][2][225],
B_[13][0][225],
B_[13][1][225],
B_[13][2][225],
B_[14][0][225],
B_[14][1][225],
B_[14][2][225],
B_[15][0][225],
B_[15][1][225],
B_[15][2][225],
B_[0][0][226],
B_[0][1][226],
B_[0][2][226],
B_[1][0][226],
B_[1][1][226],
B_[1][2][226],
B_[2][0][226],
B_[2][1][226],
B_[2][2][226],
B_[3][0][226],
B_[3][1][226],
B_[3][2][226],
B_[4][0][226],
B_[4][1][226],
B_[4][2][226],
B_[5][0][226],
B_[5][1][226],
B_[5][2][226],
B_[6][0][226],
B_[6][1][226],
B_[6][2][226],
B_[7][0][226],
B_[7][1][226],
B_[7][2][226],
B_[8][0][226],
B_[8][1][226],
B_[8][2][226],
B_[9][0][226],
B_[9][1][226],
B_[9][2][226],
B_[10][0][226],
B_[10][1][226],
B_[10][2][226],
B_[11][0][226],
B_[11][1][226],
B_[11][2][226],
B_[12][0][226],
B_[12][1][226],
B_[12][2][226],
B_[13][0][226],
B_[13][1][226],
B_[13][2][226],
B_[14][0][226],
B_[14][1][226],
B_[14][2][226],
B_[15][0][226],
B_[15][1][226],
B_[15][2][226],
B_[0][0][227],
B_[0][1][227],
B_[0][2][227],
B_[1][0][227],
B_[1][1][227],
B_[1][2][227],
B_[2][0][227],
B_[2][1][227],
B_[2][2][227],
B_[3][0][227],
B_[3][1][227],
B_[3][2][227],
B_[4][0][227],
B_[4][1][227],
B_[4][2][227],
B_[5][0][227],
B_[5][1][227],
B_[5][2][227],
B_[6][0][227],
B_[6][1][227],
B_[6][2][227],
B_[7][0][227],
B_[7][1][227],
B_[7][2][227],
B_[8][0][227],
B_[8][1][227],
B_[8][2][227],
B_[9][0][227],
B_[9][1][227],
B_[9][2][227],
B_[10][0][227],
B_[10][1][227],
B_[10][2][227],
B_[11][0][227],
B_[11][1][227],
B_[11][2][227],
B_[12][0][227],
B_[12][1][227],
B_[12][2][227],
B_[13][0][227],
B_[13][1][227],
B_[13][2][227],
B_[14][0][227],
B_[14][1][227],
B_[14][2][227],
B_[15][0][227],
B_[15][1][227],
B_[15][2][227],
B_[0][0][228],
B_[0][1][228],
B_[0][2][228],
B_[1][0][228],
B_[1][1][228],
B_[1][2][228],
B_[2][0][228],
B_[2][1][228],
B_[2][2][228],
B_[3][0][228],
B_[3][1][228],
B_[3][2][228],
B_[4][0][228],
B_[4][1][228],
B_[4][2][228],
B_[5][0][228],
B_[5][1][228],
B_[5][2][228],
B_[6][0][228],
B_[6][1][228],
B_[6][2][228],
B_[7][0][228],
B_[7][1][228],
B_[7][2][228],
B_[8][0][228],
B_[8][1][228],
B_[8][2][228],
B_[9][0][228],
B_[9][1][228],
B_[9][2][228],
B_[10][0][228],
B_[10][1][228],
B_[10][2][228],
B_[11][0][228],
B_[11][1][228],
B_[11][2][228],
B_[12][0][228],
B_[12][1][228],
B_[12][2][228],
B_[13][0][228],
B_[13][1][228],
B_[13][2][228],
B_[14][0][228],
B_[14][1][228],
B_[14][2][228],
B_[15][0][228],
B_[15][1][228],
B_[15][2][228],
B_[0][0][229],
B_[0][1][229],
B_[0][2][229],
B_[1][0][229],
B_[1][1][229],
B_[1][2][229],
B_[2][0][229],
B_[2][1][229],
B_[2][2][229],
B_[3][0][229],
B_[3][1][229],
B_[3][2][229],
B_[4][0][229],
B_[4][1][229],
B_[4][2][229],
B_[5][0][229],
B_[5][1][229],
B_[5][2][229],
B_[6][0][229],
B_[6][1][229],
B_[6][2][229],
B_[7][0][229],
B_[7][1][229],
B_[7][2][229],
B_[8][0][229],
B_[8][1][229],
B_[8][2][229],
B_[9][0][229],
B_[9][1][229],
B_[9][2][229],
B_[10][0][229],
B_[10][1][229],
B_[10][2][229],
B_[11][0][229],
B_[11][1][229],
B_[11][2][229],
B_[12][0][229],
B_[12][1][229],
B_[12][2][229],
B_[13][0][229],
B_[13][1][229],
B_[13][2][229],
B_[14][0][229],
B_[14][1][229],
B_[14][2][229],
B_[15][0][229],
B_[15][1][229],
B_[15][2][229],
B_[0][0][230],
B_[0][1][230],
B_[0][2][230],
B_[1][0][230],
B_[1][1][230],
B_[1][2][230],
B_[2][0][230],
B_[2][1][230],
B_[2][2][230],
B_[3][0][230],
B_[3][1][230],
B_[3][2][230],
B_[4][0][230],
B_[4][1][230],
B_[4][2][230],
B_[5][0][230],
B_[5][1][230],
B_[5][2][230],
B_[6][0][230],
B_[6][1][230],
B_[6][2][230],
B_[7][0][230],
B_[7][1][230],
B_[7][2][230],
B_[8][0][230],
B_[8][1][230],
B_[8][2][230],
B_[9][0][230],
B_[9][1][230],
B_[9][2][230],
B_[10][0][230],
B_[10][1][230],
B_[10][2][230],
B_[11][0][230],
B_[11][1][230],
B_[11][2][230],
B_[12][0][230],
B_[12][1][230],
B_[12][2][230],
B_[13][0][230],
B_[13][1][230],
B_[13][2][230],
B_[14][0][230],
B_[14][1][230],
B_[14][2][230],
B_[15][0][230],
B_[15][1][230],
B_[15][2][230],
B_[0][0][231],
B_[0][1][231],
B_[0][2][231],
B_[1][0][231],
B_[1][1][231],
B_[1][2][231],
B_[2][0][231],
B_[2][1][231],
B_[2][2][231],
B_[3][0][231],
B_[3][1][231],
B_[3][2][231],
B_[4][0][231],
B_[4][1][231],
B_[4][2][231],
B_[5][0][231],
B_[5][1][231],
B_[5][2][231],
B_[6][0][231],
B_[6][1][231],
B_[6][2][231],
B_[7][0][231],
B_[7][1][231],
B_[7][2][231],
B_[8][0][231],
B_[8][1][231],
B_[8][2][231],
B_[9][0][231],
B_[9][1][231],
B_[9][2][231],
B_[10][0][231],
B_[10][1][231],
B_[10][2][231],
B_[11][0][231],
B_[11][1][231],
B_[11][2][231],
B_[12][0][231],
B_[12][1][231],
B_[12][2][231],
B_[13][0][231],
B_[13][1][231],
B_[13][2][231],
B_[14][0][231],
B_[14][1][231],
B_[14][2][231],
B_[15][0][231],
B_[15][1][231],
B_[15][2][231],
B_[0][0][232],
B_[0][1][232],
B_[0][2][232],
B_[1][0][232],
B_[1][1][232],
B_[1][2][232],
B_[2][0][232],
B_[2][1][232],
B_[2][2][232],
B_[3][0][232],
B_[3][1][232],
B_[3][2][232],
B_[4][0][232],
B_[4][1][232],
B_[4][2][232],
B_[5][0][232],
B_[5][1][232],
B_[5][2][232],
B_[6][0][232],
B_[6][1][232],
B_[6][2][232],
B_[7][0][232],
B_[7][1][232],
B_[7][2][232],
B_[8][0][232],
B_[8][1][232],
B_[8][2][232],
B_[9][0][232],
B_[9][1][232],
B_[9][2][232],
B_[10][0][232],
B_[10][1][232],
B_[10][2][232],
B_[11][0][232],
B_[11][1][232],
B_[11][2][232],
B_[12][0][232],
B_[12][1][232],
B_[12][2][232],
B_[13][0][232],
B_[13][1][232],
B_[13][2][232],
B_[14][0][232],
B_[14][1][232],
B_[14][2][232],
B_[15][0][232],
B_[15][1][232],
B_[15][2][232],
B_[0][0][233],
B_[0][1][233],
B_[0][2][233],
B_[1][0][233],
B_[1][1][233],
B_[1][2][233],
B_[2][0][233],
B_[2][1][233],
B_[2][2][233],
B_[3][0][233],
B_[3][1][233],
B_[3][2][233],
B_[4][0][233],
B_[4][1][233],
B_[4][2][233],
B_[5][0][233],
B_[5][1][233],
B_[5][2][233],
B_[6][0][233],
B_[6][1][233],
B_[6][2][233],
B_[7][0][233],
B_[7][1][233],
B_[7][2][233],
B_[8][0][233],
B_[8][1][233],
B_[8][2][233],
B_[9][0][233],
B_[9][1][233],
B_[9][2][233],
B_[10][0][233],
B_[10][1][233],
B_[10][2][233],
B_[11][0][233],
B_[11][1][233],
B_[11][2][233],
B_[12][0][233],
B_[12][1][233],
B_[12][2][233],
B_[13][0][233],
B_[13][1][233],
B_[13][2][233],
B_[14][0][233],
B_[14][1][233],
B_[14][2][233],
B_[15][0][233],
B_[15][1][233],
B_[15][2][233],
B_[0][0][234],
B_[0][1][234],
B_[0][2][234],
B_[1][0][234],
B_[1][1][234],
B_[1][2][234],
B_[2][0][234],
B_[2][1][234],
B_[2][2][234],
B_[3][0][234],
B_[3][1][234],
B_[3][2][234],
B_[4][0][234],
B_[4][1][234],
B_[4][2][234],
B_[5][0][234],
B_[5][1][234],
B_[5][2][234],
B_[6][0][234],
B_[6][1][234],
B_[6][2][234],
B_[7][0][234],
B_[7][1][234],
B_[7][2][234],
B_[8][0][234],
B_[8][1][234],
B_[8][2][234],
B_[9][0][234],
B_[9][1][234],
B_[9][2][234],
B_[10][0][234],
B_[10][1][234],
B_[10][2][234],
B_[11][0][234],
B_[11][1][234],
B_[11][2][234],
B_[12][0][234],
B_[12][1][234],
B_[12][2][234],
B_[13][0][234],
B_[13][1][234],
B_[13][2][234],
B_[14][0][234],
B_[14][1][234],
B_[14][2][234],
B_[15][0][234],
B_[15][1][234],
B_[15][2][234],
B_[0][0][235],
B_[0][1][235],
B_[0][2][235],
B_[1][0][235],
B_[1][1][235],
B_[1][2][235],
B_[2][0][235],
B_[2][1][235],
B_[2][2][235],
B_[3][0][235],
B_[3][1][235],
B_[3][2][235],
B_[4][0][235],
B_[4][1][235],
B_[4][2][235],
B_[5][0][235],
B_[5][1][235],
B_[5][2][235],
B_[6][0][235],
B_[6][1][235],
B_[6][2][235],
B_[7][0][235],
B_[7][1][235],
B_[7][2][235],
B_[8][0][235],
B_[8][1][235],
B_[8][2][235],
B_[9][0][235],
B_[9][1][235],
B_[9][2][235],
B_[10][0][235],
B_[10][1][235],
B_[10][2][235],
B_[11][0][235],
B_[11][1][235],
B_[11][2][235],
B_[12][0][235],
B_[12][1][235],
B_[12][2][235],
B_[13][0][235],
B_[13][1][235],
B_[13][2][235],
B_[14][0][235],
B_[14][1][235],
B_[14][2][235],
B_[15][0][235],
B_[15][1][235],
B_[15][2][235],
B_[0][0][236],
B_[0][1][236],
B_[0][2][236],
B_[1][0][236],
B_[1][1][236],
B_[1][2][236],
B_[2][0][236],
B_[2][1][236],
B_[2][2][236],
B_[3][0][236],
B_[3][1][236],
B_[3][2][236],
B_[4][0][236],
B_[4][1][236],
B_[4][2][236],
B_[5][0][236],
B_[5][1][236],
B_[5][2][236],
B_[6][0][236],
B_[6][1][236],
B_[6][2][236],
B_[7][0][236],
B_[7][1][236],
B_[7][2][236],
B_[8][0][236],
B_[8][1][236],
B_[8][2][236],
B_[9][0][236],
B_[9][1][236],
B_[9][2][236],
B_[10][0][236],
B_[10][1][236],
B_[10][2][236],
B_[11][0][236],
B_[11][1][236],
B_[11][2][236],
B_[12][0][236],
B_[12][1][236],
B_[12][2][236],
B_[13][0][236],
B_[13][1][236],
B_[13][2][236],
B_[14][0][236],
B_[14][1][236],
B_[14][2][236],
B_[15][0][236],
B_[15][1][236],
B_[15][2][236],
B_[0][0][237],
B_[0][1][237],
B_[0][2][237],
B_[1][0][237],
B_[1][1][237],
B_[1][2][237],
B_[2][0][237],
B_[2][1][237],
B_[2][2][237],
B_[3][0][237],
B_[3][1][237],
B_[3][2][237],
B_[4][0][237],
B_[4][1][237],
B_[4][2][237],
B_[5][0][237],
B_[5][1][237],
B_[5][2][237],
B_[6][0][237],
B_[6][1][237],
B_[6][2][237],
B_[7][0][237],
B_[7][1][237],
B_[7][2][237],
B_[8][0][237],
B_[8][1][237],
B_[8][2][237],
B_[9][0][237],
B_[9][1][237],
B_[9][2][237],
B_[10][0][237],
B_[10][1][237],
B_[10][2][237],
B_[11][0][237],
B_[11][1][237],
B_[11][2][237],
B_[12][0][237],
B_[12][1][237],
B_[12][2][237],
B_[13][0][237],
B_[13][1][237],
B_[13][2][237],
B_[14][0][237],
B_[14][1][237],
B_[14][2][237],
B_[15][0][237],
B_[15][1][237],
B_[15][2][237],
B_[0][0][238],
B_[0][1][238],
B_[0][2][238],
B_[1][0][238],
B_[1][1][238],
B_[1][2][238],
B_[2][0][238],
B_[2][1][238],
B_[2][2][238],
B_[3][0][238],
B_[3][1][238],
B_[3][2][238],
B_[4][0][238],
B_[4][1][238],
B_[4][2][238],
B_[5][0][238],
B_[5][1][238],
B_[5][2][238],
B_[6][0][238],
B_[6][1][238],
B_[6][2][238],
B_[7][0][238],
B_[7][1][238],
B_[7][2][238],
B_[8][0][238],
B_[8][1][238],
B_[8][2][238],
B_[9][0][238],
B_[9][1][238],
B_[9][2][238],
B_[10][0][238],
B_[10][1][238],
B_[10][2][238],
B_[11][0][238],
B_[11][1][238],
B_[11][2][238],
B_[12][0][238],
B_[12][1][238],
B_[12][2][238],
B_[13][0][238],
B_[13][1][238],
B_[13][2][238],
B_[14][0][238],
B_[14][1][238],
B_[14][2][238],
B_[15][0][238],
B_[15][1][238],
B_[15][2][238],
B_[0][0][239],
B_[0][1][239],
B_[0][2][239],
B_[1][0][239],
B_[1][1][239],
B_[1][2][239],
B_[2][0][239],
B_[2][1][239],
B_[2][2][239],
B_[3][0][239],
B_[3][1][239],
B_[3][2][239],
B_[4][0][239],
B_[4][1][239],
B_[4][2][239],
B_[5][0][239],
B_[5][1][239],
B_[5][2][239],
B_[6][0][239],
B_[6][1][239],
B_[6][2][239],
B_[7][0][239],
B_[7][1][239],
B_[7][2][239],
B_[8][0][239],
B_[8][1][239],
B_[8][2][239],
B_[9][0][239],
B_[9][1][239],
B_[9][2][239],
B_[10][0][239],
B_[10][1][239],
B_[10][2][239],
B_[11][0][239],
B_[11][1][239],
B_[11][2][239],
B_[12][0][239],
B_[12][1][239],
B_[12][2][239],
B_[13][0][239],
B_[13][1][239],
B_[13][2][239],
B_[14][0][239],
B_[14][1][239],
B_[14][2][239],
B_[15][0][239],
B_[15][1][239],
B_[15][2][239],
B_[0][0][240],
B_[0][1][240],
B_[0][2][240],
B_[1][0][240],
B_[1][1][240],
B_[1][2][240],
B_[2][0][240],
B_[2][1][240],
B_[2][2][240],
B_[3][0][240],
B_[3][1][240],
B_[3][2][240],
B_[4][0][240],
B_[4][1][240],
B_[4][2][240],
B_[5][0][240],
B_[5][1][240],
B_[5][2][240],
B_[6][0][240],
B_[6][1][240],
B_[6][2][240],
B_[7][0][240],
B_[7][1][240],
B_[7][2][240],
B_[8][0][240],
B_[8][1][240],
B_[8][2][240],
B_[9][0][240],
B_[9][1][240],
B_[9][2][240],
B_[10][0][240],
B_[10][1][240],
B_[10][2][240],
B_[11][0][240],
B_[11][1][240],
B_[11][2][240],
B_[12][0][240],
B_[12][1][240],
B_[12][2][240],
B_[13][0][240],
B_[13][1][240],
B_[13][2][240],
B_[14][0][240],
B_[14][1][240],
B_[14][2][240],
B_[15][0][240],
B_[15][1][240],
B_[15][2][240],
B_[0][0][241],
B_[0][1][241],
B_[0][2][241],
B_[1][0][241],
B_[1][1][241],
B_[1][2][241],
B_[2][0][241],
B_[2][1][241],
B_[2][2][241],
B_[3][0][241],
B_[3][1][241],
B_[3][2][241],
B_[4][0][241],
B_[4][1][241],
B_[4][2][241],
B_[5][0][241],
B_[5][1][241],
B_[5][2][241],
B_[6][0][241],
B_[6][1][241],
B_[6][2][241],
B_[7][0][241],
B_[7][1][241],
B_[7][2][241],
B_[8][0][241],
B_[8][1][241],
B_[8][2][241],
B_[9][0][241],
B_[9][1][241],
B_[9][2][241],
B_[10][0][241],
B_[10][1][241],
B_[10][2][241],
B_[11][0][241],
B_[11][1][241],
B_[11][2][241],
B_[12][0][241],
B_[12][1][241],
B_[12][2][241],
B_[13][0][241],
B_[13][1][241],
B_[13][2][241],
B_[14][0][241],
B_[14][1][241],
B_[14][2][241],
B_[15][0][241],
B_[15][1][241],
B_[15][2][241],
B_[0][0][242],
B_[0][1][242],
B_[0][2][242],
B_[1][0][242],
B_[1][1][242],
B_[1][2][242],
B_[2][0][242],
B_[2][1][242],
B_[2][2][242],
B_[3][0][242],
B_[3][1][242],
B_[3][2][242],
B_[4][0][242],
B_[4][1][242],
B_[4][2][242],
B_[5][0][242],
B_[5][1][242],
B_[5][2][242],
B_[6][0][242],
B_[6][1][242],
B_[6][2][242],
B_[7][0][242],
B_[7][1][242],
B_[7][2][242],
B_[8][0][242],
B_[8][1][242],
B_[8][2][242],
B_[9][0][242],
B_[9][1][242],
B_[9][2][242],
B_[10][0][242],
B_[10][1][242],
B_[10][2][242],
B_[11][0][242],
B_[11][1][242],
B_[11][2][242],
B_[12][0][242],
B_[12][1][242],
B_[12][2][242],
B_[13][0][242],
B_[13][1][242],
B_[13][2][242],
B_[14][0][242],
B_[14][1][242],
B_[14][2][242],
B_[15][0][242],
B_[15][1][242],
B_[15][2][242],
B_[0][0][243],
B_[0][1][243],
B_[0][2][243],
B_[1][0][243],
B_[1][1][243],
B_[1][2][243],
B_[2][0][243],
B_[2][1][243],
B_[2][2][243],
B_[3][0][243],
B_[3][1][243],
B_[3][2][243],
B_[4][0][243],
B_[4][1][243],
B_[4][2][243],
B_[5][0][243],
B_[5][1][243],
B_[5][2][243],
B_[6][0][243],
B_[6][1][243],
B_[6][2][243],
B_[7][0][243],
B_[7][1][243],
B_[7][2][243],
B_[8][0][243],
B_[8][1][243],
B_[8][2][243],
B_[9][0][243],
B_[9][1][243],
B_[9][2][243],
B_[10][0][243],
B_[10][1][243],
B_[10][2][243],
B_[11][0][243],
B_[11][1][243],
B_[11][2][243],
B_[12][0][243],
B_[12][1][243],
B_[12][2][243],
B_[13][0][243],
B_[13][1][243],
B_[13][2][243],
B_[14][0][243],
B_[14][1][243],
B_[14][2][243],
B_[15][0][243],
B_[15][1][243],
B_[15][2][243],
B_[0][0][244],
B_[0][1][244],
B_[0][2][244],
B_[1][0][244],
B_[1][1][244],
B_[1][2][244],
B_[2][0][244],
B_[2][1][244],
B_[2][2][244],
B_[3][0][244],
B_[3][1][244],
B_[3][2][244],
B_[4][0][244],
B_[4][1][244],
B_[4][2][244],
B_[5][0][244],
B_[5][1][244],
B_[5][2][244],
B_[6][0][244],
B_[6][1][244],
B_[6][2][244],
B_[7][0][244],
B_[7][1][244],
B_[7][2][244],
B_[8][0][244],
B_[8][1][244],
B_[8][2][244],
B_[9][0][244],
B_[9][1][244],
B_[9][2][244],
B_[10][0][244],
B_[10][1][244],
B_[10][2][244],
B_[11][0][244],
B_[11][1][244],
B_[11][2][244],
B_[12][0][244],
B_[12][1][244],
B_[12][2][244],
B_[13][0][244],
B_[13][1][244],
B_[13][2][244],
B_[14][0][244],
B_[14][1][244],
B_[14][2][244],
B_[15][0][244],
B_[15][1][244],
B_[15][2][244],
B_[0][0][245],
B_[0][1][245],
B_[0][2][245],
B_[1][0][245],
B_[1][1][245],
B_[1][2][245],
B_[2][0][245],
B_[2][1][245],
B_[2][2][245],
B_[3][0][245],
B_[3][1][245],
B_[3][2][245],
B_[4][0][245],
B_[4][1][245],
B_[4][2][245],
B_[5][0][245],
B_[5][1][245],
B_[5][2][245],
B_[6][0][245],
B_[6][1][245],
B_[6][2][245],
B_[7][0][245],
B_[7][1][245],
B_[7][2][245],
B_[8][0][245],
B_[8][1][245],
B_[8][2][245],
B_[9][0][245],
B_[9][1][245],
B_[9][2][245],
B_[10][0][245],
B_[10][1][245],
B_[10][2][245],
B_[11][0][245],
B_[11][1][245],
B_[11][2][245],
B_[12][0][245],
B_[12][1][245],
B_[12][2][245],
B_[13][0][245],
B_[13][1][245],
B_[13][2][245],
B_[14][0][245],
B_[14][1][245],
B_[14][2][245],
B_[15][0][245],
B_[15][1][245],
B_[15][2][245],
B_[0][0][246],
B_[0][1][246],
B_[0][2][246],
B_[1][0][246],
B_[1][1][246],
B_[1][2][246],
B_[2][0][246],
B_[2][1][246],
B_[2][2][246],
B_[3][0][246],
B_[3][1][246],
B_[3][2][246],
B_[4][0][246],
B_[4][1][246],
B_[4][2][246],
B_[5][0][246],
B_[5][1][246],
B_[5][2][246],
B_[6][0][246],
B_[6][1][246],
B_[6][2][246],
B_[7][0][246],
B_[7][1][246],
B_[7][2][246],
B_[8][0][246],
B_[8][1][246],
B_[8][2][246],
B_[9][0][246],
B_[9][1][246],
B_[9][2][246],
B_[10][0][246],
B_[10][1][246],
B_[10][2][246],
B_[11][0][246],
B_[11][1][246],
B_[11][2][246],
B_[12][0][246],
B_[12][1][246],
B_[12][2][246],
B_[13][0][246],
B_[13][1][246],
B_[13][2][246],
B_[14][0][246],
B_[14][1][246],
B_[14][2][246],
B_[15][0][246],
B_[15][1][246],
B_[15][2][246],
B_[0][0][247],
B_[0][1][247],
B_[0][2][247],
B_[1][0][247],
B_[1][1][247],
B_[1][2][247],
B_[2][0][247],
B_[2][1][247],
B_[2][2][247],
B_[3][0][247],
B_[3][1][247],
B_[3][2][247],
B_[4][0][247],
B_[4][1][247],
B_[4][2][247],
B_[5][0][247],
B_[5][1][247],
B_[5][2][247],
B_[6][0][247],
B_[6][1][247],
B_[6][2][247],
B_[7][0][247],
B_[7][1][247],
B_[7][2][247],
B_[8][0][247],
B_[8][1][247],
B_[8][2][247],
B_[9][0][247],
B_[9][1][247],
B_[9][2][247],
B_[10][0][247],
B_[10][1][247],
B_[10][2][247],
B_[11][0][247],
B_[11][1][247],
B_[11][2][247],
B_[12][0][247],
B_[12][1][247],
B_[12][2][247],
B_[13][0][247],
B_[13][1][247],
B_[13][2][247],
B_[14][0][247],
B_[14][1][247],
B_[14][2][247],
B_[15][0][247],
B_[15][1][247],
B_[15][2][247],
B_[0][0][248],
B_[0][1][248],
B_[0][2][248],
B_[1][0][248],
B_[1][1][248],
B_[1][2][248],
B_[2][0][248],
B_[2][1][248],
B_[2][2][248],
B_[3][0][248],
B_[3][1][248],
B_[3][2][248],
B_[4][0][248],
B_[4][1][248],
B_[4][2][248],
B_[5][0][248],
B_[5][1][248],
B_[5][2][248],
B_[6][0][248],
B_[6][1][248],
B_[6][2][248],
B_[7][0][248],
B_[7][1][248],
B_[7][2][248],
B_[8][0][248],
B_[8][1][248],
B_[8][2][248],
B_[9][0][248],
B_[9][1][248],
B_[9][2][248],
B_[10][0][248],
B_[10][1][248],
B_[10][2][248],
B_[11][0][248],
B_[11][1][248],
B_[11][2][248],
B_[12][0][248],
B_[12][1][248],
B_[12][2][248],
B_[13][0][248],
B_[13][1][248],
B_[13][2][248],
B_[14][0][248],
B_[14][1][248],
B_[14][2][248],
B_[15][0][248],
B_[15][1][248],
B_[15][2][248],
B_[0][0][249],
B_[0][1][249],
B_[0][2][249],
B_[1][0][249],
B_[1][1][249],
B_[1][2][249],
B_[2][0][249],
B_[2][1][249],
B_[2][2][249],
B_[3][0][249],
B_[3][1][249],
B_[3][2][249],
B_[4][0][249],
B_[4][1][249],
B_[4][2][249],
B_[5][0][249],
B_[5][1][249],
B_[5][2][249],
B_[6][0][249],
B_[6][1][249],
B_[6][2][249],
B_[7][0][249],
B_[7][1][249],
B_[7][2][249],
B_[8][0][249],
B_[8][1][249],
B_[8][2][249],
B_[9][0][249],
B_[9][1][249],
B_[9][2][249],
B_[10][0][249],
B_[10][1][249],
B_[10][2][249],
B_[11][0][249],
B_[11][1][249],
B_[11][2][249],
B_[12][0][249],
B_[12][1][249],
B_[12][2][249],
B_[13][0][249],
B_[13][1][249],
B_[13][2][249],
B_[14][0][249],
B_[14][1][249],
B_[14][2][249],
B_[15][0][249],
B_[15][1][249],
B_[15][2][249],
B_[0][0][250],
B_[0][1][250],
B_[0][2][250],
B_[1][0][250],
B_[1][1][250],
B_[1][2][250],
B_[2][0][250],
B_[2][1][250],
B_[2][2][250],
B_[3][0][250],
B_[3][1][250],
B_[3][2][250],
B_[4][0][250],
B_[4][1][250],
B_[4][2][250],
B_[5][0][250],
B_[5][1][250],
B_[5][2][250],
B_[6][0][250],
B_[6][1][250],
B_[6][2][250],
B_[7][0][250],
B_[7][1][250],
B_[7][2][250],
B_[8][0][250],
B_[8][1][250],
B_[8][2][250],
B_[9][0][250],
B_[9][1][250],
B_[9][2][250],
B_[10][0][250],
B_[10][1][250],
B_[10][2][250],
B_[11][0][250],
B_[11][1][250],
B_[11][2][250],
B_[12][0][250],
B_[12][1][250],
B_[12][2][250],
B_[13][0][250],
B_[13][1][250],
B_[13][2][250],
B_[14][0][250],
B_[14][1][250],
B_[14][2][250],
B_[15][0][250],
B_[15][1][250],
B_[15][2][250],
B_[0][0][251],
B_[0][1][251],
B_[0][2][251],
B_[1][0][251],
B_[1][1][251],
B_[1][2][251],
B_[2][0][251],
B_[2][1][251],
B_[2][2][251],
B_[3][0][251],
B_[3][1][251],
B_[3][2][251],
B_[4][0][251],
B_[4][1][251],
B_[4][2][251],
B_[5][0][251],
B_[5][1][251],
B_[5][2][251],
B_[6][0][251],
B_[6][1][251],
B_[6][2][251],
B_[7][0][251],
B_[7][1][251],
B_[7][2][251],
B_[8][0][251],
B_[8][1][251],
B_[8][2][251],
B_[9][0][251],
B_[9][1][251],
B_[9][2][251],
B_[10][0][251],
B_[10][1][251],
B_[10][2][251],
B_[11][0][251],
B_[11][1][251],
B_[11][2][251],
B_[12][0][251],
B_[12][1][251],
B_[12][2][251],
B_[13][0][251],
B_[13][1][251],
B_[13][2][251],
B_[14][0][251],
B_[14][1][251],
B_[14][2][251],
B_[15][0][251],
B_[15][1][251],
B_[15][2][251],
B_[0][0][252],
B_[0][1][252],
B_[0][2][252],
B_[1][0][252],
B_[1][1][252],
B_[1][2][252],
B_[2][0][252],
B_[2][1][252],
B_[2][2][252],
B_[3][0][252],
B_[3][1][252],
B_[3][2][252],
B_[4][0][252],
B_[4][1][252],
B_[4][2][252],
B_[5][0][252],
B_[5][1][252],
B_[5][2][252],
B_[6][0][252],
B_[6][1][252],
B_[6][2][252],
B_[7][0][252],
B_[7][1][252],
B_[7][2][252],
B_[8][0][252],
B_[8][1][252],
B_[8][2][252],
B_[9][0][252],
B_[9][1][252],
B_[9][2][252],
B_[10][0][252],
B_[10][1][252],
B_[10][2][252],
B_[11][0][252],
B_[11][1][252],
B_[11][2][252],
B_[12][0][252],
B_[12][1][252],
B_[12][2][252],
B_[13][0][252],
B_[13][1][252],
B_[13][2][252],
B_[14][0][252],
B_[14][1][252],
B_[14][2][252],
B_[15][0][252],
B_[15][1][252],
B_[15][2][252],
B_[0][0][253],
B_[0][1][253],
B_[0][2][253],
B_[1][0][253],
B_[1][1][253],
B_[1][2][253],
B_[2][0][253],
B_[2][1][253],
B_[2][2][253],
B_[3][0][253],
B_[3][1][253],
B_[3][2][253],
B_[4][0][253],
B_[4][1][253],
B_[4][2][253],
B_[5][0][253],
B_[5][1][253],
B_[5][2][253],
B_[6][0][253],
B_[6][1][253],
B_[6][2][253],
B_[7][0][253],
B_[7][1][253],
B_[7][2][253],
B_[8][0][253],
B_[8][1][253],
B_[8][2][253],
B_[9][0][253],
B_[9][1][253],
B_[9][2][253],
B_[10][0][253],
B_[10][1][253],
B_[10][2][253],
B_[11][0][253],
B_[11][1][253],
B_[11][2][253],
B_[12][0][253],
B_[12][1][253],
B_[12][2][253],
B_[13][0][253],
B_[13][1][253],
B_[13][2][253],
B_[14][0][253],
B_[14][1][253],
B_[14][2][253],
B_[15][0][253],
B_[15][1][253],
B_[15][2][253],
B_[0][0][254],
B_[0][1][254],
B_[0][2][254],
B_[1][0][254],
B_[1][1][254],
B_[1][2][254],
B_[2][0][254],
B_[2][1][254],
B_[2][2][254],
B_[3][0][254],
B_[3][1][254],
B_[3][2][254],
B_[4][0][254],
B_[4][1][254],
B_[4][2][254],
B_[5][0][254],
B_[5][1][254],
B_[5][2][254],
B_[6][0][254],
B_[6][1][254],
B_[6][2][254],
B_[7][0][254],
B_[7][1][254],
B_[7][2][254],
B_[8][0][254],
B_[8][1][254],
B_[8][2][254],
B_[9][0][254],
B_[9][1][254],
B_[9][2][254],
B_[10][0][254],
B_[10][1][254],
B_[10][2][254],
B_[11][0][254],
B_[11][1][254],
B_[11][2][254],
B_[12][0][254],
B_[12][1][254],
B_[12][2][254],
B_[13][0][254],
B_[13][1][254],
B_[13][2][254],
B_[14][0][254],
B_[14][1][254],
B_[14][2][254],
B_[15][0][254],
B_[15][1][254],
B_[15][2][254],
B_[0][0][255],
B_[0][1][255],
B_[0][2][255],
B_[1][0][255],
B_[1][1][255],
B_[1][2][255],
B_[2][0][255],
B_[2][1][255],
B_[2][2][255],
B_[3][0][255],
B_[3][1][255],
B_[3][2][255],
B_[4][0][255],
B_[4][1][255],
B_[4][2][255],
B_[5][0][255],
B_[5][1][255],
B_[5][2][255],
B_[6][0][255],
B_[6][1][255],
B_[6][2][255],
B_[7][0][255],
B_[7][1][255],
B_[7][2][255],
B_[8][0][255],
B_[8][1][255],
B_[8][2][255],
B_[9][0][255],
B_[9][1][255],
B_[9][2][255],
B_[10][0][255],
B_[10][1][255],
B_[10][2][255],
B_[11][0][255],
B_[11][1][255],
B_[11][2][255],
B_[12][0][255],
B_[12][1][255],
B_[12][2][255],
B_[13][0][255],
B_[13][1][255],
B_[13][2][255],
B_[14][0][255],
B_[14][1][255],
B_[14][2][255],
B_[15][0][255],
B_[15][1][255],
B_[15][2][255],
F_[0][0][0],
F_[0][1][0],
F_[0][2][0],
F_[1][0][0],
F_[1][1][0],
F_[1][2][0],
F_[2][0][0],
F_[2][1][0],
F_[2][2][0],
F_[3][0][0],
F_[3][1][0],
F_[3][2][0],
F_[4][0][0],
F_[4][1][0],
F_[4][2][0],
F_[5][0][0],
F_[5][1][0],
F_[5][2][0],
F_[6][0][0],
F_[6][1][0],
F_[6][2][0],
F_[7][0][0],
F_[7][1][0],
F_[7][2][0],
F_[8][0][0],
F_[8][1][0],
F_[8][2][0],
F_[9][0][0],
F_[9][1][0],
F_[9][2][0],
F_[10][0][0],
F_[10][1][0],
F_[10][2][0],
F_[11][0][0],
F_[11][1][0],
F_[11][2][0],
F_[12][0][0],
F_[12][1][0],
F_[12][2][0],
F_[13][0][0],
F_[13][1][0],
F_[13][2][0],
F_[14][0][0],
F_[14][1][0],
F_[14][2][0],
F_[15][0][0],
F_[15][1][0],
F_[15][2][0],
F_[0][0][1],
F_[0][1][1],
F_[0][2][1],
F_[1][0][1],
F_[1][1][1],
F_[1][2][1],
F_[2][0][1],
F_[2][1][1],
F_[2][2][1],
F_[3][0][1],
F_[3][1][1],
F_[3][2][1],
F_[4][0][1],
F_[4][1][1],
F_[4][2][1],
F_[5][0][1],
F_[5][1][1],
F_[5][2][1],
F_[6][0][1],
F_[6][1][1],
F_[6][2][1],
F_[7][0][1],
F_[7][1][1],
F_[7][2][1],
F_[8][0][1],
F_[8][1][1],
F_[8][2][1],
F_[9][0][1],
F_[9][1][1],
F_[9][2][1],
F_[10][0][1],
F_[10][1][1],
F_[10][2][1],
F_[11][0][1],
F_[11][1][1],
F_[11][2][1],
F_[12][0][1],
F_[12][1][1],
F_[12][2][1],
F_[13][0][1],
F_[13][1][1],
F_[13][2][1],
F_[14][0][1],
F_[14][1][1],
F_[14][2][1],
F_[15][0][1],
F_[15][1][1],
F_[15][2][1],
F_[0][0][2],
F_[0][1][2],
F_[0][2][2],
F_[1][0][2],
F_[1][1][2],
F_[1][2][2],
F_[2][0][2],
F_[2][1][2],
F_[2][2][2],
F_[3][0][2],
F_[3][1][2],
F_[3][2][2],
F_[4][0][2],
F_[4][1][2],
F_[4][2][2],
F_[5][0][2],
F_[5][1][2],
F_[5][2][2],
F_[6][0][2],
F_[6][1][2],
F_[6][2][2],
F_[7][0][2],
F_[7][1][2],
F_[7][2][2],
F_[8][0][2],
F_[8][1][2],
F_[8][2][2],
F_[9][0][2],
F_[9][1][2],
F_[9][2][2],
F_[10][0][2],
F_[10][1][2],
F_[10][2][2],
F_[11][0][2],
F_[11][1][2],
F_[11][2][2],
F_[12][0][2],
F_[12][1][2],
F_[12][2][2],
F_[13][0][2],
F_[13][1][2],
F_[13][2][2],
F_[14][0][2],
F_[14][1][2],
F_[14][2][2],
F_[15][0][2],
F_[15][1][2],
F_[15][2][2],
F_[0][0][3],
F_[0][1][3],
F_[0][2][3],
F_[1][0][3],
F_[1][1][3],
F_[1][2][3],
F_[2][0][3],
F_[2][1][3],
F_[2][2][3],
F_[3][0][3],
F_[3][1][3],
F_[3][2][3],
F_[4][0][3],
F_[4][1][3],
F_[4][2][3],
F_[5][0][3],
F_[5][1][3],
F_[5][2][3],
F_[6][0][3],
F_[6][1][3],
F_[6][2][3],
F_[7][0][3],
F_[7][1][3],
F_[7][2][3],
F_[8][0][3],
F_[8][1][3],
F_[8][2][3],
F_[9][0][3],
F_[9][1][3],
F_[9][2][3],
F_[10][0][3],
F_[10][1][3],
F_[10][2][3],
F_[11][0][3],
F_[11][1][3],
F_[11][2][3],
F_[12][0][3],
F_[12][1][3],
F_[12][2][3],
F_[13][0][3],
F_[13][1][3],
F_[13][2][3],
F_[14][0][3],
F_[14][1][3],
F_[14][2][3],
F_[15][0][3],
F_[15][1][3],
F_[15][2][3],
F_[0][0][4],
F_[0][1][4],
F_[0][2][4],
F_[1][0][4],
F_[1][1][4],
F_[1][2][4],
F_[2][0][4],
F_[2][1][4],
F_[2][2][4],
F_[3][0][4],
F_[3][1][4],
F_[3][2][4],
F_[4][0][4],
F_[4][1][4],
F_[4][2][4],
F_[5][0][4],
F_[5][1][4],
F_[5][2][4],
F_[6][0][4],
F_[6][1][4],
F_[6][2][4],
F_[7][0][4],
F_[7][1][4],
F_[7][2][4],
F_[8][0][4],
F_[8][1][4],
F_[8][2][4],
F_[9][0][4],
F_[9][1][4],
F_[9][2][4],
F_[10][0][4],
F_[10][1][4],
F_[10][2][4],
F_[11][0][4],
F_[11][1][4],
F_[11][2][4],
F_[12][0][4],
F_[12][1][4],
F_[12][2][4],
F_[13][0][4],
F_[13][1][4],
F_[13][2][4],
F_[14][0][4],
F_[14][1][4],
F_[14][2][4],
F_[15][0][4],
F_[15][1][4],
F_[15][2][4],
F_[0][0][5],
F_[0][1][5],
F_[0][2][5],
F_[1][0][5],
F_[1][1][5],
F_[1][2][5],
F_[2][0][5],
F_[2][1][5],
F_[2][2][5],
F_[3][0][5],
F_[3][1][5],
F_[3][2][5],
F_[4][0][5],
F_[4][1][5],
F_[4][2][5],
F_[5][0][5],
F_[5][1][5],
F_[5][2][5],
F_[6][0][5],
F_[6][1][5],
F_[6][2][5],
F_[7][0][5],
F_[7][1][5],
F_[7][2][5],
F_[8][0][5],
F_[8][1][5],
F_[8][2][5],
F_[9][0][5],
F_[9][1][5],
F_[9][2][5],
F_[10][0][5],
F_[10][1][5],
F_[10][2][5],
F_[11][0][5],
F_[11][1][5],
F_[11][2][5],
F_[12][0][5],
F_[12][1][5],
F_[12][2][5],
F_[13][0][5],
F_[13][1][5],
F_[13][2][5],
F_[14][0][5],
F_[14][1][5],
F_[14][2][5],
F_[15][0][5],
F_[15][1][5],
F_[15][2][5],
F_[0][0][6],
F_[0][1][6],
F_[0][2][6],
F_[1][0][6],
F_[1][1][6],
F_[1][2][6],
F_[2][0][6],
F_[2][1][6],
F_[2][2][6],
F_[3][0][6],
F_[3][1][6],
F_[3][2][6],
F_[4][0][6],
F_[4][1][6],
F_[4][2][6],
F_[5][0][6],
F_[5][1][6],
F_[5][2][6],
F_[6][0][6],
F_[6][1][6],
F_[6][2][6],
F_[7][0][6],
F_[7][1][6],
F_[7][2][6],
F_[8][0][6],
F_[8][1][6],
F_[8][2][6],
F_[9][0][6],
F_[9][1][6],
F_[9][2][6],
F_[10][0][6],
F_[10][1][6],
F_[10][2][6],
F_[11][0][6],
F_[11][1][6],
F_[11][2][6],
F_[12][0][6],
F_[12][1][6],
F_[12][2][6],
F_[13][0][6],
F_[13][1][6],
F_[13][2][6],
F_[14][0][6],
F_[14][1][6],
F_[14][2][6],
F_[15][0][6],
F_[15][1][6],
F_[15][2][6],
F_[0][0][7],
F_[0][1][7],
F_[0][2][7],
F_[1][0][7],
F_[1][1][7],
F_[1][2][7],
F_[2][0][7],
F_[2][1][7],
F_[2][2][7],
F_[3][0][7],
F_[3][1][7],
F_[3][2][7],
F_[4][0][7],
F_[4][1][7],
F_[4][2][7],
F_[5][0][7],
F_[5][1][7],
F_[5][2][7],
F_[6][0][7],
F_[6][1][7],
F_[6][2][7],
F_[7][0][7],
F_[7][1][7],
F_[7][2][7],
F_[8][0][7],
F_[8][1][7],
F_[8][2][7],
F_[9][0][7],
F_[9][1][7],
F_[9][2][7],
F_[10][0][7],
F_[10][1][7],
F_[10][2][7],
F_[11][0][7],
F_[11][1][7],
F_[11][2][7],
F_[12][0][7],
F_[12][1][7],
F_[12][2][7],
F_[13][0][7],
F_[13][1][7],
F_[13][2][7],
F_[14][0][7],
F_[14][1][7],
F_[14][2][7],
F_[15][0][7],
F_[15][1][7],
F_[15][2][7],
F_[0][0][8],
F_[0][1][8],
F_[0][2][8],
F_[1][0][8],
F_[1][1][8],
F_[1][2][8],
F_[2][0][8],
F_[2][1][8],
F_[2][2][8],
F_[3][0][8],
F_[3][1][8],
F_[3][2][8],
F_[4][0][8],
F_[4][1][8],
F_[4][2][8],
F_[5][0][8],
F_[5][1][8],
F_[5][2][8],
F_[6][0][8],
F_[6][1][8],
F_[6][2][8],
F_[7][0][8],
F_[7][1][8],
F_[7][2][8],
F_[8][0][8],
F_[8][1][8],
F_[8][2][8],
F_[9][0][8],
F_[9][1][8],
F_[9][2][8],
F_[10][0][8],
F_[10][1][8],
F_[10][2][8],
F_[11][0][8],
F_[11][1][8],
F_[11][2][8],
F_[12][0][8],
F_[12][1][8],
F_[12][2][8],
F_[13][0][8],
F_[13][1][8],
F_[13][2][8],
F_[14][0][8],
F_[14][1][8],
F_[14][2][8],
F_[15][0][8],
F_[15][1][8],
F_[15][2][8],
F_[0][0][9],
F_[0][1][9],
F_[0][2][9],
F_[1][0][9],
F_[1][1][9],
F_[1][2][9],
F_[2][0][9],
F_[2][1][9],
F_[2][2][9],
F_[3][0][9],
F_[3][1][9],
F_[3][2][9],
F_[4][0][9],
F_[4][1][9],
F_[4][2][9],
F_[5][0][9],
F_[5][1][9],
F_[5][2][9],
F_[6][0][9],
F_[6][1][9],
F_[6][2][9],
F_[7][0][9],
F_[7][1][9],
F_[7][2][9],
F_[8][0][9],
F_[8][1][9],
F_[8][2][9],
F_[9][0][9],
F_[9][1][9],
F_[9][2][9],
F_[10][0][9],
F_[10][1][9],
F_[10][2][9],
F_[11][0][9],
F_[11][1][9],
F_[11][2][9],
F_[12][0][9],
F_[12][1][9],
F_[12][2][9],
F_[13][0][9],
F_[13][1][9],
F_[13][2][9],
F_[14][0][9],
F_[14][1][9],
F_[14][2][9],
F_[15][0][9],
F_[15][1][9],
F_[15][2][9],
F_[0][0][10],
F_[0][1][10],
F_[0][2][10],
F_[1][0][10],
F_[1][1][10],
F_[1][2][10],
F_[2][0][10],
F_[2][1][10],
F_[2][2][10],
F_[3][0][10],
F_[3][1][10],
F_[3][2][10],
F_[4][0][10],
F_[4][1][10],
F_[4][2][10],
F_[5][0][10],
F_[5][1][10],
F_[5][2][10],
F_[6][0][10],
F_[6][1][10],
F_[6][2][10],
F_[7][0][10],
F_[7][1][10],
F_[7][2][10],
F_[8][0][10],
F_[8][1][10],
F_[8][2][10],
F_[9][0][10],
F_[9][1][10],
F_[9][2][10],
F_[10][0][10],
F_[10][1][10],
F_[10][2][10],
F_[11][0][10],
F_[11][1][10],
F_[11][2][10],
F_[12][0][10],
F_[12][1][10],
F_[12][2][10],
F_[13][0][10],
F_[13][1][10],
F_[13][2][10],
F_[14][0][10],
F_[14][1][10],
F_[14][2][10],
F_[15][0][10],
F_[15][1][10],
F_[15][2][10],
F_[0][0][11],
F_[0][1][11],
F_[0][2][11],
F_[1][0][11],
F_[1][1][11],
F_[1][2][11],
F_[2][0][11],
F_[2][1][11],
F_[2][2][11],
F_[3][0][11],
F_[3][1][11],
F_[3][2][11],
F_[4][0][11],
F_[4][1][11],
F_[4][2][11],
F_[5][0][11],
F_[5][1][11],
F_[5][2][11],
F_[6][0][11],
F_[6][1][11],
F_[6][2][11],
F_[7][0][11],
F_[7][1][11],
F_[7][2][11],
F_[8][0][11],
F_[8][1][11],
F_[8][2][11],
F_[9][0][11],
F_[9][1][11],
F_[9][2][11],
F_[10][0][11],
F_[10][1][11],
F_[10][2][11],
F_[11][0][11],
F_[11][1][11],
F_[11][2][11],
F_[12][0][11],
F_[12][1][11],
F_[12][2][11],
F_[13][0][11],
F_[13][1][11],
F_[13][2][11],
F_[14][0][11],
F_[14][1][11],
F_[14][2][11],
F_[15][0][11],
F_[15][1][11],
F_[15][2][11],
F_[0][0][12],
F_[0][1][12],
F_[0][2][12],
F_[1][0][12],
F_[1][1][12],
F_[1][2][12],
F_[2][0][12],
F_[2][1][12],
F_[2][2][12],
F_[3][0][12],
F_[3][1][12],
F_[3][2][12],
F_[4][0][12],
F_[4][1][12],
F_[4][2][12],
F_[5][0][12],
F_[5][1][12],
F_[5][2][12],
F_[6][0][12],
F_[6][1][12],
F_[6][2][12],
F_[7][0][12],
F_[7][1][12],
F_[7][2][12],
F_[8][0][12],
F_[8][1][12],
F_[8][2][12],
F_[9][0][12],
F_[9][1][12],
F_[9][2][12],
F_[10][0][12],
F_[10][1][12],
F_[10][2][12],
F_[11][0][12],
F_[11][1][12],
F_[11][2][12],
F_[12][0][12],
F_[12][1][12],
F_[12][2][12],
F_[13][0][12],
F_[13][1][12],
F_[13][2][12],
F_[14][0][12],
F_[14][1][12],
F_[14][2][12],
F_[15][0][12],
F_[15][1][12],
F_[15][2][12],
F_[0][0][13],
F_[0][1][13],
F_[0][2][13],
F_[1][0][13],
F_[1][1][13],
F_[1][2][13],
F_[2][0][13],
F_[2][1][13],
F_[2][2][13],
F_[3][0][13],
F_[3][1][13],
F_[3][2][13],
F_[4][0][13],
F_[4][1][13],
F_[4][2][13],
F_[5][0][13],
F_[5][1][13],
F_[5][2][13],
F_[6][0][13],
F_[6][1][13],
F_[6][2][13],
F_[7][0][13],
F_[7][1][13],
F_[7][2][13],
F_[8][0][13],
F_[8][1][13],
F_[8][2][13],
F_[9][0][13],
F_[9][1][13],
F_[9][2][13],
F_[10][0][13],
F_[10][1][13],
F_[10][2][13],
F_[11][0][13],
F_[11][1][13],
F_[11][2][13],
F_[12][0][13],
F_[12][1][13],
F_[12][2][13],
F_[13][0][13],
F_[13][1][13],
F_[13][2][13],
F_[14][0][13],
F_[14][1][13],
F_[14][2][13],
F_[15][0][13],
F_[15][1][13],
F_[15][2][13],
F_[0][0][14],
F_[0][1][14],
F_[0][2][14],
F_[1][0][14],
F_[1][1][14],
F_[1][2][14],
F_[2][0][14],
F_[2][1][14],
F_[2][2][14],
F_[3][0][14],
F_[3][1][14],
F_[3][2][14],
F_[4][0][14],
F_[4][1][14],
F_[4][2][14],
F_[5][0][14],
F_[5][1][14],
F_[5][2][14],
F_[6][0][14],
F_[6][1][14],
F_[6][2][14],
F_[7][0][14],
F_[7][1][14],
F_[7][2][14],
F_[8][0][14],
F_[8][1][14],
F_[8][2][14],
F_[9][0][14],
F_[9][1][14],
F_[9][2][14],
F_[10][0][14],
F_[10][1][14],
F_[10][2][14],
F_[11][0][14],
F_[11][1][14],
F_[11][2][14],
F_[12][0][14],
F_[12][1][14],
F_[12][2][14],
F_[13][0][14],
F_[13][1][14],
F_[13][2][14],
F_[14][0][14],
F_[14][1][14],
F_[14][2][14],
F_[15][0][14],
F_[15][1][14],
F_[15][2][14],
F_[0][0][15],
F_[0][1][15],
F_[0][2][15],
F_[1][0][15],
F_[1][1][15],
F_[1][2][15],
F_[2][0][15],
F_[2][1][15],
F_[2][2][15],
F_[3][0][15],
F_[3][1][15],
F_[3][2][15],
F_[4][0][15],
F_[4][1][15],
F_[4][2][15],
F_[5][0][15],
F_[5][1][15],
F_[5][2][15],
F_[6][0][15],
F_[6][1][15],
F_[6][2][15],
F_[7][0][15],
F_[7][1][15],
F_[7][2][15],
F_[8][0][15],
F_[8][1][15],
F_[8][2][15],
F_[9][0][15],
F_[9][1][15],
F_[9][2][15],
F_[10][0][15],
F_[10][1][15],
F_[10][2][15],
F_[11][0][15],
F_[11][1][15],
F_[11][2][15],
F_[12][0][15],
F_[12][1][15],
F_[12][2][15],
F_[13][0][15],
F_[13][1][15],
F_[13][2][15],
F_[14][0][15],
F_[14][1][15],
F_[14][2][15],
F_[15][0][15],
F_[15][1][15],
F_[15][2][15],
F_[0][0][16],
F_[0][1][16],
F_[0][2][16],
F_[1][0][16],
F_[1][1][16],
F_[1][2][16],
F_[2][0][16],
F_[2][1][16],
F_[2][2][16],
F_[3][0][16],
F_[3][1][16],
F_[3][2][16],
F_[4][0][16],
F_[4][1][16],
F_[4][2][16],
F_[5][0][16],
F_[5][1][16],
F_[5][2][16],
F_[6][0][16],
F_[6][1][16],
F_[6][2][16],
F_[7][0][16],
F_[7][1][16],
F_[7][2][16],
F_[8][0][16],
F_[8][1][16],
F_[8][2][16],
F_[9][0][16],
F_[9][1][16],
F_[9][2][16],
F_[10][0][16],
F_[10][1][16],
F_[10][2][16],
F_[11][0][16],
F_[11][1][16],
F_[11][2][16],
F_[12][0][16],
F_[12][1][16],
F_[12][2][16],
F_[13][0][16],
F_[13][1][16],
F_[13][2][16],
F_[14][0][16],
F_[14][1][16],
F_[14][2][16],
F_[15][0][16],
F_[15][1][16],
F_[15][2][16],
F_[0][0][17],
F_[0][1][17],
F_[0][2][17],
F_[1][0][17],
F_[1][1][17],
F_[1][2][17],
F_[2][0][17],
F_[2][1][17],
F_[2][2][17],
F_[3][0][17],
F_[3][1][17],
F_[3][2][17],
F_[4][0][17],
F_[4][1][17],
F_[4][2][17],
F_[5][0][17],
F_[5][1][17],
F_[5][2][17],
F_[6][0][17],
F_[6][1][17],
F_[6][2][17],
F_[7][0][17],
F_[7][1][17],
F_[7][2][17],
F_[8][0][17],
F_[8][1][17],
F_[8][2][17],
F_[9][0][17],
F_[9][1][17],
F_[9][2][17],
F_[10][0][17],
F_[10][1][17],
F_[10][2][17],
F_[11][0][17],
F_[11][1][17],
F_[11][2][17],
F_[12][0][17],
F_[12][1][17],
F_[12][2][17],
F_[13][0][17],
F_[13][1][17],
F_[13][2][17],
F_[14][0][17],
F_[14][1][17],
F_[14][2][17],
F_[15][0][17],
F_[15][1][17],
F_[15][2][17],
F_[0][0][18],
F_[0][1][18],
F_[0][2][18],
F_[1][0][18],
F_[1][1][18],
F_[1][2][18],
F_[2][0][18],
F_[2][1][18],
F_[2][2][18],
F_[3][0][18],
F_[3][1][18],
F_[3][2][18],
F_[4][0][18],
F_[4][1][18],
F_[4][2][18],
F_[5][0][18],
F_[5][1][18],
F_[5][2][18],
F_[6][0][18],
F_[6][1][18],
F_[6][2][18],
F_[7][0][18],
F_[7][1][18],
F_[7][2][18],
F_[8][0][18],
F_[8][1][18],
F_[8][2][18],
F_[9][0][18],
F_[9][1][18],
F_[9][2][18],
F_[10][0][18],
F_[10][1][18],
F_[10][2][18],
F_[11][0][18],
F_[11][1][18],
F_[11][2][18],
F_[12][0][18],
F_[12][1][18],
F_[12][2][18],
F_[13][0][18],
F_[13][1][18],
F_[13][2][18],
F_[14][0][18],
F_[14][1][18],
F_[14][2][18],
F_[15][0][18],
F_[15][1][18],
F_[15][2][18],
F_[0][0][19],
F_[0][1][19],
F_[0][2][19],
F_[1][0][19],
F_[1][1][19],
F_[1][2][19],
F_[2][0][19],
F_[2][1][19],
F_[2][2][19],
F_[3][0][19],
F_[3][1][19],
F_[3][2][19],
F_[4][0][19],
F_[4][1][19],
F_[4][2][19],
F_[5][0][19],
F_[5][1][19],
F_[5][2][19],
F_[6][0][19],
F_[6][1][19],
F_[6][2][19],
F_[7][0][19],
F_[7][1][19],
F_[7][2][19],
F_[8][0][19],
F_[8][1][19],
F_[8][2][19],
F_[9][0][19],
F_[9][1][19],
F_[9][2][19],
F_[10][0][19],
F_[10][1][19],
F_[10][2][19],
F_[11][0][19],
F_[11][1][19],
F_[11][2][19],
F_[12][0][19],
F_[12][1][19],
F_[12][2][19],
F_[13][0][19],
F_[13][1][19],
F_[13][2][19],
F_[14][0][19],
F_[14][1][19],
F_[14][2][19],
F_[15][0][19],
F_[15][1][19],
F_[15][2][19],
F_[0][0][20],
F_[0][1][20],
F_[0][2][20],
F_[1][0][20],
F_[1][1][20],
F_[1][2][20],
F_[2][0][20],
F_[2][1][20],
F_[2][2][20],
F_[3][0][20],
F_[3][1][20],
F_[3][2][20],
F_[4][0][20],
F_[4][1][20],
F_[4][2][20],
F_[5][0][20],
F_[5][1][20],
F_[5][2][20],
F_[6][0][20],
F_[6][1][20],
F_[6][2][20],
F_[7][0][20],
F_[7][1][20],
F_[7][2][20],
F_[8][0][20],
F_[8][1][20],
F_[8][2][20],
F_[9][0][20],
F_[9][1][20],
F_[9][2][20],
F_[10][0][20],
F_[10][1][20],
F_[10][2][20],
F_[11][0][20],
F_[11][1][20],
F_[11][2][20],
F_[12][0][20],
F_[12][1][20],
F_[12][2][20],
F_[13][0][20],
F_[13][1][20],
F_[13][2][20],
F_[14][0][20],
F_[14][1][20],
F_[14][2][20],
F_[15][0][20],
F_[15][1][20],
F_[15][2][20],
F_[0][0][21],
F_[0][1][21],
F_[0][2][21],
F_[1][0][21],
F_[1][1][21],
F_[1][2][21],
F_[2][0][21],
F_[2][1][21],
F_[2][2][21],
F_[3][0][21],
F_[3][1][21],
F_[3][2][21],
F_[4][0][21],
F_[4][1][21],
F_[4][2][21],
F_[5][0][21],
F_[5][1][21],
F_[5][2][21],
F_[6][0][21],
F_[6][1][21],
F_[6][2][21],
F_[7][0][21],
F_[7][1][21],
F_[7][2][21],
F_[8][0][21],
F_[8][1][21],
F_[8][2][21],
F_[9][0][21],
F_[9][1][21],
F_[9][2][21],
F_[10][0][21],
F_[10][1][21],
F_[10][2][21],
F_[11][0][21],
F_[11][1][21],
F_[11][2][21],
F_[12][0][21],
F_[12][1][21],
F_[12][2][21],
F_[13][0][21],
F_[13][1][21],
F_[13][2][21],
F_[14][0][21],
F_[14][1][21],
F_[14][2][21],
F_[15][0][21],
F_[15][1][21],
F_[15][2][21],
F_[0][0][22],
F_[0][1][22],
F_[0][2][22],
F_[1][0][22],
F_[1][1][22],
F_[1][2][22],
F_[2][0][22],
F_[2][1][22],
F_[2][2][22],
F_[3][0][22],
F_[3][1][22],
F_[3][2][22],
F_[4][0][22],
F_[4][1][22],
F_[4][2][22],
F_[5][0][22],
F_[5][1][22],
F_[5][2][22],
F_[6][0][22],
F_[6][1][22],
F_[6][2][22],
F_[7][0][22],
F_[7][1][22],
F_[7][2][22],
F_[8][0][22],
F_[8][1][22],
F_[8][2][22],
F_[9][0][22],
F_[9][1][22],
F_[9][2][22],
F_[10][0][22],
F_[10][1][22],
F_[10][2][22],
F_[11][0][22],
F_[11][1][22],
F_[11][2][22],
F_[12][0][22],
F_[12][1][22],
F_[12][2][22],
F_[13][0][22],
F_[13][1][22],
F_[13][2][22],
F_[14][0][22],
F_[14][1][22],
F_[14][2][22],
F_[15][0][22],
F_[15][1][22],
F_[15][2][22],
F_[0][0][23],
F_[0][1][23],
F_[0][2][23],
F_[1][0][23],
F_[1][1][23],
F_[1][2][23],
F_[2][0][23],
F_[2][1][23],
F_[2][2][23],
F_[3][0][23],
F_[3][1][23],
F_[3][2][23],
F_[4][0][23],
F_[4][1][23],
F_[4][2][23],
F_[5][0][23],
F_[5][1][23],
F_[5][2][23],
F_[6][0][23],
F_[6][1][23],
F_[6][2][23],
F_[7][0][23],
F_[7][1][23],
F_[7][2][23],
F_[8][0][23],
F_[8][1][23],
F_[8][2][23],
F_[9][0][23],
F_[9][1][23],
F_[9][2][23],
F_[10][0][23],
F_[10][1][23],
F_[10][2][23],
F_[11][0][23],
F_[11][1][23],
F_[11][2][23],
F_[12][0][23],
F_[12][1][23],
F_[12][2][23],
F_[13][0][23],
F_[13][1][23],
F_[13][2][23],
F_[14][0][23],
F_[14][1][23],
F_[14][2][23],
F_[15][0][23],
F_[15][1][23],
F_[15][2][23],
F_[0][0][24],
F_[0][1][24],
F_[0][2][24],
F_[1][0][24],
F_[1][1][24],
F_[1][2][24],
F_[2][0][24],
F_[2][1][24],
F_[2][2][24],
F_[3][0][24],
F_[3][1][24],
F_[3][2][24],
F_[4][0][24],
F_[4][1][24],
F_[4][2][24],
F_[5][0][24],
F_[5][1][24],
F_[5][2][24],
F_[6][0][24],
F_[6][1][24],
F_[6][2][24],
F_[7][0][24],
F_[7][1][24],
F_[7][2][24],
F_[8][0][24],
F_[8][1][24],
F_[8][2][24],
F_[9][0][24],
F_[9][1][24],
F_[9][2][24],
F_[10][0][24],
F_[10][1][24],
F_[10][2][24],
F_[11][0][24],
F_[11][1][24],
F_[11][2][24],
F_[12][0][24],
F_[12][1][24],
F_[12][2][24],
F_[13][0][24],
F_[13][1][24],
F_[13][2][24],
F_[14][0][24],
F_[14][1][24],
F_[14][2][24],
F_[15][0][24],
F_[15][1][24],
F_[15][2][24],
F_[0][0][25],
F_[0][1][25],
F_[0][2][25],
F_[1][0][25],
F_[1][1][25],
F_[1][2][25],
F_[2][0][25],
F_[2][1][25],
F_[2][2][25],
F_[3][0][25],
F_[3][1][25],
F_[3][2][25],
F_[4][0][25],
F_[4][1][25],
F_[4][2][25],
F_[5][0][25],
F_[5][1][25],
F_[5][2][25],
F_[6][0][25],
F_[6][1][25],
F_[6][2][25],
F_[7][0][25],
F_[7][1][25],
F_[7][2][25],
F_[8][0][25],
F_[8][1][25],
F_[8][2][25],
F_[9][0][25],
F_[9][1][25],
F_[9][2][25],
F_[10][0][25],
F_[10][1][25],
F_[10][2][25],
F_[11][0][25],
F_[11][1][25],
F_[11][2][25],
F_[12][0][25],
F_[12][1][25],
F_[12][2][25],
F_[13][0][25],
F_[13][1][25],
F_[13][2][25],
F_[14][0][25],
F_[14][1][25],
F_[14][2][25],
F_[15][0][25],
F_[15][1][25],
F_[15][2][25],
F_[0][0][26],
F_[0][1][26],
F_[0][2][26],
F_[1][0][26],
F_[1][1][26],
F_[1][2][26],
F_[2][0][26],
F_[2][1][26],
F_[2][2][26],
F_[3][0][26],
F_[3][1][26],
F_[3][2][26],
F_[4][0][26],
F_[4][1][26],
F_[4][2][26],
F_[5][0][26],
F_[5][1][26],
F_[5][2][26],
F_[6][0][26],
F_[6][1][26],
F_[6][2][26],
F_[7][0][26],
F_[7][1][26],
F_[7][2][26],
F_[8][0][26],
F_[8][1][26],
F_[8][2][26],
F_[9][0][26],
F_[9][1][26],
F_[9][2][26],
F_[10][0][26],
F_[10][1][26],
F_[10][2][26],
F_[11][0][26],
F_[11][1][26],
F_[11][2][26],
F_[12][0][26],
F_[12][1][26],
F_[12][2][26],
F_[13][0][26],
F_[13][1][26],
F_[13][2][26],
F_[14][0][26],
F_[14][1][26],
F_[14][2][26],
F_[15][0][26],
F_[15][1][26],
F_[15][2][26],
F_[0][0][27],
F_[0][1][27],
F_[0][2][27],
F_[1][0][27],
F_[1][1][27],
F_[1][2][27],
F_[2][0][27],
F_[2][1][27],
F_[2][2][27],
F_[3][0][27],
F_[3][1][27],
F_[3][2][27],
F_[4][0][27],
F_[4][1][27],
F_[4][2][27],
F_[5][0][27],
F_[5][1][27],
F_[5][2][27],
F_[6][0][27],
F_[6][1][27],
F_[6][2][27],
F_[7][0][27],
F_[7][1][27],
F_[7][2][27],
F_[8][0][27],
F_[8][1][27],
F_[8][2][27],
F_[9][0][27],
F_[9][1][27],
F_[9][2][27],
F_[10][0][27],
F_[10][1][27],
F_[10][2][27],
F_[11][0][27],
F_[11][1][27],
F_[11][2][27],
F_[12][0][27],
F_[12][1][27],
F_[12][2][27],
F_[13][0][27],
F_[13][1][27],
F_[13][2][27],
F_[14][0][27],
F_[14][1][27],
F_[14][2][27],
F_[15][0][27],
F_[15][1][27],
F_[15][2][27],
F_[0][0][28],
F_[0][1][28],
F_[0][2][28],
F_[1][0][28],
F_[1][1][28],
F_[1][2][28],
F_[2][0][28],
F_[2][1][28],
F_[2][2][28],
F_[3][0][28],
F_[3][1][28],
F_[3][2][28],
F_[4][0][28],
F_[4][1][28],
F_[4][2][28],
F_[5][0][28],
F_[5][1][28],
F_[5][2][28],
F_[6][0][28],
F_[6][1][28],
F_[6][2][28],
F_[7][0][28],
F_[7][1][28],
F_[7][2][28],
F_[8][0][28],
F_[8][1][28],
F_[8][2][28],
F_[9][0][28],
F_[9][1][28],
F_[9][2][28],
F_[10][0][28],
F_[10][1][28],
F_[10][2][28],
F_[11][0][28],
F_[11][1][28],
F_[11][2][28],
F_[12][0][28],
F_[12][1][28],
F_[12][2][28],
F_[13][0][28],
F_[13][1][28],
F_[13][2][28],
F_[14][0][28],
F_[14][1][28],
F_[14][2][28],
F_[15][0][28],
F_[15][1][28],
F_[15][2][28],
F_[0][0][29],
F_[0][1][29],
F_[0][2][29],
F_[1][0][29],
F_[1][1][29],
F_[1][2][29],
F_[2][0][29],
F_[2][1][29],
F_[2][2][29],
F_[3][0][29],
F_[3][1][29],
F_[3][2][29],
F_[4][0][29],
F_[4][1][29],
F_[4][2][29],
F_[5][0][29],
F_[5][1][29],
F_[5][2][29],
F_[6][0][29],
F_[6][1][29],
F_[6][2][29],
F_[7][0][29],
F_[7][1][29],
F_[7][2][29],
F_[8][0][29],
F_[8][1][29],
F_[8][2][29],
F_[9][0][29],
F_[9][1][29],
F_[9][2][29],
F_[10][0][29],
F_[10][1][29],
F_[10][2][29],
F_[11][0][29],
F_[11][1][29],
F_[11][2][29],
F_[12][0][29],
F_[12][1][29],
F_[12][2][29],
F_[13][0][29],
F_[13][1][29],
F_[13][2][29],
F_[14][0][29],
F_[14][1][29],
F_[14][2][29],
F_[15][0][29],
F_[15][1][29],
F_[15][2][29],
F_[0][0][30],
F_[0][1][30],
F_[0][2][30],
F_[1][0][30],
F_[1][1][30],
F_[1][2][30],
F_[2][0][30],
F_[2][1][30],
F_[2][2][30],
F_[3][0][30],
F_[3][1][30],
F_[3][2][30],
F_[4][0][30],
F_[4][1][30],
F_[4][2][30],
F_[5][0][30],
F_[5][1][30],
F_[5][2][30],
F_[6][0][30],
F_[6][1][30],
F_[6][2][30],
F_[7][0][30],
F_[7][1][30],
F_[7][2][30],
F_[8][0][30],
F_[8][1][30],
F_[8][2][30],
F_[9][0][30],
F_[9][1][30],
F_[9][2][30],
F_[10][0][30],
F_[10][1][30],
F_[10][2][30],
F_[11][0][30],
F_[11][1][30],
F_[11][2][30],
F_[12][0][30],
F_[12][1][30],
F_[12][2][30],
F_[13][0][30],
F_[13][1][30],
F_[13][2][30],
F_[14][0][30],
F_[14][1][30],
F_[14][2][30],
F_[15][0][30],
F_[15][1][30],
F_[15][2][30],
F_[0][0][31],
F_[0][1][31],
F_[0][2][31],
F_[1][0][31],
F_[1][1][31],
F_[1][2][31],
F_[2][0][31],
F_[2][1][31],
F_[2][2][31],
F_[3][0][31],
F_[3][1][31],
F_[3][2][31],
F_[4][0][31],
F_[4][1][31],
F_[4][2][31],
F_[5][0][31],
F_[5][1][31],
F_[5][2][31],
F_[6][0][31],
F_[6][1][31],
F_[6][2][31],
F_[7][0][31],
F_[7][1][31],
F_[7][2][31],
F_[8][0][31],
F_[8][1][31],
F_[8][2][31],
F_[9][0][31],
F_[9][1][31],
F_[9][2][31],
F_[10][0][31],
F_[10][1][31],
F_[10][2][31],
F_[11][0][31],
F_[11][1][31],
F_[11][2][31],
F_[12][0][31],
F_[12][1][31],
F_[12][2][31],
F_[13][0][31],
F_[13][1][31],
F_[13][2][31],
F_[14][0][31],
F_[14][1][31],
F_[14][2][31],
F_[15][0][31],
F_[15][1][31],
F_[15][2][31],
F_[0][0][32],
F_[0][1][32],
F_[0][2][32],
F_[1][0][32],
F_[1][1][32],
F_[1][2][32],
F_[2][0][32],
F_[2][1][32],
F_[2][2][32],
F_[3][0][32],
F_[3][1][32],
F_[3][2][32],
F_[4][0][32],
F_[4][1][32],
F_[4][2][32],
F_[5][0][32],
F_[5][1][32],
F_[5][2][32],
F_[6][0][32],
F_[6][1][32],
F_[6][2][32],
F_[7][0][32],
F_[7][1][32],
F_[7][2][32],
F_[8][0][32],
F_[8][1][32],
F_[8][2][32],
F_[9][0][32],
F_[9][1][32],
F_[9][2][32],
F_[10][0][32],
F_[10][1][32],
F_[10][2][32],
F_[11][0][32],
F_[11][1][32],
F_[11][2][32],
F_[12][0][32],
F_[12][1][32],
F_[12][2][32],
F_[13][0][32],
F_[13][1][32],
F_[13][2][32],
F_[14][0][32],
F_[14][1][32],
F_[14][2][32],
F_[15][0][32],
F_[15][1][32],
F_[15][2][32],
F_[0][0][33],
F_[0][1][33],
F_[0][2][33],
F_[1][0][33],
F_[1][1][33],
F_[1][2][33],
F_[2][0][33],
F_[2][1][33],
F_[2][2][33],
F_[3][0][33],
F_[3][1][33],
F_[3][2][33],
F_[4][0][33],
F_[4][1][33],
F_[4][2][33],
F_[5][0][33],
F_[5][1][33],
F_[5][2][33],
F_[6][0][33],
F_[6][1][33],
F_[6][2][33],
F_[7][0][33],
F_[7][1][33],
F_[7][2][33],
F_[8][0][33],
F_[8][1][33],
F_[8][2][33],
F_[9][0][33],
F_[9][1][33],
F_[9][2][33],
F_[10][0][33],
F_[10][1][33],
F_[10][2][33],
F_[11][0][33],
F_[11][1][33],
F_[11][2][33],
F_[12][0][33],
F_[12][1][33],
F_[12][2][33],
F_[13][0][33],
F_[13][1][33],
F_[13][2][33],
F_[14][0][33],
F_[14][1][33],
F_[14][2][33],
F_[15][0][33],
F_[15][1][33],
F_[15][2][33],
F_[0][0][34],
F_[0][1][34],
F_[0][2][34],
F_[1][0][34],
F_[1][1][34],
F_[1][2][34],
F_[2][0][34],
F_[2][1][34],
F_[2][2][34],
F_[3][0][34],
F_[3][1][34],
F_[3][2][34],
F_[4][0][34],
F_[4][1][34],
F_[4][2][34],
F_[5][0][34],
F_[5][1][34],
F_[5][2][34],
F_[6][0][34],
F_[6][1][34],
F_[6][2][34],
F_[7][0][34],
F_[7][1][34],
F_[7][2][34],
F_[8][0][34],
F_[8][1][34],
F_[8][2][34],
F_[9][0][34],
F_[9][1][34],
F_[9][2][34],
F_[10][0][34],
F_[10][1][34],
F_[10][2][34],
F_[11][0][34],
F_[11][1][34],
F_[11][2][34],
F_[12][0][34],
F_[12][1][34],
F_[12][2][34],
F_[13][0][34],
F_[13][1][34],
F_[13][2][34],
F_[14][0][34],
F_[14][1][34],
F_[14][2][34],
F_[15][0][34],
F_[15][1][34],
F_[15][2][34],
F_[0][0][35],
F_[0][1][35],
F_[0][2][35],
F_[1][0][35],
F_[1][1][35],
F_[1][2][35],
F_[2][0][35],
F_[2][1][35],
F_[2][2][35],
F_[3][0][35],
F_[3][1][35],
F_[3][2][35],
F_[4][0][35],
F_[4][1][35],
F_[4][2][35],
F_[5][0][35],
F_[5][1][35],
F_[5][2][35],
F_[6][0][35],
F_[6][1][35],
F_[6][2][35],
F_[7][0][35],
F_[7][1][35],
F_[7][2][35],
F_[8][0][35],
F_[8][1][35],
F_[8][2][35],
F_[9][0][35],
F_[9][1][35],
F_[9][2][35],
F_[10][0][35],
F_[10][1][35],
F_[10][2][35],
F_[11][0][35],
F_[11][1][35],
F_[11][2][35],
F_[12][0][35],
F_[12][1][35],
F_[12][2][35],
F_[13][0][35],
F_[13][1][35],
F_[13][2][35],
F_[14][0][35],
F_[14][1][35],
F_[14][2][35],
F_[15][0][35],
F_[15][1][35],
F_[15][2][35],
F_[0][0][36],
F_[0][1][36],
F_[0][2][36],
F_[1][0][36],
F_[1][1][36],
F_[1][2][36],
F_[2][0][36],
F_[2][1][36],
F_[2][2][36],
F_[3][0][36],
F_[3][1][36],
F_[3][2][36],
F_[4][0][36],
F_[4][1][36],
F_[4][2][36],
F_[5][0][36],
F_[5][1][36],
F_[5][2][36],
F_[6][0][36],
F_[6][1][36],
F_[6][2][36],
F_[7][0][36],
F_[7][1][36],
F_[7][2][36],
F_[8][0][36],
F_[8][1][36],
F_[8][2][36],
F_[9][0][36],
F_[9][1][36],
F_[9][2][36],
F_[10][0][36],
F_[10][1][36],
F_[10][2][36],
F_[11][0][36],
F_[11][1][36],
F_[11][2][36],
F_[12][0][36],
F_[12][1][36],
F_[12][2][36],
F_[13][0][36],
F_[13][1][36],
F_[13][2][36],
F_[14][0][36],
F_[14][1][36],
F_[14][2][36],
F_[15][0][36],
F_[15][1][36],
F_[15][2][36],
F_[0][0][37],
F_[0][1][37],
F_[0][2][37],
F_[1][0][37],
F_[1][1][37],
F_[1][2][37],
F_[2][0][37],
F_[2][1][37],
F_[2][2][37],
F_[3][0][37],
F_[3][1][37],
F_[3][2][37],
F_[4][0][37],
F_[4][1][37],
F_[4][2][37],
F_[5][0][37],
F_[5][1][37],
F_[5][2][37],
F_[6][0][37],
F_[6][1][37],
F_[6][2][37],
F_[7][0][37],
F_[7][1][37],
F_[7][2][37],
F_[8][0][37],
F_[8][1][37],
F_[8][2][37],
F_[9][0][37],
F_[9][1][37],
F_[9][2][37],
F_[10][0][37],
F_[10][1][37],
F_[10][2][37],
F_[11][0][37],
F_[11][1][37],
F_[11][2][37],
F_[12][0][37],
F_[12][1][37],
F_[12][2][37],
F_[13][0][37],
F_[13][1][37],
F_[13][2][37],
F_[14][0][37],
F_[14][1][37],
F_[14][2][37],
F_[15][0][37],
F_[15][1][37],
F_[15][2][37],
F_[0][0][38],
F_[0][1][38],
F_[0][2][38],
F_[1][0][38],
F_[1][1][38],
F_[1][2][38],
F_[2][0][38],
F_[2][1][38],
F_[2][2][38],
F_[3][0][38],
F_[3][1][38],
F_[3][2][38],
F_[4][0][38],
F_[4][1][38],
F_[4][2][38],
F_[5][0][38],
F_[5][1][38],
F_[5][2][38],
F_[6][0][38],
F_[6][1][38],
F_[6][2][38],
F_[7][0][38],
F_[7][1][38],
F_[7][2][38],
F_[8][0][38],
F_[8][1][38],
F_[8][2][38],
F_[9][0][38],
F_[9][1][38],
F_[9][2][38],
F_[10][0][38],
F_[10][1][38],
F_[10][2][38],
F_[11][0][38],
F_[11][1][38],
F_[11][2][38],
F_[12][0][38],
F_[12][1][38],
F_[12][2][38],
F_[13][0][38],
F_[13][1][38],
F_[13][2][38],
F_[14][0][38],
F_[14][1][38],
F_[14][2][38],
F_[15][0][38],
F_[15][1][38],
F_[15][2][38],
F_[0][0][39],
F_[0][1][39],
F_[0][2][39],
F_[1][0][39],
F_[1][1][39],
F_[1][2][39],
F_[2][0][39],
F_[2][1][39],
F_[2][2][39],
F_[3][0][39],
F_[3][1][39],
F_[3][2][39],
F_[4][0][39],
F_[4][1][39],
F_[4][2][39],
F_[5][0][39],
F_[5][1][39],
F_[5][2][39],
F_[6][0][39],
F_[6][1][39],
F_[6][2][39],
F_[7][0][39],
F_[7][1][39],
F_[7][2][39],
F_[8][0][39],
F_[8][1][39],
F_[8][2][39],
F_[9][0][39],
F_[9][1][39],
F_[9][2][39],
F_[10][0][39],
F_[10][1][39],
F_[10][2][39],
F_[11][0][39],
F_[11][1][39],
F_[11][2][39],
F_[12][0][39],
F_[12][1][39],
F_[12][2][39],
F_[13][0][39],
F_[13][1][39],
F_[13][2][39],
F_[14][0][39],
F_[14][1][39],
F_[14][2][39],
F_[15][0][39],
F_[15][1][39],
F_[15][2][39],
F_[0][0][40],
F_[0][1][40],
F_[0][2][40],
F_[1][0][40],
F_[1][1][40],
F_[1][2][40],
F_[2][0][40],
F_[2][1][40],
F_[2][2][40],
F_[3][0][40],
F_[3][1][40],
F_[3][2][40],
F_[4][0][40],
F_[4][1][40],
F_[4][2][40],
F_[5][0][40],
F_[5][1][40],
F_[5][2][40],
F_[6][0][40],
F_[6][1][40],
F_[6][2][40],
F_[7][0][40],
F_[7][1][40],
F_[7][2][40],
F_[8][0][40],
F_[8][1][40],
F_[8][2][40],
F_[9][0][40],
F_[9][1][40],
F_[9][2][40],
F_[10][0][40],
F_[10][1][40],
F_[10][2][40],
F_[11][0][40],
F_[11][1][40],
F_[11][2][40],
F_[12][0][40],
F_[12][1][40],
F_[12][2][40],
F_[13][0][40],
F_[13][1][40],
F_[13][2][40],
F_[14][0][40],
F_[14][1][40],
F_[14][2][40],
F_[15][0][40],
F_[15][1][40],
F_[15][2][40],
F_[0][0][41],
F_[0][1][41],
F_[0][2][41],
F_[1][0][41],
F_[1][1][41],
F_[1][2][41],
F_[2][0][41],
F_[2][1][41],
F_[2][2][41],
F_[3][0][41],
F_[3][1][41],
F_[3][2][41],
F_[4][0][41],
F_[4][1][41],
F_[4][2][41],
F_[5][0][41],
F_[5][1][41],
F_[5][2][41],
F_[6][0][41],
F_[6][1][41],
F_[6][2][41],
F_[7][0][41],
F_[7][1][41],
F_[7][2][41],
F_[8][0][41],
F_[8][1][41],
F_[8][2][41],
F_[9][0][41],
F_[9][1][41],
F_[9][2][41],
F_[10][0][41],
F_[10][1][41],
F_[10][2][41],
F_[11][0][41],
F_[11][1][41],
F_[11][2][41],
F_[12][0][41],
F_[12][1][41],
F_[12][2][41],
F_[13][0][41],
F_[13][1][41],
F_[13][2][41],
F_[14][0][41],
F_[14][1][41],
F_[14][2][41],
F_[15][0][41],
F_[15][1][41],
F_[15][2][41],
F_[0][0][42],
F_[0][1][42],
F_[0][2][42],
F_[1][0][42],
F_[1][1][42],
F_[1][2][42],
F_[2][0][42],
F_[2][1][42],
F_[2][2][42],
F_[3][0][42],
F_[3][1][42],
F_[3][2][42],
F_[4][0][42],
F_[4][1][42],
F_[4][2][42],
F_[5][0][42],
F_[5][1][42],
F_[5][2][42],
F_[6][0][42],
F_[6][1][42],
F_[6][2][42],
F_[7][0][42],
F_[7][1][42],
F_[7][2][42],
F_[8][0][42],
F_[8][1][42],
F_[8][2][42],
F_[9][0][42],
F_[9][1][42],
F_[9][2][42],
F_[10][0][42],
F_[10][1][42],
F_[10][2][42],
F_[11][0][42],
F_[11][1][42],
F_[11][2][42],
F_[12][0][42],
F_[12][1][42],
F_[12][2][42],
F_[13][0][42],
F_[13][1][42],
F_[13][2][42],
F_[14][0][42],
F_[14][1][42],
F_[14][2][42],
F_[15][0][42],
F_[15][1][42],
F_[15][2][42],
F_[0][0][43],
F_[0][1][43],
F_[0][2][43],
F_[1][0][43],
F_[1][1][43],
F_[1][2][43],
F_[2][0][43],
F_[2][1][43],
F_[2][2][43],
F_[3][0][43],
F_[3][1][43],
F_[3][2][43],
F_[4][0][43],
F_[4][1][43],
F_[4][2][43],
F_[5][0][43],
F_[5][1][43],
F_[5][2][43],
F_[6][0][43],
F_[6][1][43],
F_[6][2][43],
F_[7][0][43],
F_[7][1][43],
F_[7][2][43],
F_[8][0][43],
F_[8][1][43],
F_[8][2][43],
F_[9][0][43],
F_[9][1][43],
F_[9][2][43],
F_[10][0][43],
F_[10][1][43],
F_[10][2][43],
F_[11][0][43],
F_[11][1][43],
F_[11][2][43],
F_[12][0][43],
F_[12][1][43],
F_[12][2][43],
F_[13][0][43],
F_[13][1][43],
F_[13][2][43],
F_[14][0][43],
F_[14][1][43],
F_[14][2][43],
F_[15][0][43],
F_[15][1][43],
F_[15][2][43],
F_[0][0][44],
F_[0][1][44],
F_[0][2][44],
F_[1][0][44],
F_[1][1][44],
F_[1][2][44],
F_[2][0][44],
F_[2][1][44],
F_[2][2][44],
F_[3][0][44],
F_[3][1][44],
F_[3][2][44],
F_[4][0][44],
F_[4][1][44],
F_[4][2][44],
F_[5][0][44],
F_[5][1][44],
F_[5][2][44],
F_[6][0][44],
F_[6][1][44],
F_[6][2][44],
F_[7][0][44],
F_[7][1][44],
F_[7][2][44],
F_[8][0][44],
F_[8][1][44],
F_[8][2][44],
F_[9][0][44],
F_[9][1][44],
F_[9][2][44],
F_[10][0][44],
F_[10][1][44],
F_[10][2][44],
F_[11][0][44],
F_[11][1][44],
F_[11][2][44],
F_[12][0][44],
F_[12][1][44],
F_[12][2][44],
F_[13][0][44],
F_[13][1][44],
F_[13][2][44],
F_[14][0][44],
F_[14][1][44],
F_[14][2][44],
F_[15][0][44],
F_[15][1][44],
F_[15][2][44],
F_[0][0][45],
F_[0][1][45],
F_[0][2][45],
F_[1][0][45],
F_[1][1][45],
F_[1][2][45],
F_[2][0][45],
F_[2][1][45],
F_[2][2][45],
F_[3][0][45],
F_[3][1][45],
F_[3][2][45],
F_[4][0][45],
F_[4][1][45],
F_[4][2][45],
F_[5][0][45],
F_[5][1][45],
F_[5][2][45],
F_[6][0][45],
F_[6][1][45],
F_[6][2][45],
F_[7][0][45],
F_[7][1][45],
F_[7][2][45],
F_[8][0][45],
F_[8][1][45],
F_[8][2][45],
F_[9][0][45],
F_[9][1][45],
F_[9][2][45],
F_[10][0][45],
F_[10][1][45],
F_[10][2][45],
F_[11][0][45],
F_[11][1][45],
F_[11][2][45],
F_[12][0][45],
F_[12][1][45],
F_[12][2][45],
F_[13][0][45],
F_[13][1][45],
F_[13][2][45],
F_[14][0][45],
F_[14][1][45],
F_[14][2][45],
F_[15][0][45],
F_[15][1][45],
F_[15][2][45],
F_[0][0][46],
F_[0][1][46],
F_[0][2][46],
F_[1][0][46],
F_[1][1][46],
F_[1][2][46],
F_[2][0][46],
F_[2][1][46],
F_[2][2][46],
F_[3][0][46],
F_[3][1][46],
F_[3][2][46],
F_[4][0][46],
F_[4][1][46],
F_[4][2][46],
F_[5][0][46],
F_[5][1][46],
F_[5][2][46],
F_[6][0][46],
F_[6][1][46],
F_[6][2][46],
F_[7][0][46],
F_[7][1][46],
F_[7][2][46],
F_[8][0][46],
F_[8][1][46],
F_[8][2][46],
F_[9][0][46],
F_[9][1][46],
F_[9][2][46],
F_[10][0][46],
F_[10][1][46],
F_[10][2][46],
F_[11][0][46],
F_[11][1][46],
F_[11][2][46],
F_[12][0][46],
F_[12][1][46],
F_[12][2][46],
F_[13][0][46],
F_[13][1][46],
F_[13][2][46],
F_[14][0][46],
F_[14][1][46],
F_[14][2][46],
F_[15][0][46],
F_[15][1][46],
F_[15][2][46],
F_[0][0][47],
F_[0][1][47],
F_[0][2][47],
F_[1][0][47],
F_[1][1][47],
F_[1][2][47],
F_[2][0][47],
F_[2][1][47],
F_[2][2][47],
F_[3][0][47],
F_[3][1][47],
F_[3][2][47],
F_[4][0][47],
F_[4][1][47],
F_[4][2][47],
F_[5][0][47],
F_[5][1][47],
F_[5][2][47],
F_[6][0][47],
F_[6][1][47],
F_[6][2][47],
F_[7][0][47],
F_[7][1][47],
F_[7][2][47],
F_[8][0][47],
F_[8][1][47],
F_[8][2][47],
F_[9][0][47],
F_[9][1][47],
F_[9][2][47],
F_[10][0][47],
F_[10][1][47],
F_[10][2][47],
F_[11][0][47],
F_[11][1][47],
F_[11][2][47],
F_[12][0][47],
F_[12][1][47],
F_[12][2][47],
F_[13][0][47],
F_[13][1][47],
F_[13][2][47],
F_[14][0][47],
F_[14][1][47],
F_[14][2][47],
F_[15][0][47],
F_[15][1][47],
F_[15][2][47],
F_[0][0][48],
F_[0][1][48],
F_[0][2][48],
F_[1][0][48],
F_[1][1][48],
F_[1][2][48],
F_[2][0][48],
F_[2][1][48],
F_[2][2][48],
F_[3][0][48],
F_[3][1][48],
F_[3][2][48],
F_[4][0][48],
F_[4][1][48],
F_[4][2][48],
F_[5][0][48],
F_[5][1][48],
F_[5][2][48],
F_[6][0][48],
F_[6][1][48],
F_[6][2][48],
F_[7][0][48],
F_[7][1][48],
F_[7][2][48],
F_[8][0][48],
F_[8][1][48],
F_[8][2][48],
F_[9][0][48],
F_[9][1][48],
F_[9][2][48],
F_[10][0][48],
F_[10][1][48],
F_[10][2][48],
F_[11][0][48],
F_[11][1][48],
F_[11][2][48],
F_[12][0][48],
F_[12][1][48],
F_[12][2][48],
F_[13][0][48],
F_[13][1][48],
F_[13][2][48],
F_[14][0][48],
F_[14][1][48],
F_[14][2][48],
F_[15][0][48],
F_[15][1][48],
F_[15][2][48],
F_[0][0][49],
F_[0][1][49],
F_[0][2][49],
F_[1][0][49],
F_[1][1][49],
F_[1][2][49],
F_[2][0][49],
F_[2][1][49],
F_[2][2][49],
F_[3][0][49],
F_[3][1][49],
F_[3][2][49],
F_[4][0][49],
F_[4][1][49],
F_[4][2][49],
F_[5][0][49],
F_[5][1][49],
F_[5][2][49],
F_[6][0][49],
F_[6][1][49],
F_[6][2][49],
F_[7][0][49],
F_[7][1][49],
F_[7][2][49],
F_[8][0][49],
F_[8][1][49],
F_[8][2][49],
F_[9][0][49],
F_[9][1][49],
F_[9][2][49],
F_[10][0][49],
F_[10][1][49],
F_[10][2][49],
F_[11][0][49],
F_[11][1][49],
F_[11][2][49],
F_[12][0][49],
F_[12][1][49],
F_[12][2][49],
F_[13][0][49],
F_[13][1][49],
F_[13][2][49],
F_[14][0][49],
F_[14][1][49],
F_[14][2][49],
F_[15][0][49],
F_[15][1][49],
F_[15][2][49],
F_[0][0][50],
F_[0][1][50],
F_[0][2][50],
F_[1][0][50],
F_[1][1][50],
F_[1][2][50],
F_[2][0][50],
F_[2][1][50],
F_[2][2][50],
F_[3][0][50],
F_[3][1][50],
F_[3][2][50],
F_[4][0][50],
F_[4][1][50],
F_[4][2][50],
F_[5][0][50],
F_[5][1][50],
F_[5][2][50],
F_[6][0][50],
F_[6][1][50],
F_[6][2][50],
F_[7][0][50],
F_[7][1][50],
F_[7][2][50],
F_[8][0][50],
F_[8][1][50],
F_[8][2][50],
F_[9][0][50],
F_[9][1][50],
F_[9][2][50],
F_[10][0][50],
F_[10][1][50],
F_[10][2][50],
F_[11][0][50],
F_[11][1][50],
F_[11][2][50],
F_[12][0][50],
F_[12][1][50],
F_[12][2][50],
F_[13][0][50],
F_[13][1][50],
F_[13][2][50],
F_[14][0][50],
F_[14][1][50],
F_[14][2][50],
F_[15][0][50],
F_[15][1][50],
F_[15][2][50],
F_[0][0][51],
F_[0][1][51],
F_[0][2][51],
F_[1][0][51],
F_[1][1][51],
F_[1][2][51],
F_[2][0][51],
F_[2][1][51],
F_[2][2][51],
F_[3][0][51],
F_[3][1][51],
F_[3][2][51],
F_[4][0][51],
F_[4][1][51],
F_[4][2][51],
F_[5][0][51],
F_[5][1][51],
F_[5][2][51],
F_[6][0][51],
F_[6][1][51],
F_[6][2][51],
F_[7][0][51],
F_[7][1][51],
F_[7][2][51],
F_[8][0][51],
F_[8][1][51],
F_[8][2][51],
F_[9][0][51],
F_[9][1][51],
F_[9][2][51],
F_[10][0][51],
F_[10][1][51],
F_[10][2][51],
F_[11][0][51],
F_[11][1][51],
F_[11][2][51],
F_[12][0][51],
F_[12][1][51],
F_[12][2][51],
F_[13][0][51],
F_[13][1][51],
F_[13][2][51],
F_[14][0][51],
F_[14][1][51],
F_[14][2][51],
F_[15][0][51],
F_[15][1][51],
F_[15][2][51],
F_[0][0][52],
F_[0][1][52],
F_[0][2][52],
F_[1][0][52],
F_[1][1][52],
F_[1][2][52],
F_[2][0][52],
F_[2][1][52],
F_[2][2][52],
F_[3][0][52],
F_[3][1][52],
F_[3][2][52],
F_[4][0][52],
F_[4][1][52],
F_[4][2][52],
F_[5][0][52],
F_[5][1][52],
F_[5][2][52],
F_[6][0][52],
F_[6][1][52],
F_[6][2][52],
F_[7][0][52],
F_[7][1][52],
F_[7][2][52],
F_[8][0][52],
F_[8][1][52],
F_[8][2][52],
F_[9][0][52],
F_[9][1][52],
F_[9][2][52],
F_[10][0][52],
F_[10][1][52],
F_[10][2][52],
F_[11][0][52],
F_[11][1][52],
F_[11][2][52],
F_[12][0][52],
F_[12][1][52],
F_[12][2][52],
F_[13][0][52],
F_[13][1][52],
F_[13][2][52],
F_[14][0][52],
F_[14][1][52],
F_[14][2][52],
F_[15][0][52],
F_[15][1][52],
F_[15][2][52],
F_[0][0][53],
F_[0][1][53],
F_[0][2][53],
F_[1][0][53],
F_[1][1][53],
F_[1][2][53],
F_[2][0][53],
F_[2][1][53],
F_[2][2][53],
F_[3][0][53],
F_[3][1][53],
F_[3][2][53],
F_[4][0][53],
F_[4][1][53],
F_[4][2][53],
F_[5][0][53],
F_[5][1][53],
F_[5][2][53],
F_[6][0][53],
F_[6][1][53],
F_[6][2][53],
F_[7][0][53],
F_[7][1][53],
F_[7][2][53],
F_[8][0][53],
F_[8][1][53],
F_[8][2][53],
F_[9][0][53],
F_[9][1][53],
F_[9][2][53],
F_[10][0][53],
F_[10][1][53],
F_[10][2][53],
F_[11][0][53],
F_[11][1][53],
F_[11][2][53],
F_[12][0][53],
F_[12][1][53],
F_[12][2][53],
F_[13][0][53],
F_[13][1][53],
F_[13][2][53],
F_[14][0][53],
F_[14][1][53],
F_[14][2][53],
F_[15][0][53],
F_[15][1][53],
F_[15][2][53],
F_[0][0][54],
F_[0][1][54],
F_[0][2][54],
F_[1][0][54],
F_[1][1][54],
F_[1][2][54],
F_[2][0][54],
F_[2][1][54],
F_[2][2][54],
F_[3][0][54],
F_[3][1][54],
F_[3][2][54],
F_[4][0][54],
F_[4][1][54],
F_[4][2][54],
F_[5][0][54],
F_[5][1][54],
F_[5][2][54],
F_[6][0][54],
F_[6][1][54],
F_[6][2][54],
F_[7][0][54],
F_[7][1][54],
F_[7][2][54],
F_[8][0][54],
F_[8][1][54],
F_[8][2][54],
F_[9][0][54],
F_[9][1][54],
F_[9][2][54],
F_[10][0][54],
F_[10][1][54],
F_[10][2][54],
F_[11][0][54],
F_[11][1][54],
F_[11][2][54],
F_[12][0][54],
F_[12][1][54],
F_[12][2][54],
F_[13][0][54],
F_[13][1][54],
F_[13][2][54],
F_[14][0][54],
F_[14][1][54],
F_[14][2][54],
F_[15][0][54],
F_[15][1][54],
F_[15][2][54],
F_[0][0][55],
F_[0][1][55],
F_[0][2][55],
F_[1][0][55],
F_[1][1][55],
F_[1][2][55],
F_[2][0][55],
F_[2][1][55],
F_[2][2][55],
F_[3][0][55],
F_[3][1][55],
F_[3][2][55],
F_[4][0][55],
F_[4][1][55],
F_[4][2][55],
F_[5][0][55],
F_[5][1][55],
F_[5][2][55],
F_[6][0][55],
F_[6][1][55],
F_[6][2][55],
F_[7][0][55],
F_[7][1][55],
F_[7][2][55],
F_[8][0][55],
F_[8][1][55],
F_[8][2][55],
F_[9][0][55],
F_[9][1][55],
F_[9][2][55],
F_[10][0][55],
F_[10][1][55],
F_[10][2][55],
F_[11][0][55],
F_[11][1][55],
F_[11][2][55],
F_[12][0][55],
F_[12][1][55],
F_[12][2][55],
F_[13][0][55],
F_[13][1][55],
F_[13][2][55],
F_[14][0][55],
F_[14][1][55],
F_[14][2][55],
F_[15][0][55],
F_[15][1][55],
F_[15][2][55],
F_[0][0][56],
F_[0][1][56],
F_[0][2][56],
F_[1][0][56],
F_[1][1][56],
F_[1][2][56],
F_[2][0][56],
F_[2][1][56],
F_[2][2][56],
F_[3][0][56],
F_[3][1][56],
F_[3][2][56],
F_[4][0][56],
F_[4][1][56],
F_[4][2][56],
F_[5][0][56],
F_[5][1][56],
F_[5][2][56],
F_[6][0][56],
F_[6][1][56],
F_[6][2][56],
F_[7][0][56],
F_[7][1][56],
F_[7][2][56],
F_[8][0][56],
F_[8][1][56],
F_[8][2][56],
F_[9][0][56],
F_[9][1][56],
F_[9][2][56],
F_[10][0][56],
F_[10][1][56],
F_[10][2][56],
F_[11][0][56],
F_[11][1][56],
F_[11][2][56],
F_[12][0][56],
F_[12][1][56],
F_[12][2][56],
F_[13][0][56],
F_[13][1][56],
F_[13][2][56],
F_[14][0][56],
F_[14][1][56],
F_[14][2][56],
F_[15][0][56],
F_[15][1][56],
F_[15][2][56],
F_[0][0][57],
F_[0][1][57],
F_[0][2][57],
F_[1][0][57],
F_[1][1][57],
F_[1][2][57],
F_[2][0][57],
F_[2][1][57],
F_[2][2][57],
F_[3][0][57],
F_[3][1][57],
F_[3][2][57],
F_[4][0][57],
F_[4][1][57],
F_[4][2][57],
F_[5][0][57],
F_[5][1][57],
F_[5][2][57],
F_[6][0][57],
F_[6][1][57],
F_[6][2][57],
F_[7][0][57],
F_[7][1][57],
F_[7][2][57],
F_[8][0][57],
F_[8][1][57],
F_[8][2][57],
F_[9][0][57],
F_[9][1][57],
F_[9][2][57],
F_[10][0][57],
F_[10][1][57],
F_[10][2][57],
F_[11][0][57],
F_[11][1][57],
F_[11][2][57],
F_[12][0][57],
F_[12][1][57],
F_[12][2][57],
F_[13][0][57],
F_[13][1][57],
F_[13][2][57],
F_[14][0][57],
F_[14][1][57],
F_[14][2][57],
F_[15][0][57],
F_[15][1][57],
F_[15][2][57],
F_[0][0][58],
F_[0][1][58],
F_[0][2][58],
F_[1][0][58],
F_[1][1][58],
F_[1][2][58],
F_[2][0][58],
F_[2][1][58],
F_[2][2][58],
F_[3][0][58],
F_[3][1][58],
F_[3][2][58],
F_[4][0][58],
F_[4][1][58],
F_[4][2][58],
F_[5][0][58],
F_[5][1][58],
F_[5][2][58],
F_[6][0][58],
F_[6][1][58],
F_[6][2][58],
F_[7][0][58],
F_[7][1][58],
F_[7][2][58],
F_[8][0][58],
F_[8][1][58],
F_[8][2][58],
F_[9][0][58],
F_[9][1][58],
F_[9][2][58],
F_[10][0][58],
F_[10][1][58],
F_[10][2][58],
F_[11][0][58],
F_[11][1][58],
F_[11][2][58],
F_[12][0][58],
F_[12][1][58],
F_[12][2][58],
F_[13][0][58],
F_[13][1][58],
F_[13][2][58],
F_[14][0][58],
F_[14][1][58],
F_[14][2][58],
F_[15][0][58],
F_[15][1][58],
F_[15][2][58],
F_[0][0][59],
F_[0][1][59],
F_[0][2][59],
F_[1][0][59],
F_[1][1][59],
F_[1][2][59],
F_[2][0][59],
F_[2][1][59],
F_[2][2][59],
F_[3][0][59],
F_[3][1][59],
F_[3][2][59],
F_[4][0][59],
F_[4][1][59],
F_[4][2][59],
F_[5][0][59],
F_[5][1][59],
F_[5][2][59],
F_[6][0][59],
F_[6][1][59],
F_[6][2][59],
F_[7][0][59],
F_[7][1][59],
F_[7][2][59],
F_[8][0][59],
F_[8][1][59],
F_[8][2][59],
F_[9][0][59],
F_[9][1][59],
F_[9][2][59],
F_[10][0][59],
F_[10][1][59],
F_[10][2][59],
F_[11][0][59],
F_[11][1][59],
F_[11][2][59],
F_[12][0][59],
F_[12][1][59],
F_[12][2][59],
F_[13][0][59],
F_[13][1][59],
F_[13][2][59],
F_[14][0][59],
F_[14][1][59],
F_[14][2][59],
F_[15][0][59],
F_[15][1][59],
F_[15][2][59],
F_[0][0][60],
F_[0][1][60],
F_[0][2][60],
F_[1][0][60],
F_[1][1][60],
F_[1][2][60],
F_[2][0][60],
F_[2][1][60],
F_[2][2][60],
F_[3][0][60],
F_[3][1][60],
F_[3][2][60],
F_[4][0][60],
F_[4][1][60],
F_[4][2][60],
F_[5][0][60],
F_[5][1][60],
F_[5][2][60],
F_[6][0][60],
F_[6][1][60],
F_[6][2][60],
F_[7][0][60],
F_[7][1][60],
F_[7][2][60],
F_[8][0][60],
F_[8][1][60],
F_[8][2][60],
F_[9][0][60],
F_[9][1][60],
F_[9][2][60],
F_[10][0][60],
F_[10][1][60],
F_[10][2][60],
F_[11][0][60],
F_[11][1][60],
F_[11][2][60],
F_[12][0][60],
F_[12][1][60],
F_[12][2][60],
F_[13][0][60],
F_[13][1][60],
F_[13][2][60],
F_[14][0][60],
F_[14][1][60],
F_[14][2][60],
F_[15][0][60],
F_[15][1][60],
F_[15][2][60],
F_[0][0][61],
F_[0][1][61],
F_[0][2][61],
F_[1][0][61],
F_[1][1][61],
F_[1][2][61],
F_[2][0][61],
F_[2][1][61],
F_[2][2][61],
F_[3][0][61],
F_[3][1][61],
F_[3][2][61],
F_[4][0][61],
F_[4][1][61],
F_[4][2][61],
F_[5][0][61],
F_[5][1][61],
F_[5][2][61],
F_[6][0][61],
F_[6][1][61],
F_[6][2][61],
F_[7][0][61],
F_[7][1][61],
F_[7][2][61],
F_[8][0][61],
F_[8][1][61],
F_[8][2][61],
F_[9][0][61],
F_[9][1][61],
F_[9][2][61],
F_[10][0][61],
F_[10][1][61],
F_[10][2][61],
F_[11][0][61],
F_[11][1][61],
F_[11][2][61],
F_[12][0][61],
F_[12][1][61],
F_[12][2][61],
F_[13][0][61],
F_[13][1][61],
F_[13][2][61],
F_[14][0][61],
F_[14][1][61],
F_[14][2][61],
F_[15][0][61],
F_[15][1][61],
F_[15][2][61],
F_[0][0][62],
F_[0][1][62],
F_[0][2][62],
F_[1][0][62],
F_[1][1][62],
F_[1][2][62],
F_[2][0][62],
F_[2][1][62],
F_[2][2][62],
F_[3][0][62],
F_[3][1][62],
F_[3][2][62],
F_[4][0][62],
F_[4][1][62],
F_[4][2][62],
F_[5][0][62],
F_[5][1][62],
F_[5][2][62],
F_[6][0][62],
F_[6][1][62],
F_[6][2][62],
F_[7][0][62],
F_[7][1][62],
F_[7][2][62],
F_[8][0][62],
F_[8][1][62],
F_[8][2][62],
F_[9][0][62],
F_[9][1][62],
F_[9][2][62],
F_[10][0][62],
F_[10][1][62],
F_[10][2][62],
F_[11][0][62],
F_[11][1][62],
F_[11][2][62],
F_[12][0][62],
F_[12][1][62],
F_[12][2][62],
F_[13][0][62],
F_[13][1][62],
F_[13][2][62],
F_[14][0][62],
F_[14][1][62],
F_[14][2][62],
F_[15][0][62],
F_[15][1][62],
F_[15][2][62],
F_[0][0][63],
F_[0][1][63],
F_[0][2][63],
F_[1][0][63],
F_[1][1][63],
F_[1][2][63],
F_[2][0][63],
F_[2][1][63],
F_[2][2][63],
F_[3][0][63],
F_[3][1][63],
F_[3][2][63],
F_[4][0][63],
F_[4][1][63],
F_[4][2][63],
F_[5][0][63],
F_[5][1][63],
F_[5][2][63],
F_[6][0][63],
F_[6][1][63],
F_[6][2][63],
F_[7][0][63],
F_[7][1][63],
F_[7][2][63],
F_[8][0][63],
F_[8][1][63],
F_[8][2][63],
F_[9][0][63],
F_[9][1][63],
F_[9][2][63],
F_[10][0][63],
F_[10][1][63],
F_[10][2][63],
F_[11][0][63],
F_[11][1][63],
F_[11][2][63],
F_[12][0][63],
F_[12][1][63],
F_[12][2][63],
F_[13][0][63],
F_[13][1][63],
F_[13][2][63],
F_[14][0][63],
F_[14][1][63],
F_[14][2][63],
F_[15][0][63],
F_[15][1][63],
F_[15][2][63],
F_[0][0][64],
F_[0][1][64],
F_[0][2][64],
F_[1][0][64],
F_[1][1][64],
F_[1][2][64],
F_[2][0][64],
F_[2][1][64],
F_[2][2][64],
F_[3][0][64],
F_[3][1][64],
F_[3][2][64],
F_[4][0][64],
F_[4][1][64],
F_[4][2][64],
F_[5][0][64],
F_[5][1][64],
F_[5][2][64],
F_[6][0][64],
F_[6][1][64],
F_[6][2][64],
F_[7][0][64],
F_[7][1][64],
F_[7][2][64],
F_[8][0][64],
F_[8][1][64],
F_[8][2][64],
F_[9][0][64],
F_[9][1][64],
F_[9][2][64],
F_[10][0][64],
F_[10][1][64],
F_[10][2][64],
F_[11][0][64],
F_[11][1][64],
F_[11][2][64],
F_[12][0][64],
F_[12][1][64],
F_[12][2][64],
F_[13][0][64],
F_[13][1][64],
F_[13][2][64],
F_[14][0][64],
F_[14][1][64],
F_[14][2][64],
F_[15][0][64],
F_[15][1][64],
F_[15][2][64],
F_[0][0][65],
F_[0][1][65],
F_[0][2][65],
F_[1][0][65],
F_[1][1][65],
F_[1][2][65],
F_[2][0][65],
F_[2][1][65],
F_[2][2][65],
F_[3][0][65],
F_[3][1][65],
F_[3][2][65],
F_[4][0][65],
F_[4][1][65],
F_[4][2][65],
F_[5][0][65],
F_[5][1][65],
F_[5][2][65],
F_[6][0][65],
F_[6][1][65],
F_[6][2][65],
F_[7][0][65],
F_[7][1][65],
F_[7][2][65],
F_[8][0][65],
F_[8][1][65],
F_[8][2][65],
F_[9][0][65],
F_[9][1][65],
F_[9][2][65],
F_[10][0][65],
F_[10][1][65],
F_[10][2][65],
F_[11][0][65],
F_[11][1][65],
F_[11][2][65],
F_[12][0][65],
F_[12][1][65],
F_[12][2][65],
F_[13][0][65],
F_[13][1][65],
F_[13][2][65],
F_[14][0][65],
F_[14][1][65],
F_[14][2][65],
F_[15][0][65],
F_[15][1][65],
F_[15][2][65],
F_[0][0][66],
F_[0][1][66],
F_[0][2][66],
F_[1][0][66],
F_[1][1][66],
F_[1][2][66],
F_[2][0][66],
F_[2][1][66],
F_[2][2][66],
F_[3][0][66],
F_[3][1][66],
F_[3][2][66],
F_[4][0][66],
F_[4][1][66],
F_[4][2][66],
F_[5][0][66],
F_[5][1][66],
F_[5][2][66],
F_[6][0][66],
F_[6][1][66],
F_[6][2][66],
F_[7][0][66],
F_[7][1][66],
F_[7][2][66],
F_[8][0][66],
F_[8][1][66],
F_[8][2][66],
F_[9][0][66],
F_[9][1][66],
F_[9][2][66],
F_[10][0][66],
F_[10][1][66],
F_[10][2][66],
F_[11][0][66],
F_[11][1][66],
F_[11][2][66],
F_[12][0][66],
F_[12][1][66],
F_[12][2][66],
F_[13][0][66],
F_[13][1][66],
F_[13][2][66],
F_[14][0][66],
F_[14][1][66],
F_[14][2][66],
F_[15][0][66],
F_[15][1][66],
F_[15][2][66],
F_[0][0][67],
F_[0][1][67],
F_[0][2][67],
F_[1][0][67],
F_[1][1][67],
F_[1][2][67],
F_[2][0][67],
F_[2][1][67],
F_[2][2][67],
F_[3][0][67],
F_[3][1][67],
F_[3][2][67],
F_[4][0][67],
F_[4][1][67],
F_[4][2][67],
F_[5][0][67],
F_[5][1][67],
F_[5][2][67],
F_[6][0][67],
F_[6][1][67],
F_[6][2][67],
F_[7][0][67],
F_[7][1][67],
F_[7][2][67],
F_[8][0][67],
F_[8][1][67],
F_[8][2][67],
F_[9][0][67],
F_[9][1][67],
F_[9][2][67],
F_[10][0][67],
F_[10][1][67],
F_[10][2][67],
F_[11][0][67],
F_[11][1][67],
F_[11][2][67],
F_[12][0][67],
F_[12][1][67],
F_[12][2][67],
F_[13][0][67],
F_[13][1][67],
F_[13][2][67],
F_[14][0][67],
F_[14][1][67],
F_[14][2][67],
F_[15][0][67],
F_[15][1][67],
F_[15][2][67],
F_[0][0][68],
F_[0][1][68],
F_[0][2][68],
F_[1][0][68],
F_[1][1][68],
F_[1][2][68],
F_[2][0][68],
F_[2][1][68],
F_[2][2][68],
F_[3][0][68],
F_[3][1][68],
F_[3][2][68],
F_[4][0][68],
F_[4][1][68],
F_[4][2][68],
F_[5][0][68],
F_[5][1][68],
F_[5][2][68],
F_[6][0][68],
F_[6][1][68],
F_[6][2][68],
F_[7][0][68],
F_[7][1][68],
F_[7][2][68],
F_[8][0][68],
F_[8][1][68],
F_[8][2][68],
F_[9][0][68],
F_[9][1][68],
F_[9][2][68],
F_[10][0][68],
F_[10][1][68],
F_[10][2][68],
F_[11][0][68],
F_[11][1][68],
F_[11][2][68],
F_[12][0][68],
F_[12][1][68],
F_[12][2][68],
F_[13][0][68],
F_[13][1][68],
F_[13][2][68],
F_[14][0][68],
F_[14][1][68],
F_[14][2][68],
F_[15][0][68],
F_[15][1][68],
F_[15][2][68],
F_[0][0][69],
F_[0][1][69],
F_[0][2][69],
F_[1][0][69],
F_[1][1][69],
F_[1][2][69],
F_[2][0][69],
F_[2][1][69],
F_[2][2][69],
F_[3][0][69],
F_[3][1][69],
F_[3][2][69],
F_[4][0][69],
F_[4][1][69],
F_[4][2][69],
F_[5][0][69],
F_[5][1][69],
F_[5][2][69],
F_[6][0][69],
F_[6][1][69],
F_[6][2][69],
F_[7][0][69],
F_[7][1][69],
F_[7][2][69],
F_[8][0][69],
F_[8][1][69],
F_[8][2][69],
F_[9][0][69],
F_[9][1][69],
F_[9][2][69],
F_[10][0][69],
F_[10][1][69],
F_[10][2][69],
F_[11][0][69],
F_[11][1][69],
F_[11][2][69],
F_[12][0][69],
F_[12][1][69],
F_[12][2][69],
F_[13][0][69],
F_[13][1][69],
F_[13][2][69],
F_[14][0][69],
F_[14][1][69],
F_[14][2][69],
F_[15][0][69],
F_[15][1][69],
F_[15][2][69],
F_[0][0][70],
F_[0][1][70],
F_[0][2][70],
F_[1][0][70],
F_[1][1][70],
F_[1][2][70],
F_[2][0][70],
F_[2][1][70],
F_[2][2][70],
F_[3][0][70],
F_[3][1][70],
F_[3][2][70],
F_[4][0][70],
F_[4][1][70],
F_[4][2][70],
F_[5][0][70],
F_[5][1][70],
F_[5][2][70],
F_[6][0][70],
F_[6][1][70],
F_[6][2][70],
F_[7][0][70],
F_[7][1][70],
F_[7][2][70],
F_[8][0][70],
F_[8][1][70],
F_[8][2][70],
F_[9][0][70],
F_[9][1][70],
F_[9][2][70],
F_[10][0][70],
F_[10][1][70],
F_[10][2][70],
F_[11][0][70],
F_[11][1][70],
F_[11][2][70],
F_[12][0][70],
F_[12][1][70],
F_[12][2][70],
F_[13][0][70],
F_[13][1][70],
F_[13][2][70],
F_[14][0][70],
F_[14][1][70],
F_[14][2][70],
F_[15][0][70],
F_[15][1][70],
F_[15][2][70],
F_[0][0][71],
F_[0][1][71],
F_[0][2][71],
F_[1][0][71],
F_[1][1][71],
F_[1][2][71],
F_[2][0][71],
F_[2][1][71],
F_[2][2][71],
F_[3][0][71],
F_[3][1][71],
F_[3][2][71],
F_[4][0][71],
F_[4][1][71],
F_[4][2][71],
F_[5][0][71],
F_[5][1][71],
F_[5][2][71],
F_[6][0][71],
F_[6][1][71],
F_[6][2][71],
F_[7][0][71],
F_[7][1][71],
F_[7][2][71],
F_[8][0][71],
F_[8][1][71],
F_[8][2][71],
F_[9][0][71],
F_[9][1][71],
F_[9][2][71],
F_[10][0][71],
F_[10][1][71],
F_[10][2][71],
F_[11][0][71],
F_[11][1][71],
F_[11][2][71],
F_[12][0][71],
F_[12][1][71],
F_[12][2][71],
F_[13][0][71],
F_[13][1][71],
F_[13][2][71],
F_[14][0][71],
F_[14][1][71],
F_[14][2][71],
F_[15][0][71],
F_[15][1][71],
F_[15][2][71],
F_[0][0][72],
F_[0][1][72],
F_[0][2][72],
F_[1][0][72],
F_[1][1][72],
F_[1][2][72],
F_[2][0][72],
F_[2][1][72],
F_[2][2][72],
F_[3][0][72],
F_[3][1][72],
F_[3][2][72],
F_[4][0][72],
F_[4][1][72],
F_[4][2][72],
F_[5][0][72],
F_[5][1][72],
F_[5][2][72],
F_[6][0][72],
F_[6][1][72],
F_[6][2][72],
F_[7][0][72],
F_[7][1][72],
F_[7][2][72],
F_[8][0][72],
F_[8][1][72],
F_[8][2][72],
F_[9][0][72],
F_[9][1][72],
F_[9][2][72],
F_[10][0][72],
F_[10][1][72],
F_[10][2][72],
F_[11][0][72],
F_[11][1][72],
F_[11][2][72],
F_[12][0][72],
F_[12][1][72],
F_[12][2][72],
F_[13][0][72],
F_[13][1][72],
F_[13][2][72],
F_[14][0][72],
F_[14][1][72],
F_[14][2][72],
F_[15][0][72],
F_[15][1][72],
F_[15][2][72],
F_[0][0][73],
F_[0][1][73],
F_[0][2][73],
F_[1][0][73],
F_[1][1][73],
F_[1][2][73],
F_[2][0][73],
F_[2][1][73],
F_[2][2][73],
F_[3][0][73],
F_[3][1][73],
F_[3][2][73],
F_[4][0][73],
F_[4][1][73],
F_[4][2][73],
F_[5][0][73],
F_[5][1][73],
F_[5][2][73],
F_[6][0][73],
F_[6][1][73],
F_[6][2][73],
F_[7][0][73],
F_[7][1][73],
F_[7][2][73],
F_[8][0][73],
F_[8][1][73],
F_[8][2][73],
F_[9][0][73],
F_[9][1][73],
F_[9][2][73],
F_[10][0][73],
F_[10][1][73],
F_[10][2][73],
F_[11][0][73],
F_[11][1][73],
F_[11][2][73],
F_[12][0][73],
F_[12][1][73],
F_[12][2][73],
F_[13][0][73],
F_[13][1][73],
F_[13][2][73],
F_[14][0][73],
F_[14][1][73],
F_[14][2][73],
F_[15][0][73],
F_[15][1][73],
F_[15][2][73],
F_[0][0][74],
F_[0][1][74],
F_[0][2][74],
F_[1][0][74],
F_[1][1][74],
F_[1][2][74],
F_[2][0][74],
F_[2][1][74],
F_[2][2][74],
F_[3][0][74],
F_[3][1][74],
F_[3][2][74],
F_[4][0][74],
F_[4][1][74],
F_[4][2][74],
F_[5][0][74],
F_[5][1][74],
F_[5][2][74],
F_[6][0][74],
F_[6][1][74],
F_[6][2][74],
F_[7][0][74],
F_[7][1][74],
F_[7][2][74],
F_[8][0][74],
F_[8][1][74],
F_[8][2][74],
F_[9][0][74],
F_[9][1][74],
F_[9][2][74],
F_[10][0][74],
F_[10][1][74],
F_[10][2][74],
F_[11][0][74],
F_[11][1][74],
F_[11][2][74],
F_[12][0][74],
F_[12][1][74],
F_[12][2][74],
F_[13][0][74],
F_[13][1][74],
F_[13][2][74],
F_[14][0][74],
F_[14][1][74],
F_[14][2][74],
F_[15][0][74],
F_[15][1][74],
F_[15][2][74],
F_[0][0][75],
F_[0][1][75],
F_[0][2][75],
F_[1][0][75],
F_[1][1][75],
F_[1][2][75],
F_[2][0][75],
F_[2][1][75],
F_[2][2][75],
F_[3][0][75],
F_[3][1][75],
F_[3][2][75],
F_[4][0][75],
F_[4][1][75],
F_[4][2][75],
F_[5][0][75],
F_[5][1][75],
F_[5][2][75],
F_[6][0][75],
F_[6][1][75],
F_[6][2][75],
F_[7][0][75],
F_[7][1][75],
F_[7][2][75],
F_[8][0][75],
F_[8][1][75],
F_[8][2][75],
F_[9][0][75],
F_[9][1][75],
F_[9][2][75],
F_[10][0][75],
F_[10][1][75],
F_[10][2][75],
F_[11][0][75],
F_[11][1][75],
F_[11][2][75],
F_[12][0][75],
F_[12][1][75],
F_[12][2][75],
F_[13][0][75],
F_[13][1][75],
F_[13][2][75],
F_[14][0][75],
F_[14][1][75],
F_[14][2][75],
F_[15][0][75],
F_[15][1][75],
F_[15][2][75],
F_[0][0][76],
F_[0][1][76],
F_[0][2][76],
F_[1][0][76],
F_[1][1][76],
F_[1][2][76],
F_[2][0][76],
F_[2][1][76],
F_[2][2][76],
F_[3][0][76],
F_[3][1][76],
F_[3][2][76],
F_[4][0][76],
F_[4][1][76],
F_[4][2][76],
F_[5][0][76],
F_[5][1][76],
F_[5][2][76],
F_[6][0][76],
F_[6][1][76],
F_[6][2][76],
F_[7][0][76],
F_[7][1][76],
F_[7][2][76],
F_[8][0][76],
F_[8][1][76],
F_[8][2][76],
F_[9][0][76],
F_[9][1][76],
F_[9][2][76],
F_[10][0][76],
F_[10][1][76],
F_[10][2][76],
F_[11][0][76],
F_[11][1][76],
F_[11][2][76],
F_[12][0][76],
F_[12][1][76],
F_[12][2][76],
F_[13][0][76],
F_[13][1][76],
F_[13][2][76],
F_[14][0][76],
F_[14][1][76],
F_[14][2][76],
F_[15][0][76],
F_[15][1][76],
F_[15][2][76],
F_[0][0][77],
F_[0][1][77],
F_[0][2][77],
F_[1][0][77],
F_[1][1][77],
F_[1][2][77],
F_[2][0][77],
F_[2][1][77],
F_[2][2][77],
F_[3][0][77],
F_[3][1][77],
F_[3][2][77],
F_[4][0][77],
F_[4][1][77],
F_[4][2][77],
F_[5][0][77],
F_[5][1][77],
F_[5][2][77],
F_[6][0][77],
F_[6][1][77],
F_[6][2][77],
F_[7][0][77],
F_[7][1][77],
F_[7][2][77],
F_[8][0][77],
F_[8][1][77],
F_[8][2][77],
F_[9][0][77],
F_[9][1][77],
F_[9][2][77],
F_[10][0][77],
F_[10][1][77],
F_[10][2][77],
F_[11][0][77],
F_[11][1][77],
F_[11][2][77],
F_[12][0][77],
F_[12][1][77],
F_[12][2][77],
F_[13][0][77],
F_[13][1][77],
F_[13][2][77],
F_[14][0][77],
F_[14][1][77],
F_[14][2][77],
F_[15][0][77],
F_[15][1][77],
F_[15][2][77],
F_[0][0][78],
F_[0][1][78],
F_[0][2][78],
F_[1][0][78],
F_[1][1][78],
F_[1][2][78],
F_[2][0][78],
F_[2][1][78],
F_[2][2][78],
F_[3][0][78],
F_[3][1][78],
F_[3][2][78],
F_[4][0][78],
F_[4][1][78],
F_[4][2][78],
F_[5][0][78],
F_[5][1][78],
F_[5][2][78],
F_[6][0][78],
F_[6][1][78],
F_[6][2][78],
F_[7][0][78],
F_[7][1][78],
F_[7][2][78],
F_[8][0][78],
F_[8][1][78],
F_[8][2][78],
F_[9][0][78],
F_[9][1][78],
F_[9][2][78],
F_[10][0][78],
F_[10][1][78],
F_[10][2][78],
F_[11][0][78],
F_[11][1][78],
F_[11][2][78],
F_[12][0][78],
F_[12][1][78],
F_[12][2][78],
F_[13][0][78],
F_[13][1][78],
F_[13][2][78],
F_[14][0][78],
F_[14][1][78],
F_[14][2][78],
F_[15][0][78],
F_[15][1][78],
F_[15][2][78],
F_[0][0][79],
F_[0][1][79],
F_[0][2][79],
F_[1][0][79],
F_[1][1][79],
F_[1][2][79],
F_[2][0][79],
F_[2][1][79],
F_[2][2][79],
F_[3][0][79],
F_[3][1][79],
F_[3][2][79],
F_[4][0][79],
F_[4][1][79],
F_[4][2][79],
F_[5][0][79],
F_[5][1][79],
F_[5][2][79],
F_[6][0][79],
F_[6][1][79],
F_[6][2][79],
F_[7][0][79],
F_[7][1][79],
F_[7][2][79],
F_[8][0][79],
F_[8][1][79],
F_[8][2][79],
F_[9][0][79],
F_[9][1][79],
F_[9][2][79],
F_[10][0][79],
F_[10][1][79],
F_[10][2][79],
F_[11][0][79],
F_[11][1][79],
F_[11][2][79],
F_[12][0][79],
F_[12][1][79],
F_[12][2][79],
F_[13][0][79],
F_[13][1][79],
F_[13][2][79],
F_[14][0][79],
F_[14][1][79],
F_[14][2][79],
F_[15][0][79],
F_[15][1][79],
F_[15][2][79],
F_[0][0][80],
F_[0][1][80],
F_[0][2][80],
F_[1][0][80],
F_[1][1][80],
F_[1][2][80],
F_[2][0][80],
F_[2][1][80],
F_[2][2][80],
F_[3][0][80],
F_[3][1][80],
F_[3][2][80],
F_[4][0][80],
F_[4][1][80],
F_[4][2][80],
F_[5][0][80],
F_[5][1][80],
F_[5][2][80],
F_[6][0][80],
F_[6][1][80],
F_[6][2][80],
F_[7][0][80],
F_[7][1][80],
F_[7][2][80],
F_[8][0][80],
F_[8][1][80],
F_[8][2][80],
F_[9][0][80],
F_[9][1][80],
F_[9][2][80],
F_[10][0][80],
F_[10][1][80],
F_[10][2][80],
F_[11][0][80],
F_[11][1][80],
F_[11][2][80],
F_[12][0][80],
F_[12][1][80],
F_[12][2][80],
F_[13][0][80],
F_[13][1][80],
F_[13][2][80],
F_[14][0][80],
F_[14][1][80],
F_[14][2][80],
F_[15][0][80],
F_[15][1][80],
F_[15][2][80],
F_[0][0][81],
F_[0][1][81],
F_[0][2][81],
F_[1][0][81],
F_[1][1][81],
F_[1][2][81],
F_[2][0][81],
F_[2][1][81],
F_[2][2][81],
F_[3][0][81],
F_[3][1][81],
F_[3][2][81],
F_[4][0][81],
F_[4][1][81],
F_[4][2][81],
F_[5][0][81],
F_[5][1][81],
F_[5][2][81],
F_[6][0][81],
F_[6][1][81],
F_[6][2][81],
F_[7][0][81],
F_[7][1][81],
F_[7][2][81],
F_[8][0][81],
F_[8][1][81],
F_[8][2][81],
F_[9][0][81],
F_[9][1][81],
F_[9][2][81],
F_[10][0][81],
F_[10][1][81],
F_[10][2][81],
F_[11][0][81],
F_[11][1][81],
F_[11][2][81],
F_[12][0][81],
F_[12][1][81],
F_[12][2][81],
F_[13][0][81],
F_[13][1][81],
F_[13][2][81],
F_[14][0][81],
F_[14][1][81],
F_[14][2][81],
F_[15][0][81],
F_[15][1][81],
F_[15][2][81],
F_[0][0][82],
F_[0][1][82],
F_[0][2][82],
F_[1][0][82],
F_[1][1][82],
F_[1][2][82],
F_[2][0][82],
F_[2][1][82],
F_[2][2][82],
F_[3][0][82],
F_[3][1][82],
F_[3][2][82],
F_[4][0][82],
F_[4][1][82],
F_[4][2][82],
F_[5][0][82],
F_[5][1][82],
F_[5][2][82],
F_[6][0][82],
F_[6][1][82],
F_[6][2][82],
F_[7][0][82],
F_[7][1][82],
F_[7][2][82],
F_[8][0][82],
F_[8][1][82],
F_[8][2][82],
F_[9][0][82],
F_[9][1][82],
F_[9][2][82],
F_[10][0][82],
F_[10][1][82],
F_[10][2][82],
F_[11][0][82],
F_[11][1][82],
F_[11][2][82],
F_[12][0][82],
F_[12][1][82],
F_[12][2][82],
F_[13][0][82],
F_[13][1][82],
F_[13][2][82],
F_[14][0][82],
F_[14][1][82],
F_[14][2][82],
F_[15][0][82],
F_[15][1][82],
F_[15][2][82],
F_[0][0][83],
F_[0][1][83],
F_[0][2][83],
F_[1][0][83],
F_[1][1][83],
F_[1][2][83],
F_[2][0][83],
F_[2][1][83],
F_[2][2][83],
F_[3][0][83],
F_[3][1][83],
F_[3][2][83],
F_[4][0][83],
F_[4][1][83],
F_[4][2][83],
F_[5][0][83],
F_[5][1][83],
F_[5][2][83],
F_[6][0][83],
F_[6][1][83],
F_[6][2][83],
F_[7][0][83],
F_[7][1][83],
F_[7][2][83],
F_[8][0][83],
F_[8][1][83],
F_[8][2][83],
F_[9][0][83],
F_[9][1][83],
F_[9][2][83],
F_[10][0][83],
F_[10][1][83],
F_[10][2][83],
F_[11][0][83],
F_[11][1][83],
F_[11][2][83],
F_[12][0][83],
F_[12][1][83],
F_[12][2][83],
F_[13][0][83],
F_[13][1][83],
F_[13][2][83],
F_[14][0][83],
F_[14][1][83],
F_[14][2][83],
F_[15][0][83],
F_[15][1][83],
F_[15][2][83],
F_[0][0][84],
F_[0][1][84],
F_[0][2][84],
F_[1][0][84],
F_[1][1][84],
F_[1][2][84],
F_[2][0][84],
F_[2][1][84],
F_[2][2][84],
F_[3][0][84],
F_[3][1][84],
F_[3][2][84],
F_[4][0][84],
F_[4][1][84],
F_[4][2][84],
F_[5][0][84],
F_[5][1][84],
F_[5][2][84],
F_[6][0][84],
F_[6][1][84],
F_[6][2][84],
F_[7][0][84],
F_[7][1][84],
F_[7][2][84],
F_[8][0][84],
F_[8][1][84],
F_[8][2][84],
F_[9][0][84],
F_[9][1][84],
F_[9][2][84],
F_[10][0][84],
F_[10][1][84],
F_[10][2][84],
F_[11][0][84],
F_[11][1][84],
F_[11][2][84],
F_[12][0][84],
F_[12][1][84],
F_[12][2][84],
F_[13][0][84],
F_[13][1][84],
F_[13][2][84],
F_[14][0][84],
F_[14][1][84],
F_[14][2][84],
F_[15][0][84],
F_[15][1][84],
F_[15][2][84],
F_[0][0][85],
F_[0][1][85],
F_[0][2][85],
F_[1][0][85],
F_[1][1][85],
F_[1][2][85],
F_[2][0][85],
F_[2][1][85],
F_[2][2][85],
F_[3][0][85],
F_[3][1][85],
F_[3][2][85],
F_[4][0][85],
F_[4][1][85],
F_[4][2][85],
F_[5][0][85],
F_[5][1][85],
F_[5][2][85],
F_[6][0][85],
F_[6][1][85],
F_[6][2][85],
F_[7][0][85],
F_[7][1][85],
F_[7][2][85],
F_[8][0][85],
F_[8][1][85],
F_[8][2][85],
F_[9][0][85],
F_[9][1][85],
F_[9][2][85],
F_[10][0][85],
F_[10][1][85],
F_[10][2][85],
F_[11][0][85],
F_[11][1][85],
F_[11][2][85],
F_[12][0][85],
F_[12][1][85],
F_[12][2][85],
F_[13][0][85],
F_[13][1][85],
F_[13][2][85],
F_[14][0][85],
F_[14][1][85],
F_[14][2][85],
F_[15][0][85],
F_[15][1][85],
F_[15][2][85],
F_[0][0][86],
F_[0][1][86],
F_[0][2][86],
F_[1][0][86],
F_[1][1][86],
F_[1][2][86],
F_[2][0][86],
F_[2][1][86],
F_[2][2][86],
F_[3][0][86],
F_[3][1][86],
F_[3][2][86],
F_[4][0][86],
F_[4][1][86],
F_[4][2][86],
F_[5][0][86],
F_[5][1][86],
F_[5][2][86],
F_[6][0][86],
F_[6][1][86],
F_[6][2][86],
F_[7][0][86],
F_[7][1][86],
F_[7][2][86],
F_[8][0][86],
F_[8][1][86],
F_[8][2][86],
F_[9][0][86],
F_[9][1][86],
F_[9][2][86],
F_[10][0][86],
F_[10][1][86],
F_[10][2][86],
F_[11][0][86],
F_[11][1][86],
F_[11][2][86],
F_[12][0][86],
F_[12][1][86],
F_[12][2][86],
F_[13][0][86],
F_[13][1][86],
F_[13][2][86],
F_[14][0][86],
F_[14][1][86],
F_[14][2][86],
F_[15][0][86],
F_[15][1][86],
F_[15][2][86],
F_[0][0][87],
F_[0][1][87],
F_[0][2][87],
F_[1][0][87],
F_[1][1][87],
F_[1][2][87],
F_[2][0][87],
F_[2][1][87],
F_[2][2][87],
F_[3][0][87],
F_[3][1][87],
F_[3][2][87],
F_[4][0][87],
F_[4][1][87],
F_[4][2][87],
F_[5][0][87],
F_[5][1][87],
F_[5][2][87],
F_[6][0][87],
F_[6][1][87],
F_[6][2][87],
F_[7][0][87],
F_[7][1][87],
F_[7][2][87],
F_[8][0][87],
F_[8][1][87],
F_[8][2][87],
F_[9][0][87],
F_[9][1][87],
F_[9][2][87],
F_[10][0][87],
F_[10][1][87],
F_[10][2][87],
F_[11][0][87],
F_[11][1][87],
F_[11][2][87],
F_[12][0][87],
F_[12][1][87],
F_[12][2][87],
F_[13][0][87],
F_[13][1][87],
F_[13][2][87],
F_[14][0][87],
F_[14][1][87],
F_[14][2][87],
F_[15][0][87],
F_[15][1][87],
F_[15][2][87],
F_[0][0][88],
F_[0][1][88],
F_[0][2][88],
F_[1][0][88],
F_[1][1][88],
F_[1][2][88],
F_[2][0][88],
F_[2][1][88],
F_[2][2][88],
F_[3][0][88],
F_[3][1][88],
F_[3][2][88],
F_[4][0][88],
F_[4][1][88],
F_[4][2][88],
F_[5][0][88],
F_[5][1][88],
F_[5][2][88],
F_[6][0][88],
F_[6][1][88],
F_[6][2][88],
F_[7][0][88],
F_[7][1][88],
F_[7][2][88],
F_[8][0][88],
F_[8][1][88],
F_[8][2][88],
F_[9][0][88],
F_[9][1][88],
F_[9][2][88],
F_[10][0][88],
F_[10][1][88],
F_[10][2][88],
F_[11][0][88],
F_[11][1][88],
F_[11][2][88],
F_[12][0][88],
F_[12][1][88],
F_[12][2][88],
F_[13][0][88],
F_[13][1][88],
F_[13][2][88],
F_[14][0][88],
F_[14][1][88],
F_[14][2][88],
F_[15][0][88],
F_[15][1][88],
F_[15][2][88],
F_[0][0][89],
F_[0][1][89],
F_[0][2][89],
F_[1][0][89],
F_[1][1][89],
F_[1][2][89],
F_[2][0][89],
F_[2][1][89],
F_[2][2][89],
F_[3][0][89],
F_[3][1][89],
F_[3][2][89],
F_[4][0][89],
F_[4][1][89],
F_[4][2][89],
F_[5][0][89],
F_[5][1][89],
F_[5][2][89],
F_[6][0][89],
F_[6][1][89],
F_[6][2][89],
F_[7][0][89],
F_[7][1][89],
F_[7][2][89],
F_[8][0][89],
F_[8][1][89],
F_[8][2][89],
F_[9][0][89],
F_[9][1][89],
F_[9][2][89],
F_[10][0][89],
F_[10][1][89],
F_[10][2][89],
F_[11][0][89],
F_[11][1][89],
F_[11][2][89],
F_[12][0][89],
F_[12][1][89],
F_[12][2][89],
F_[13][0][89],
F_[13][1][89],
F_[13][2][89],
F_[14][0][89],
F_[14][1][89],
F_[14][2][89],
F_[15][0][89],
F_[15][1][89],
F_[15][2][89],
F_[0][0][90],
F_[0][1][90],
F_[0][2][90],
F_[1][0][90],
F_[1][1][90],
F_[1][2][90],
F_[2][0][90],
F_[2][1][90],
F_[2][2][90],
F_[3][0][90],
F_[3][1][90],
F_[3][2][90],
F_[4][0][90],
F_[4][1][90],
F_[4][2][90],
F_[5][0][90],
F_[5][1][90],
F_[5][2][90],
F_[6][0][90],
F_[6][1][90],
F_[6][2][90],
F_[7][0][90],
F_[7][1][90],
F_[7][2][90],
F_[8][0][90],
F_[8][1][90],
F_[8][2][90],
F_[9][0][90],
F_[9][1][90],
F_[9][2][90],
F_[10][0][90],
F_[10][1][90],
F_[10][2][90],
F_[11][0][90],
F_[11][1][90],
F_[11][2][90],
F_[12][0][90],
F_[12][1][90],
F_[12][2][90],
F_[13][0][90],
F_[13][1][90],
F_[13][2][90],
F_[14][0][90],
F_[14][1][90],
F_[14][2][90],
F_[15][0][90],
F_[15][1][90],
F_[15][2][90],
F_[0][0][91],
F_[0][1][91],
F_[0][2][91],
F_[1][0][91],
F_[1][1][91],
F_[1][2][91],
F_[2][0][91],
F_[2][1][91],
F_[2][2][91],
F_[3][0][91],
F_[3][1][91],
F_[3][2][91],
F_[4][0][91],
F_[4][1][91],
F_[4][2][91],
F_[5][0][91],
F_[5][1][91],
F_[5][2][91],
F_[6][0][91],
F_[6][1][91],
F_[6][2][91],
F_[7][0][91],
F_[7][1][91],
F_[7][2][91],
F_[8][0][91],
F_[8][1][91],
F_[8][2][91],
F_[9][0][91],
F_[9][1][91],
F_[9][2][91],
F_[10][0][91],
F_[10][1][91],
F_[10][2][91],
F_[11][0][91],
F_[11][1][91],
F_[11][2][91],
F_[12][0][91],
F_[12][1][91],
F_[12][2][91],
F_[13][0][91],
F_[13][1][91],
F_[13][2][91],
F_[14][0][91],
F_[14][1][91],
F_[14][2][91],
F_[15][0][91],
F_[15][1][91],
F_[15][2][91],
F_[0][0][92],
F_[0][1][92],
F_[0][2][92],
F_[1][0][92],
F_[1][1][92],
F_[1][2][92],
F_[2][0][92],
F_[2][1][92],
F_[2][2][92],
F_[3][0][92],
F_[3][1][92],
F_[3][2][92],
F_[4][0][92],
F_[4][1][92],
F_[4][2][92],
F_[5][0][92],
F_[5][1][92],
F_[5][2][92],
F_[6][0][92],
F_[6][1][92],
F_[6][2][92],
F_[7][0][92],
F_[7][1][92],
F_[7][2][92],
F_[8][0][92],
F_[8][1][92],
F_[8][2][92],
F_[9][0][92],
F_[9][1][92],
F_[9][2][92],
F_[10][0][92],
F_[10][1][92],
F_[10][2][92],
F_[11][0][92],
F_[11][1][92],
F_[11][2][92],
F_[12][0][92],
F_[12][1][92],
F_[12][2][92],
F_[13][0][92],
F_[13][1][92],
F_[13][2][92],
F_[14][0][92],
F_[14][1][92],
F_[14][2][92],
F_[15][0][92],
F_[15][1][92],
F_[15][2][92],
F_[0][0][93],
F_[0][1][93],
F_[0][2][93],
F_[1][0][93],
F_[1][1][93],
F_[1][2][93],
F_[2][0][93],
F_[2][1][93],
F_[2][2][93],
F_[3][0][93],
F_[3][1][93],
F_[3][2][93],
F_[4][0][93],
F_[4][1][93],
F_[4][2][93],
F_[5][0][93],
F_[5][1][93],
F_[5][2][93],
F_[6][0][93],
F_[6][1][93],
F_[6][2][93],
F_[7][0][93],
F_[7][1][93],
F_[7][2][93],
F_[8][0][93],
F_[8][1][93],
F_[8][2][93],
F_[9][0][93],
F_[9][1][93],
F_[9][2][93],
F_[10][0][93],
F_[10][1][93],
F_[10][2][93],
F_[11][0][93],
F_[11][1][93],
F_[11][2][93],
F_[12][0][93],
F_[12][1][93],
F_[12][2][93],
F_[13][0][93],
F_[13][1][93],
F_[13][2][93],
F_[14][0][93],
F_[14][1][93],
F_[14][2][93],
F_[15][0][93],
F_[15][1][93],
F_[15][2][93],
F_[0][0][94],
F_[0][1][94],
F_[0][2][94],
F_[1][0][94],
F_[1][1][94],
F_[1][2][94],
F_[2][0][94],
F_[2][1][94],
F_[2][2][94],
F_[3][0][94],
F_[3][1][94],
F_[3][2][94],
F_[4][0][94],
F_[4][1][94],
F_[4][2][94],
F_[5][0][94],
F_[5][1][94],
F_[5][2][94],
F_[6][0][94],
F_[6][1][94],
F_[6][2][94],
F_[7][0][94],
F_[7][1][94],
F_[7][2][94],
F_[8][0][94],
F_[8][1][94],
F_[8][2][94],
F_[9][0][94],
F_[9][1][94],
F_[9][2][94],
F_[10][0][94],
F_[10][1][94],
F_[10][2][94],
F_[11][0][94],
F_[11][1][94],
F_[11][2][94],
F_[12][0][94],
F_[12][1][94],
F_[12][2][94],
F_[13][0][94],
F_[13][1][94],
F_[13][2][94],
F_[14][0][94],
F_[14][1][94],
F_[14][2][94],
F_[15][0][94],
F_[15][1][94],
F_[15][2][94],
F_[0][0][95],
F_[0][1][95],
F_[0][2][95],
F_[1][0][95],
F_[1][1][95],
F_[1][2][95],
F_[2][0][95],
F_[2][1][95],
F_[2][2][95],
F_[3][0][95],
F_[3][1][95],
F_[3][2][95],
F_[4][0][95],
F_[4][1][95],
F_[4][2][95],
F_[5][0][95],
F_[5][1][95],
F_[5][2][95],
F_[6][0][95],
F_[6][1][95],
F_[6][2][95],
F_[7][0][95],
F_[7][1][95],
F_[7][2][95],
F_[8][0][95],
F_[8][1][95],
F_[8][2][95],
F_[9][0][95],
F_[9][1][95],
F_[9][2][95],
F_[10][0][95],
F_[10][1][95],
F_[10][2][95],
F_[11][0][95],
F_[11][1][95],
F_[11][2][95],
F_[12][0][95],
F_[12][1][95],
F_[12][2][95],
F_[13][0][95],
F_[13][1][95],
F_[13][2][95],
F_[14][0][95],
F_[14][1][95],
F_[14][2][95],
F_[15][0][95],
F_[15][1][95],
F_[15][2][95],
F_[0][0][96],
F_[0][1][96],
F_[0][2][96],
F_[1][0][96],
F_[1][1][96],
F_[1][2][96],
F_[2][0][96],
F_[2][1][96],
F_[2][2][96],
F_[3][0][96],
F_[3][1][96],
F_[3][2][96],
F_[4][0][96],
F_[4][1][96],
F_[4][2][96],
F_[5][0][96],
F_[5][1][96],
F_[5][2][96],
F_[6][0][96],
F_[6][1][96],
F_[6][2][96],
F_[7][0][96],
F_[7][1][96],
F_[7][2][96],
F_[8][0][96],
F_[8][1][96],
F_[8][2][96],
F_[9][0][96],
F_[9][1][96],
F_[9][2][96],
F_[10][0][96],
F_[10][1][96],
F_[10][2][96],
F_[11][0][96],
F_[11][1][96],
F_[11][2][96],
F_[12][0][96],
F_[12][1][96],
F_[12][2][96],
F_[13][0][96],
F_[13][1][96],
F_[13][2][96],
F_[14][0][96],
F_[14][1][96],
F_[14][2][96],
F_[15][0][96],
F_[15][1][96],
F_[15][2][96],
F_[0][0][97],
F_[0][1][97],
F_[0][2][97],
F_[1][0][97],
F_[1][1][97],
F_[1][2][97],
F_[2][0][97],
F_[2][1][97],
F_[2][2][97],
F_[3][0][97],
F_[3][1][97],
F_[3][2][97],
F_[4][0][97],
F_[4][1][97],
F_[4][2][97],
F_[5][0][97],
F_[5][1][97],
F_[5][2][97],
F_[6][0][97],
F_[6][1][97],
F_[6][2][97],
F_[7][0][97],
F_[7][1][97],
F_[7][2][97],
F_[8][0][97],
F_[8][1][97],
F_[8][2][97],
F_[9][0][97],
F_[9][1][97],
F_[9][2][97],
F_[10][0][97],
F_[10][1][97],
F_[10][2][97],
F_[11][0][97],
F_[11][1][97],
F_[11][2][97],
F_[12][0][97],
F_[12][1][97],
F_[12][2][97],
F_[13][0][97],
F_[13][1][97],
F_[13][2][97],
F_[14][0][97],
F_[14][1][97],
F_[14][2][97],
F_[15][0][97],
F_[15][1][97],
F_[15][2][97],
F_[0][0][98],
F_[0][1][98],
F_[0][2][98],
F_[1][0][98],
F_[1][1][98],
F_[1][2][98],
F_[2][0][98],
F_[2][1][98],
F_[2][2][98],
F_[3][0][98],
F_[3][1][98],
F_[3][2][98],
F_[4][0][98],
F_[4][1][98],
F_[4][2][98],
F_[5][0][98],
F_[5][1][98],
F_[5][2][98],
F_[6][0][98],
F_[6][1][98],
F_[6][2][98],
F_[7][0][98],
F_[7][1][98],
F_[7][2][98],
F_[8][0][98],
F_[8][1][98],
F_[8][2][98],
F_[9][0][98],
F_[9][1][98],
F_[9][2][98],
F_[10][0][98],
F_[10][1][98],
F_[10][2][98],
F_[11][0][98],
F_[11][1][98],
F_[11][2][98],
F_[12][0][98],
F_[12][1][98],
F_[12][2][98],
F_[13][0][98],
F_[13][1][98],
F_[13][2][98],
F_[14][0][98],
F_[14][1][98],
F_[14][2][98],
F_[15][0][98],
F_[15][1][98],
F_[15][2][98],
F_[0][0][99],
F_[0][1][99],
F_[0][2][99],
F_[1][0][99],
F_[1][1][99],
F_[1][2][99],
F_[2][0][99],
F_[2][1][99],
F_[2][2][99],
F_[3][0][99],
F_[3][1][99],
F_[3][2][99],
F_[4][0][99],
F_[4][1][99],
F_[4][2][99],
F_[5][0][99],
F_[5][1][99],
F_[5][2][99],
F_[6][0][99],
F_[6][1][99],
F_[6][2][99],
F_[7][0][99],
F_[7][1][99],
F_[7][2][99],
F_[8][0][99],
F_[8][1][99],
F_[8][2][99],
F_[9][0][99],
F_[9][1][99],
F_[9][2][99],
F_[10][0][99],
F_[10][1][99],
F_[10][2][99],
F_[11][0][99],
F_[11][1][99],
F_[11][2][99],
F_[12][0][99],
F_[12][1][99],
F_[12][2][99],
F_[13][0][99],
F_[13][1][99],
F_[13][2][99],
F_[14][0][99],
F_[14][1][99],
F_[14][2][99],
F_[15][0][99],
F_[15][1][99],
F_[15][2][99],
F_[0][0][100],
F_[0][1][100],
F_[0][2][100],
F_[1][0][100],
F_[1][1][100],
F_[1][2][100],
F_[2][0][100],
F_[2][1][100],
F_[2][2][100],
F_[3][0][100],
F_[3][1][100],
F_[3][2][100],
F_[4][0][100],
F_[4][1][100],
F_[4][2][100],
F_[5][0][100],
F_[5][1][100],
F_[5][2][100],
F_[6][0][100],
F_[6][1][100],
F_[6][2][100],
F_[7][0][100],
F_[7][1][100],
F_[7][2][100],
F_[8][0][100],
F_[8][1][100],
F_[8][2][100],
F_[9][0][100],
F_[9][1][100],
F_[9][2][100],
F_[10][0][100],
F_[10][1][100],
F_[10][2][100],
F_[11][0][100],
F_[11][1][100],
F_[11][2][100],
F_[12][0][100],
F_[12][1][100],
F_[12][2][100],
F_[13][0][100],
F_[13][1][100],
F_[13][2][100],
F_[14][0][100],
F_[14][1][100],
F_[14][2][100],
F_[15][0][100],
F_[15][1][100],
F_[15][2][100],
F_[0][0][101],
F_[0][1][101],
F_[0][2][101],
F_[1][0][101],
F_[1][1][101],
F_[1][2][101],
F_[2][0][101],
F_[2][1][101],
F_[2][2][101],
F_[3][0][101],
F_[3][1][101],
F_[3][2][101],
F_[4][0][101],
F_[4][1][101],
F_[4][2][101],
F_[5][0][101],
F_[5][1][101],
F_[5][2][101],
F_[6][0][101],
F_[6][1][101],
F_[6][2][101],
F_[7][0][101],
F_[7][1][101],
F_[7][2][101],
F_[8][0][101],
F_[8][1][101],
F_[8][2][101],
F_[9][0][101],
F_[9][1][101],
F_[9][2][101],
F_[10][0][101],
F_[10][1][101],
F_[10][2][101],
F_[11][0][101],
F_[11][1][101],
F_[11][2][101],
F_[12][0][101],
F_[12][1][101],
F_[12][2][101],
F_[13][0][101],
F_[13][1][101],
F_[13][2][101],
F_[14][0][101],
F_[14][1][101],
F_[14][2][101],
F_[15][0][101],
F_[15][1][101],
F_[15][2][101],
F_[0][0][102],
F_[0][1][102],
F_[0][2][102],
F_[1][0][102],
F_[1][1][102],
F_[1][2][102],
F_[2][0][102],
F_[2][1][102],
F_[2][2][102],
F_[3][0][102],
F_[3][1][102],
F_[3][2][102],
F_[4][0][102],
F_[4][1][102],
F_[4][2][102],
F_[5][0][102],
F_[5][1][102],
F_[5][2][102],
F_[6][0][102],
F_[6][1][102],
F_[6][2][102],
F_[7][0][102],
F_[7][1][102],
F_[7][2][102],
F_[8][0][102],
F_[8][1][102],
F_[8][2][102],
F_[9][0][102],
F_[9][1][102],
F_[9][2][102],
F_[10][0][102],
F_[10][1][102],
F_[10][2][102],
F_[11][0][102],
F_[11][1][102],
F_[11][2][102],
F_[12][0][102],
F_[12][1][102],
F_[12][2][102],
F_[13][0][102],
F_[13][1][102],
F_[13][2][102],
F_[14][0][102],
F_[14][1][102],
F_[14][2][102],
F_[15][0][102],
F_[15][1][102],
F_[15][2][102],
F_[0][0][103],
F_[0][1][103],
F_[0][2][103],
F_[1][0][103],
F_[1][1][103],
F_[1][2][103],
F_[2][0][103],
F_[2][1][103],
F_[2][2][103],
F_[3][0][103],
F_[3][1][103],
F_[3][2][103],
F_[4][0][103],
F_[4][1][103],
F_[4][2][103],
F_[5][0][103],
F_[5][1][103],
F_[5][2][103],
F_[6][0][103],
F_[6][1][103],
F_[6][2][103],
F_[7][0][103],
F_[7][1][103],
F_[7][2][103],
F_[8][0][103],
F_[8][1][103],
F_[8][2][103],
F_[9][0][103],
F_[9][1][103],
F_[9][2][103],
F_[10][0][103],
F_[10][1][103],
F_[10][2][103],
F_[11][0][103],
F_[11][1][103],
F_[11][2][103],
F_[12][0][103],
F_[12][1][103],
F_[12][2][103],
F_[13][0][103],
F_[13][1][103],
F_[13][2][103],
F_[14][0][103],
F_[14][1][103],
F_[14][2][103],
F_[15][0][103],
F_[15][1][103],
F_[15][2][103],
F_[0][0][104],
F_[0][1][104],
F_[0][2][104],
F_[1][0][104],
F_[1][1][104],
F_[1][2][104],
F_[2][0][104],
F_[2][1][104],
F_[2][2][104],
F_[3][0][104],
F_[3][1][104],
F_[3][2][104],
F_[4][0][104],
F_[4][1][104],
F_[4][2][104],
F_[5][0][104],
F_[5][1][104],
F_[5][2][104],
F_[6][0][104],
F_[6][1][104],
F_[6][2][104],
F_[7][0][104],
F_[7][1][104],
F_[7][2][104],
F_[8][0][104],
F_[8][1][104],
F_[8][2][104],
F_[9][0][104],
F_[9][1][104],
F_[9][2][104],
F_[10][0][104],
F_[10][1][104],
F_[10][2][104],
F_[11][0][104],
F_[11][1][104],
F_[11][2][104],
F_[12][0][104],
F_[12][1][104],
F_[12][2][104],
F_[13][0][104],
F_[13][1][104],
F_[13][2][104],
F_[14][0][104],
F_[14][1][104],
F_[14][2][104],
F_[15][0][104],
F_[15][1][104],
F_[15][2][104],
F_[0][0][105],
F_[0][1][105],
F_[0][2][105],
F_[1][0][105],
F_[1][1][105],
F_[1][2][105],
F_[2][0][105],
F_[2][1][105],
F_[2][2][105],
F_[3][0][105],
F_[3][1][105],
F_[3][2][105],
F_[4][0][105],
F_[4][1][105],
F_[4][2][105],
F_[5][0][105],
F_[5][1][105],
F_[5][2][105],
F_[6][0][105],
F_[6][1][105],
F_[6][2][105],
F_[7][0][105],
F_[7][1][105],
F_[7][2][105],
F_[8][0][105],
F_[8][1][105],
F_[8][2][105],
F_[9][0][105],
F_[9][1][105],
F_[9][2][105],
F_[10][0][105],
F_[10][1][105],
F_[10][2][105],
F_[11][0][105],
F_[11][1][105],
F_[11][2][105],
F_[12][0][105],
F_[12][1][105],
F_[12][2][105],
F_[13][0][105],
F_[13][1][105],
F_[13][2][105],
F_[14][0][105],
F_[14][1][105],
F_[14][2][105],
F_[15][0][105],
F_[15][1][105],
F_[15][2][105],
F_[0][0][106],
F_[0][1][106],
F_[0][2][106],
F_[1][0][106],
F_[1][1][106],
F_[1][2][106],
F_[2][0][106],
F_[2][1][106],
F_[2][2][106],
F_[3][0][106],
F_[3][1][106],
F_[3][2][106],
F_[4][0][106],
F_[4][1][106],
F_[4][2][106],
F_[5][0][106],
F_[5][1][106],
F_[5][2][106],
F_[6][0][106],
F_[6][1][106],
F_[6][2][106],
F_[7][0][106],
F_[7][1][106],
F_[7][2][106],
F_[8][0][106],
F_[8][1][106],
F_[8][2][106],
F_[9][0][106],
F_[9][1][106],
F_[9][2][106],
F_[10][0][106],
F_[10][1][106],
F_[10][2][106],
F_[11][0][106],
F_[11][1][106],
F_[11][2][106],
F_[12][0][106],
F_[12][1][106],
F_[12][2][106],
F_[13][0][106],
F_[13][1][106],
F_[13][2][106],
F_[14][0][106],
F_[14][1][106],
F_[14][2][106],
F_[15][0][106],
F_[15][1][106],
F_[15][2][106],
F_[0][0][107],
F_[0][1][107],
F_[0][2][107],
F_[1][0][107],
F_[1][1][107],
F_[1][2][107],
F_[2][0][107],
F_[2][1][107],
F_[2][2][107],
F_[3][0][107],
F_[3][1][107],
F_[3][2][107],
F_[4][0][107],
F_[4][1][107],
F_[4][2][107],
F_[5][0][107],
F_[5][1][107],
F_[5][2][107],
F_[6][0][107],
F_[6][1][107],
F_[6][2][107],
F_[7][0][107],
F_[7][1][107],
F_[7][2][107],
F_[8][0][107],
F_[8][1][107],
F_[8][2][107],
F_[9][0][107],
F_[9][1][107],
F_[9][2][107],
F_[10][0][107],
F_[10][1][107],
F_[10][2][107],
F_[11][0][107],
F_[11][1][107],
F_[11][2][107],
F_[12][0][107],
F_[12][1][107],
F_[12][2][107],
F_[13][0][107],
F_[13][1][107],
F_[13][2][107],
F_[14][0][107],
F_[14][1][107],
F_[14][2][107],
F_[15][0][107],
F_[15][1][107],
F_[15][2][107],
F_[0][0][108],
F_[0][1][108],
F_[0][2][108],
F_[1][0][108],
F_[1][1][108],
F_[1][2][108],
F_[2][0][108],
F_[2][1][108],
F_[2][2][108],
F_[3][0][108],
F_[3][1][108],
F_[3][2][108],
F_[4][0][108],
F_[4][1][108],
F_[4][2][108],
F_[5][0][108],
F_[5][1][108],
F_[5][2][108],
F_[6][0][108],
F_[6][1][108],
F_[6][2][108],
F_[7][0][108],
F_[7][1][108],
F_[7][2][108],
F_[8][0][108],
F_[8][1][108],
F_[8][2][108],
F_[9][0][108],
F_[9][1][108],
F_[9][2][108],
F_[10][0][108],
F_[10][1][108],
F_[10][2][108],
F_[11][0][108],
F_[11][1][108],
F_[11][2][108],
F_[12][0][108],
F_[12][1][108],
F_[12][2][108],
F_[13][0][108],
F_[13][1][108],
F_[13][2][108],
F_[14][0][108],
F_[14][1][108],
F_[14][2][108],
F_[15][0][108],
F_[15][1][108],
F_[15][2][108],
F_[0][0][109],
F_[0][1][109],
F_[0][2][109],
F_[1][0][109],
F_[1][1][109],
F_[1][2][109],
F_[2][0][109],
F_[2][1][109],
F_[2][2][109],
F_[3][0][109],
F_[3][1][109],
F_[3][2][109],
F_[4][0][109],
F_[4][1][109],
F_[4][2][109],
F_[5][0][109],
F_[5][1][109],
F_[5][2][109],
F_[6][0][109],
F_[6][1][109],
F_[6][2][109],
F_[7][0][109],
F_[7][1][109],
F_[7][2][109],
F_[8][0][109],
F_[8][1][109],
F_[8][2][109],
F_[9][0][109],
F_[9][1][109],
F_[9][2][109],
F_[10][0][109],
F_[10][1][109],
F_[10][2][109],
F_[11][0][109],
F_[11][1][109],
F_[11][2][109],
F_[12][0][109],
F_[12][1][109],
F_[12][2][109],
F_[13][0][109],
F_[13][1][109],
F_[13][2][109],
F_[14][0][109],
F_[14][1][109],
F_[14][2][109],
F_[15][0][109],
F_[15][1][109],
F_[15][2][109],
F_[0][0][110],
F_[0][1][110],
F_[0][2][110],
F_[1][0][110],
F_[1][1][110],
F_[1][2][110],
F_[2][0][110],
F_[2][1][110],
F_[2][2][110],
F_[3][0][110],
F_[3][1][110],
F_[3][2][110],
F_[4][0][110],
F_[4][1][110],
F_[4][2][110],
F_[5][0][110],
F_[5][1][110],
F_[5][2][110],
F_[6][0][110],
F_[6][1][110],
F_[6][2][110],
F_[7][0][110],
F_[7][1][110],
F_[7][2][110],
F_[8][0][110],
F_[8][1][110],
F_[8][2][110],
F_[9][0][110],
F_[9][1][110],
F_[9][2][110],
F_[10][0][110],
F_[10][1][110],
F_[10][2][110],
F_[11][0][110],
F_[11][1][110],
F_[11][2][110],
F_[12][0][110],
F_[12][1][110],
F_[12][2][110],
F_[13][0][110],
F_[13][1][110],
F_[13][2][110],
F_[14][0][110],
F_[14][1][110],
F_[14][2][110],
F_[15][0][110],
F_[15][1][110],
F_[15][2][110],
F_[0][0][111],
F_[0][1][111],
F_[0][2][111],
F_[1][0][111],
F_[1][1][111],
F_[1][2][111],
F_[2][0][111],
F_[2][1][111],
F_[2][2][111],
F_[3][0][111],
F_[3][1][111],
F_[3][2][111],
F_[4][0][111],
F_[4][1][111],
F_[4][2][111],
F_[5][0][111],
F_[5][1][111],
F_[5][2][111],
F_[6][0][111],
F_[6][1][111],
F_[6][2][111],
F_[7][0][111],
F_[7][1][111],
F_[7][2][111],
F_[8][0][111],
F_[8][1][111],
F_[8][2][111],
F_[9][0][111],
F_[9][1][111],
F_[9][2][111],
F_[10][0][111],
F_[10][1][111],
F_[10][2][111],
F_[11][0][111],
F_[11][1][111],
F_[11][2][111],
F_[12][0][111],
F_[12][1][111],
F_[12][2][111],
F_[13][0][111],
F_[13][1][111],
F_[13][2][111],
F_[14][0][111],
F_[14][1][111],
F_[14][2][111],
F_[15][0][111],
F_[15][1][111],
F_[15][2][111],
F_[0][0][112],
F_[0][1][112],
F_[0][2][112],
F_[1][0][112],
F_[1][1][112],
F_[1][2][112],
F_[2][0][112],
F_[2][1][112],
F_[2][2][112],
F_[3][0][112],
F_[3][1][112],
F_[3][2][112],
F_[4][0][112],
F_[4][1][112],
F_[4][2][112],
F_[5][0][112],
F_[5][1][112],
F_[5][2][112],
F_[6][0][112],
F_[6][1][112],
F_[6][2][112],
F_[7][0][112],
F_[7][1][112],
F_[7][2][112],
F_[8][0][112],
F_[8][1][112],
F_[8][2][112],
F_[9][0][112],
F_[9][1][112],
F_[9][2][112],
F_[10][0][112],
F_[10][1][112],
F_[10][2][112],
F_[11][0][112],
F_[11][1][112],
F_[11][2][112],
F_[12][0][112],
F_[12][1][112],
F_[12][2][112],
F_[13][0][112],
F_[13][1][112],
F_[13][2][112],
F_[14][0][112],
F_[14][1][112],
F_[14][2][112],
F_[15][0][112],
F_[15][1][112],
F_[15][2][112],
F_[0][0][113],
F_[0][1][113],
F_[0][2][113],
F_[1][0][113],
F_[1][1][113],
F_[1][2][113],
F_[2][0][113],
F_[2][1][113],
F_[2][2][113],
F_[3][0][113],
F_[3][1][113],
F_[3][2][113],
F_[4][0][113],
F_[4][1][113],
F_[4][2][113],
F_[5][0][113],
F_[5][1][113],
F_[5][2][113],
F_[6][0][113],
F_[6][1][113],
F_[6][2][113],
F_[7][0][113],
F_[7][1][113],
F_[7][2][113],
F_[8][0][113],
F_[8][1][113],
F_[8][2][113],
F_[9][0][113],
F_[9][1][113],
F_[9][2][113],
F_[10][0][113],
F_[10][1][113],
F_[10][2][113],
F_[11][0][113],
F_[11][1][113],
F_[11][2][113],
F_[12][0][113],
F_[12][1][113],
F_[12][2][113],
F_[13][0][113],
F_[13][1][113],
F_[13][2][113],
F_[14][0][113],
F_[14][1][113],
F_[14][2][113],
F_[15][0][113],
F_[15][1][113],
F_[15][2][113],
F_[0][0][114],
F_[0][1][114],
F_[0][2][114],
F_[1][0][114],
F_[1][1][114],
F_[1][2][114],
F_[2][0][114],
F_[2][1][114],
F_[2][2][114],
F_[3][0][114],
F_[3][1][114],
F_[3][2][114],
F_[4][0][114],
F_[4][1][114],
F_[4][2][114],
F_[5][0][114],
F_[5][1][114],
F_[5][2][114],
F_[6][0][114],
F_[6][1][114],
F_[6][2][114],
F_[7][0][114],
F_[7][1][114],
F_[7][2][114],
F_[8][0][114],
F_[8][1][114],
F_[8][2][114],
F_[9][0][114],
F_[9][1][114],
F_[9][2][114],
F_[10][0][114],
F_[10][1][114],
F_[10][2][114],
F_[11][0][114],
F_[11][1][114],
F_[11][2][114],
F_[12][0][114],
F_[12][1][114],
F_[12][2][114],
F_[13][0][114],
F_[13][1][114],
F_[13][2][114],
F_[14][0][114],
F_[14][1][114],
F_[14][2][114],
F_[15][0][114],
F_[15][1][114],
F_[15][2][114],
F_[0][0][115],
F_[0][1][115],
F_[0][2][115],
F_[1][0][115],
F_[1][1][115],
F_[1][2][115],
F_[2][0][115],
F_[2][1][115],
F_[2][2][115],
F_[3][0][115],
F_[3][1][115],
F_[3][2][115],
F_[4][0][115],
F_[4][1][115],
F_[4][2][115],
F_[5][0][115],
F_[5][1][115],
F_[5][2][115],
F_[6][0][115],
F_[6][1][115],
F_[6][2][115],
F_[7][0][115],
F_[7][1][115],
F_[7][2][115],
F_[8][0][115],
F_[8][1][115],
F_[8][2][115],
F_[9][0][115],
F_[9][1][115],
F_[9][2][115],
F_[10][0][115],
F_[10][1][115],
F_[10][2][115],
F_[11][0][115],
F_[11][1][115],
F_[11][2][115],
F_[12][0][115],
F_[12][1][115],
F_[12][2][115],
F_[13][0][115],
F_[13][1][115],
F_[13][2][115],
F_[14][0][115],
F_[14][1][115],
F_[14][2][115],
F_[15][0][115],
F_[15][1][115],
F_[15][2][115],
F_[0][0][116],
F_[0][1][116],
F_[0][2][116],
F_[1][0][116],
F_[1][1][116],
F_[1][2][116],
F_[2][0][116],
F_[2][1][116],
F_[2][2][116],
F_[3][0][116],
F_[3][1][116],
F_[3][2][116],
F_[4][0][116],
F_[4][1][116],
F_[4][2][116],
F_[5][0][116],
F_[5][1][116],
F_[5][2][116],
F_[6][0][116],
F_[6][1][116],
F_[6][2][116],
F_[7][0][116],
F_[7][1][116],
F_[7][2][116],
F_[8][0][116],
F_[8][1][116],
F_[8][2][116],
F_[9][0][116],
F_[9][1][116],
F_[9][2][116],
F_[10][0][116],
F_[10][1][116],
F_[10][2][116],
F_[11][0][116],
F_[11][1][116],
F_[11][2][116],
F_[12][0][116],
F_[12][1][116],
F_[12][2][116],
F_[13][0][116],
F_[13][1][116],
F_[13][2][116],
F_[14][0][116],
F_[14][1][116],
F_[14][2][116],
F_[15][0][116],
F_[15][1][116],
F_[15][2][116],
F_[0][0][117],
F_[0][1][117],
F_[0][2][117],
F_[1][0][117],
F_[1][1][117],
F_[1][2][117],
F_[2][0][117],
F_[2][1][117],
F_[2][2][117],
F_[3][0][117],
F_[3][1][117],
F_[3][2][117],
F_[4][0][117],
F_[4][1][117],
F_[4][2][117],
F_[5][0][117],
F_[5][1][117],
F_[5][2][117],
F_[6][0][117],
F_[6][1][117],
F_[6][2][117],
F_[7][0][117],
F_[7][1][117],
F_[7][2][117],
F_[8][0][117],
F_[8][1][117],
F_[8][2][117],
F_[9][0][117],
F_[9][1][117],
F_[9][2][117],
F_[10][0][117],
F_[10][1][117],
F_[10][2][117],
F_[11][0][117],
F_[11][1][117],
F_[11][2][117],
F_[12][0][117],
F_[12][1][117],
F_[12][2][117],
F_[13][0][117],
F_[13][1][117],
F_[13][2][117],
F_[14][0][117],
F_[14][1][117],
F_[14][2][117],
F_[15][0][117],
F_[15][1][117],
F_[15][2][117],
F_[0][0][118],
F_[0][1][118],
F_[0][2][118],
F_[1][0][118],
F_[1][1][118],
F_[1][2][118],
F_[2][0][118],
F_[2][1][118],
F_[2][2][118],
F_[3][0][118],
F_[3][1][118],
F_[3][2][118],
F_[4][0][118],
F_[4][1][118],
F_[4][2][118],
F_[5][0][118],
F_[5][1][118],
F_[5][2][118],
F_[6][0][118],
F_[6][1][118],
F_[6][2][118],
F_[7][0][118],
F_[7][1][118],
F_[7][2][118],
F_[8][0][118],
F_[8][1][118],
F_[8][2][118],
F_[9][0][118],
F_[9][1][118],
F_[9][2][118],
F_[10][0][118],
F_[10][1][118],
F_[10][2][118],
F_[11][0][118],
F_[11][1][118],
F_[11][2][118],
F_[12][0][118],
F_[12][1][118],
F_[12][2][118],
F_[13][0][118],
F_[13][1][118],
F_[13][2][118],
F_[14][0][118],
F_[14][1][118],
F_[14][2][118],
F_[15][0][118],
F_[15][1][118],
F_[15][2][118],
F_[0][0][119],
F_[0][1][119],
F_[0][2][119],
F_[1][0][119],
F_[1][1][119],
F_[1][2][119],
F_[2][0][119],
F_[2][1][119],
F_[2][2][119],
F_[3][0][119],
F_[3][1][119],
F_[3][2][119],
F_[4][0][119],
F_[4][1][119],
F_[4][2][119],
F_[5][0][119],
F_[5][1][119],
F_[5][2][119],
F_[6][0][119],
F_[6][1][119],
F_[6][2][119],
F_[7][0][119],
F_[7][1][119],
F_[7][2][119],
F_[8][0][119],
F_[8][1][119],
F_[8][2][119],
F_[9][0][119],
F_[9][1][119],
F_[9][2][119],
F_[10][0][119],
F_[10][1][119],
F_[10][2][119],
F_[11][0][119],
F_[11][1][119],
F_[11][2][119],
F_[12][0][119],
F_[12][1][119],
F_[12][2][119],
F_[13][0][119],
F_[13][1][119],
F_[13][2][119],
F_[14][0][119],
F_[14][1][119],
F_[14][2][119],
F_[15][0][119],
F_[15][1][119],
F_[15][2][119],
F_[0][0][120],
F_[0][1][120],
F_[0][2][120],
F_[1][0][120],
F_[1][1][120],
F_[1][2][120],
F_[2][0][120],
F_[2][1][120],
F_[2][2][120],
F_[3][0][120],
F_[3][1][120],
F_[3][2][120],
F_[4][0][120],
F_[4][1][120],
F_[4][2][120],
F_[5][0][120],
F_[5][1][120],
F_[5][2][120],
F_[6][0][120],
F_[6][1][120],
F_[6][2][120],
F_[7][0][120],
F_[7][1][120],
F_[7][2][120],
F_[8][0][120],
F_[8][1][120],
F_[8][2][120],
F_[9][0][120],
F_[9][1][120],
F_[9][2][120],
F_[10][0][120],
F_[10][1][120],
F_[10][2][120],
F_[11][0][120],
F_[11][1][120],
F_[11][2][120],
F_[12][0][120],
F_[12][1][120],
F_[12][2][120],
F_[13][0][120],
F_[13][1][120],
F_[13][2][120],
F_[14][0][120],
F_[14][1][120],
F_[14][2][120],
F_[15][0][120],
F_[15][1][120],
F_[15][2][120],
F_[0][0][121],
F_[0][1][121],
F_[0][2][121],
F_[1][0][121],
F_[1][1][121],
F_[1][2][121],
F_[2][0][121],
F_[2][1][121],
F_[2][2][121],
F_[3][0][121],
F_[3][1][121],
F_[3][2][121],
F_[4][0][121],
F_[4][1][121],
F_[4][2][121],
F_[5][0][121],
F_[5][1][121],
F_[5][2][121],
F_[6][0][121],
F_[6][1][121],
F_[6][2][121],
F_[7][0][121],
F_[7][1][121],
F_[7][2][121],
F_[8][0][121],
F_[8][1][121],
F_[8][2][121],
F_[9][0][121],
F_[9][1][121],
F_[9][2][121],
F_[10][0][121],
F_[10][1][121],
F_[10][2][121],
F_[11][0][121],
F_[11][1][121],
F_[11][2][121],
F_[12][0][121],
F_[12][1][121],
F_[12][2][121],
F_[13][0][121],
F_[13][1][121],
F_[13][2][121],
F_[14][0][121],
F_[14][1][121],
F_[14][2][121],
F_[15][0][121],
F_[15][1][121],
F_[15][2][121],
F_[0][0][122],
F_[0][1][122],
F_[0][2][122],
F_[1][0][122],
F_[1][1][122],
F_[1][2][122],
F_[2][0][122],
F_[2][1][122],
F_[2][2][122],
F_[3][0][122],
F_[3][1][122],
F_[3][2][122],
F_[4][0][122],
F_[4][1][122],
F_[4][2][122],
F_[5][0][122],
F_[5][1][122],
F_[5][2][122],
F_[6][0][122],
F_[6][1][122],
F_[6][2][122],
F_[7][0][122],
F_[7][1][122],
F_[7][2][122],
F_[8][0][122],
F_[8][1][122],
F_[8][2][122],
F_[9][0][122],
F_[9][1][122],
F_[9][2][122],
F_[10][0][122],
F_[10][1][122],
F_[10][2][122],
F_[11][0][122],
F_[11][1][122],
F_[11][2][122],
F_[12][0][122],
F_[12][1][122],
F_[12][2][122],
F_[13][0][122],
F_[13][1][122],
F_[13][2][122],
F_[14][0][122],
F_[14][1][122],
F_[14][2][122],
F_[15][0][122],
F_[15][1][122],
F_[15][2][122],
F_[0][0][123],
F_[0][1][123],
F_[0][2][123],
F_[1][0][123],
F_[1][1][123],
F_[1][2][123],
F_[2][0][123],
F_[2][1][123],
F_[2][2][123],
F_[3][0][123],
F_[3][1][123],
F_[3][2][123],
F_[4][0][123],
F_[4][1][123],
F_[4][2][123],
F_[5][0][123],
F_[5][1][123],
F_[5][2][123],
F_[6][0][123],
F_[6][1][123],
F_[6][2][123],
F_[7][0][123],
F_[7][1][123],
F_[7][2][123],
F_[8][0][123],
F_[8][1][123],
F_[8][2][123],
F_[9][0][123],
F_[9][1][123],
F_[9][2][123],
F_[10][0][123],
F_[10][1][123],
F_[10][2][123],
F_[11][0][123],
F_[11][1][123],
F_[11][2][123],
F_[12][0][123],
F_[12][1][123],
F_[12][2][123],
F_[13][0][123],
F_[13][1][123],
F_[13][2][123],
F_[14][0][123],
F_[14][1][123],
F_[14][2][123],
F_[15][0][123],
F_[15][1][123],
F_[15][2][123],
F_[0][0][124],
F_[0][1][124],
F_[0][2][124],
F_[1][0][124],
F_[1][1][124],
F_[1][2][124],
F_[2][0][124],
F_[2][1][124],
F_[2][2][124],
F_[3][0][124],
F_[3][1][124],
F_[3][2][124],
F_[4][0][124],
F_[4][1][124],
F_[4][2][124],
F_[5][0][124],
F_[5][1][124],
F_[5][2][124],
F_[6][0][124],
F_[6][1][124],
F_[6][2][124],
F_[7][0][124],
F_[7][1][124],
F_[7][2][124],
F_[8][0][124],
F_[8][1][124],
F_[8][2][124],
F_[9][0][124],
F_[9][1][124],
F_[9][2][124],
F_[10][0][124],
F_[10][1][124],
F_[10][2][124],
F_[11][0][124],
F_[11][1][124],
F_[11][2][124],
F_[12][0][124],
F_[12][1][124],
F_[12][2][124],
F_[13][0][124],
F_[13][1][124],
F_[13][2][124],
F_[14][0][124],
F_[14][1][124],
F_[14][2][124],
F_[15][0][124],
F_[15][1][124],
F_[15][2][124],
F_[0][0][125],
F_[0][1][125],
F_[0][2][125],
F_[1][0][125],
F_[1][1][125],
F_[1][2][125],
F_[2][0][125],
F_[2][1][125],
F_[2][2][125],
F_[3][0][125],
F_[3][1][125],
F_[3][2][125],
F_[4][0][125],
F_[4][1][125],
F_[4][2][125],
F_[5][0][125],
F_[5][1][125],
F_[5][2][125],
F_[6][0][125],
F_[6][1][125],
F_[6][2][125],
F_[7][0][125],
F_[7][1][125],
F_[7][2][125],
F_[8][0][125],
F_[8][1][125],
F_[8][2][125],
F_[9][0][125],
F_[9][1][125],
F_[9][2][125],
F_[10][0][125],
F_[10][1][125],
F_[10][2][125],
F_[11][0][125],
F_[11][1][125],
F_[11][2][125],
F_[12][0][125],
F_[12][1][125],
F_[12][2][125],
F_[13][0][125],
F_[13][1][125],
F_[13][2][125],
F_[14][0][125],
F_[14][1][125],
F_[14][2][125],
F_[15][0][125],
F_[15][1][125],
F_[15][2][125],
F_[0][0][126],
F_[0][1][126],
F_[0][2][126],
F_[1][0][126],
F_[1][1][126],
F_[1][2][126],
F_[2][0][126],
F_[2][1][126],
F_[2][2][126],
F_[3][0][126],
F_[3][1][126],
F_[3][2][126],
F_[4][0][126],
F_[4][1][126],
F_[4][2][126],
F_[5][0][126],
F_[5][1][126],
F_[5][2][126],
F_[6][0][126],
F_[6][1][126],
F_[6][2][126],
F_[7][0][126],
F_[7][1][126],
F_[7][2][126],
F_[8][0][126],
F_[8][1][126],
F_[8][2][126],
F_[9][0][126],
F_[9][1][126],
F_[9][2][126],
F_[10][0][126],
F_[10][1][126],
F_[10][2][126],
F_[11][0][126],
F_[11][1][126],
F_[11][2][126],
F_[12][0][126],
F_[12][1][126],
F_[12][2][126],
F_[13][0][126],
F_[13][1][126],
F_[13][2][126],
F_[14][0][126],
F_[14][1][126],
F_[14][2][126],
F_[15][0][126],
F_[15][1][126],
F_[15][2][126],
F_[0][0][127],
F_[0][1][127],
F_[0][2][127],
F_[1][0][127],
F_[1][1][127],
F_[1][2][127],
F_[2][0][127],
F_[2][1][127],
F_[2][2][127],
F_[3][0][127],
F_[3][1][127],
F_[3][2][127],
F_[4][0][127],
F_[4][1][127],
F_[4][2][127],
F_[5][0][127],
F_[5][1][127],
F_[5][2][127],
F_[6][0][127],
F_[6][1][127],
F_[6][2][127],
F_[7][0][127],
F_[7][1][127],
F_[7][2][127],
F_[8][0][127],
F_[8][1][127],
F_[8][2][127],
F_[9][0][127],
F_[9][1][127],
F_[9][2][127],
F_[10][0][127],
F_[10][1][127],
F_[10][2][127],
F_[11][0][127],
F_[11][1][127],
F_[11][2][127],
F_[12][0][127],
F_[12][1][127],
F_[12][2][127],
F_[13][0][127],
F_[13][1][127],
F_[13][2][127],
F_[14][0][127],
F_[14][1][127],
F_[14][2][127],
F_[15][0][127],
F_[15][1][127],
F_[15][2][127],
F_[0][0][128],
F_[0][1][128],
F_[0][2][128],
F_[1][0][128],
F_[1][1][128],
F_[1][2][128],
F_[2][0][128],
F_[2][1][128],
F_[2][2][128],
F_[3][0][128],
F_[3][1][128],
F_[3][2][128],
F_[4][0][128],
F_[4][1][128],
F_[4][2][128],
F_[5][0][128],
F_[5][1][128],
F_[5][2][128],
F_[6][0][128],
F_[6][1][128],
F_[6][2][128],
F_[7][0][128],
F_[7][1][128],
F_[7][2][128],
F_[8][0][128],
F_[8][1][128],
F_[8][2][128],
F_[9][0][128],
F_[9][1][128],
F_[9][2][128],
F_[10][0][128],
F_[10][1][128],
F_[10][2][128],
F_[11][0][128],
F_[11][1][128],
F_[11][2][128],
F_[12][0][128],
F_[12][1][128],
F_[12][2][128],
F_[13][0][128],
F_[13][1][128],
F_[13][2][128],
F_[14][0][128],
F_[14][1][128],
F_[14][2][128],
F_[15][0][128],
F_[15][1][128],
F_[15][2][128],
F_[0][0][129],
F_[0][1][129],
F_[0][2][129],
F_[1][0][129],
F_[1][1][129],
F_[1][2][129],
F_[2][0][129],
F_[2][1][129],
F_[2][2][129],
F_[3][0][129],
F_[3][1][129],
F_[3][2][129],
F_[4][0][129],
F_[4][1][129],
F_[4][2][129],
F_[5][0][129],
F_[5][1][129],
F_[5][2][129],
F_[6][0][129],
F_[6][1][129],
F_[6][2][129],
F_[7][0][129],
F_[7][1][129],
F_[7][2][129],
F_[8][0][129],
F_[8][1][129],
F_[8][2][129],
F_[9][0][129],
F_[9][1][129],
F_[9][2][129],
F_[10][0][129],
F_[10][1][129],
F_[10][2][129],
F_[11][0][129],
F_[11][1][129],
F_[11][2][129],
F_[12][0][129],
F_[12][1][129],
F_[12][2][129],
F_[13][0][129],
F_[13][1][129],
F_[13][2][129],
F_[14][0][129],
F_[14][1][129],
F_[14][2][129],
F_[15][0][129],
F_[15][1][129],
F_[15][2][129],
F_[0][0][130],
F_[0][1][130],
F_[0][2][130],
F_[1][0][130],
F_[1][1][130],
F_[1][2][130],
F_[2][0][130],
F_[2][1][130],
F_[2][2][130],
F_[3][0][130],
F_[3][1][130],
F_[3][2][130],
F_[4][0][130],
F_[4][1][130],
F_[4][2][130],
F_[5][0][130],
F_[5][1][130],
F_[5][2][130],
F_[6][0][130],
F_[6][1][130],
F_[6][2][130],
F_[7][0][130],
F_[7][1][130],
F_[7][2][130],
F_[8][0][130],
F_[8][1][130],
F_[8][2][130],
F_[9][0][130],
F_[9][1][130],
F_[9][2][130],
F_[10][0][130],
F_[10][1][130],
F_[10][2][130],
F_[11][0][130],
F_[11][1][130],
F_[11][2][130],
F_[12][0][130],
F_[12][1][130],
F_[12][2][130],
F_[13][0][130],
F_[13][1][130],
F_[13][2][130],
F_[14][0][130],
F_[14][1][130],
F_[14][2][130],
F_[15][0][130],
F_[15][1][130],
F_[15][2][130],
F_[0][0][131],
F_[0][1][131],
F_[0][2][131],
F_[1][0][131],
F_[1][1][131],
F_[1][2][131],
F_[2][0][131],
F_[2][1][131],
F_[2][2][131],
F_[3][0][131],
F_[3][1][131],
F_[3][2][131],
F_[4][0][131],
F_[4][1][131],
F_[4][2][131],
F_[5][0][131],
F_[5][1][131],
F_[5][2][131],
F_[6][0][131],
F_[6][1][131],
F_[6][2][131],
F_[7][0][131],
F_[7][1][131],
F_[7][2][131],
F_[8][0][131],
F_[8][1][131],
F_[8][2][131],
F_[9][0][131],
F_[9][1][131],
F_[9][2][131],
F_[10][0][131],
F_[10][1][131],
F_[10][2][131],
F_[11][0][131],
F_[11][1][131],
F_[11][2][131],
F_[12][0][131],
F_[12][1][131],
F_[12][2][131],
F_[13][0][131],
F_[13][1][131],
F_[13][2][131],
F_[14][0][131],
F_[14][1][131],
F_[14][2][131],
F_[15][0][131],
F_[15][1][131],
F_[15][2][131],
F_[0][0][132],
F_[0][1][132],
F_[0][2][132],
F_[1][0][132],
F_[1][1][132],
F_[1][2][132],
F_[2][0][132],
F_[2][1][132],
F_[2][2][132],
F_[3][0][132],
F_[3][1][132],
F_[3][2][132],
F_[4][0][132],
F_[4][1][132],
F_[4][2][132],
F_[5][0][132],
F_[5][1][132],
F_[5][2][132],
F_[6][0][132],
F_[6][1][132],
F_[6][2][132],
F_[7][0][132],
F_[7][1][132],
F_[7][2][132],
F_[8][0][132],
F_[8][1][132],
F_[8][2][132],
F_[9][0][132],
F_[9][1][132],
F_[9][2][132],
F_[10][0][132],
F_[10][1][132],
F_[10][2][132],
F_[11][0][132],
F_[11][1][132],
F_[11][2][132],
F_[12][0][132],
F_[12][1][132],
F_[12][2][132],
F_[13][0][132],
F_[13][1][132],
F_[13][2][132],
F_[14][0][132],
F_[14][1][132],
F_[14][2][132],
F_[15][0][132],
F_[15][1][132],
F_[15][2][132],
F_[0][0][133],
F_[0][1][133],
F_[0][2][133],
F_[1][0][133],
F_[1][1][133],
F_[1][2][133],
F_[2][0][133],
F_[2][1][133],
F_[2][2][133],
F_[3][0][133],
F_[3][1][133],
F_[3][2][133],
F_[4][0][133],
F_[4][1][133],
F_[4][2][133],
F_[5][0][133],
F_[5][1][133],
F_[5][2][133],
F_[6][0][133],
F_[6][1][133],
F_[6][2][133],
F_[7][0][133],
F_[7][1][133],
F_[7][2][133],
F_[8][0][133],
F_[8][1][133],
F_[8][2][133],
F_[9][0][133],
F_[9][1][133],
F_[9][2][133],
F_[10][0][133],
F_[10][1][133],
F_[10][2][133],
F_[11][0][133],
F_[11][1][133],
F_[11][2][133],
F_[12][0][133],
F_[12][1][133],
F_[12][2][133],
F_[13][0][133],
F_[13][1][133],
F_[13][2][133],
F_[14][0][133],
F_[14][1][133],
F_[14][2][133],
F_[15][0][133],
F_[15][1][133],
F_[15][2][133],
F_[0][0][134],
F_[0][1][134],
F_[0][2][134],
F_[1][0][134],
F_[1][1][134],
F_[1][2][134],
F_[2][0][134],
F_[2][1][134],
F_[2][2][134],
F_[3][0][134],
F_[3][1][134],
F_[3][2][134],
F_[4][0][134],
F_[4][1][134],
F_[4][2][134],
F_[5][0][134],
F_[5][1][134],
F_[5][2][134],
F_[6][0][134],
F_[6][1][134],
F_[6][2][134],
F_[7][0][134],
F_[7][1][134],
F_[7][2][134],
F_[8][0][134],
F_[8][1][134],
F_[8][2][134],
F_[9][0][134],
F_[9][1][134],
F_[9][2][134],
F_[10][0][134],
F_[10][1][134],
F_[10][2][134],
F_[11][0][134],
F_[11][1][134],
F_[11][2][134],
F_[12][0][134],
F_[12][1][134],
F_[12][2][134],
F_[13][0][134],
F_[13][1][134],
F_[13][2][134],
F_[14][0][134],
F_[14][1][134],
F_[14][2][134],
F_[15][0][134],
F_[15][1][134],
F_[15][2][134],
F_[0][0][135],
F_[0][1][135],
F_[0][2][135],
F_[1][0][135],
F_[1][1][135],
F_[1][2][135],
F_[2][0][135],
F_[2][1][135],
F_[2][2][135],
F_[3][0][135],
F_[3][1][135],
F_[3][2][135],
F_[4][0][135],
F_[4][1][135],
F_[4][2][135],
F_[5][0][135],
F_[5][1][135],
F_[5][2][135],
F_[6][0][135],
F_[6][1][135],
F_[6][2][135],
F_[7][0][135],
F_[7][1][135],
F_[7][2][135],
F_[8][0][135],
F_[8][1][135],
F_[8][2][135],
F_[9][0][135],
F_[9][1][135],
F_[9][2][135],
F_[10][0][135],
F_[10][1][135],
F_[10][2][135],
F_[11][0][135],
F_[11][1][135],
F_[11][2][135],
F_[12][0][135],
F_[12][1][135],
F_[12][2][135],
F_[13][0][135],
F_[13][1][135],
F_[13][2][135],
F_[14][0][135],
F_[14][1][135],
F_[14][2][135],
F_[15][0][135],
F_[15][1][135],
F_[15][2][135],
F_[0][0][136],
F_[0][1][136],
F_[0][2][136],
F_[1][0][136],
F_[1][1][136],
F_[1][2][136],
F_[2][0][136],
F_[2][1][136],
F_[2][2][136],
F_[3][0][136],
F_[3][1][136],
F_[3][2][136],
F_[4][0][136],
F_[4][1][136],
F_[4][2][136],
F_[5][0][136],
F_[5][1][136],
F_[5][2][136],
F_[6][0][136],
F_[6][1][136],
F_[6][2][136],
F_[7][0][136],
F_[7][1][136],
F_[7][2][136],
F_[8][0][136],
F_[8][1][136],
F_[8][2][136],
F_[9][0][136],
F_[9][1][136],
F_[9][2][136],
F_[10][0][136],
F_[10][1][136],
F_[10][2][136],
F_[11][0][136],
F_[11][1][136],
F_[11][2][136],
F_[12][0][136],
F_[12][1][136],
F_[12][2][136],
F_[13][0][136],
F_[13][1][136],
F_[13][2][136],
F_[14][0][136],
F_[14][1][136],
F_[14][2][136],
F_[15][0][136],
F_[15][1][136],
F_[15][2][136],
F_[0][0][137],
F_[0][1][137],
F_[0][2][137],
F_[1][0][137],
F_[1][1][137],
F_[1][2][137],
F_[2][0][137],
F_[2][1][137],
F_[2][2][137],
F_[3][0][137],
F_[3][1][137],
F_[3][2][137],
F_[4][0][137],
F_[4][1][137],
F_[4][2][137],
F_[5][0][137],
F_[5][1][137],
F_[5][2][137],
F_[6][0][137],
F_[6][1][137],
F_[6][2][137],
F_[7][0][137],
F_[7][1][137],
F_[7][2][137],
F_[8][0][137],
F_[8][1][137],
F_[8][2][137],
F_[9][0][137],
F_[9][1][137],
F_[9][2][137],
F_[10][0][137],
F_[10][1][137],
F_[10][2][137],
F_[11][0][137],
F_[11][1][137],
F_[11][2][137],
F_[12][0][137],
F_[12][1][137],
F_[12][2][137],
F_[13][0][137],
F_[13][1][137],
F_[13][2][137],
F_[14][0][137],
F_[14][1][137],
F_[14][2][137],
F_[15][0][137],
F_[15][1][137],
F_[15][2][137],
F_[0][0][138],
F_[0][1][138],
F_[0][2][138],
F_[1][0][138],
F_[1][1][138],
F_[1][2][138],
F_[2][0][138],
F_[2][1][138],
F_[2][2][138],
F_[3][0][138],
F_[3][1][138],
F_[3][2][138],
F_[4][0][138],
F_[4][1][138],
F_[4][2][138],
F_[5][0][138],
F_[5][1][138],
F_[5][2][138],
F_[6][0][138],
F_[6][1][138],
F_[6][2][138],
F_[7][0][138],
F_[7][1][138],
F_[7][2][138],
F_[8][0][138],
F_[8][1][138],
F_[8][2][138],
F_[9][0][138],
F_[9][1][138],
F_[9][2][138],
F_[10][0][138],
F_[10][1][138],
F_[10][2][138],
F_[11][0][138],
F_[11][1][138],
F_[11][2][138],
F_[12][0][138],
F_[12][1][138],
F_[12][2][138],
F_[13][0][138],
F_[13][1][138],
F_[13][2][138],
F_[14][0][138],
F_[14][1][138],
F_[14][2][138],
F_[15][0][138],
F_[15][1][138],
F_[15][2][138],
F_[0][0][139],
F_[0][1][139],
F_[0][2][139],
F_[1][0][139],
F_[1][1][139],
F_[1][2][139],
F_[2][0][139],
F_[2][1][139],
F_[2][2][139],
F_[3][0][139],
F_[3][1][139],
F_[3][2][139],
F_[4][0][139],
F_[4][1][139],
F_[4][2][139],
F_[5][0][139],
F_[5][1][139],
F_[5][2][139],
F_[6][0][139],
F_[6][1][139],
F_[6][2][139],
F_[7][0][139],
F_[7][1][139],
F_[7][2][139],
F_[8][0][139],
F_[8][1][139],
F_[8][2][139],
F_[9][0][139],
F_[9][1][139],
F_[9][2][139],
F_[10][0][139],
F_[10][1][139],
F_[10][2][139],
F_[11][0][139],
F_[11][1][139],
F_[11][2][139],
F_[12][0][139],
F_[12][1][139],
F_[12][2][139],
F_[13][0][139],
F_[13][1][139],
F_[13][2][139],
F_[14][0][139],
F_[14][1][139],
F_[14][2][139],
F_[15][0][139],
F_[15][1][139],
F_[15][2][139],
F_[0][0][140],
F_[0][1][140],
F_[0][2][140],
F_[1][0][140],
F_[1][1][140],
F_[1][2][140],
F_[2][0][140],
F_[2][1][140],
F_[2][2][140],
F_[3][0][140],
F_[3][1][140],
F_[3][2][140],
F_[4][0][140],
F_[4][1][140],
F_[4][2][140],
F_[5][0][140],
F_[5][1][140],
F_[5][2][140],
F_[6][0][140],
F_[6][1][140],
F_[6][2][140],
F_[7][0][140],
F_[7][1][140],
F_[7][2][140],
F_[8][0][140],
F_[8][1][140],
F_[8][2][140],
F_[9][0][140],
F_[9][1][140],
F_[9][2][140],
F_[10][0][140],
F_[10][1][140],
F_[10][2][140],
F_[11][0][140],
F_[11][1][140],
F_[11][2][140],
F_[12][0][140],
F_[12][1][140],
F_[12][2][140],
F_[13][0][140],
F_[13][1][140],
F_[13][2][140],
F_[14][0][140],
F_[14][1][140],
F_[14][2][140],
F_[15][0][140],
F_[15][1][140],
F_[15][2][140],
F_[0][0][141],
F_[0][1][141],
F_[0][2][141],
F_[1][0][141],
F_[1][1][141],
F_[1][2][141],
F_[2][0][141],
F_[2][1][141],
F_[2][2][141],
F_[3][0][141],
F_[3][1][141],
F_[3][2][141],
F_[4][0][141],
F_[4][1][141],
F_[4][2][141],
F_[5][0][141],
F_[5][1][141],
F_[5][2][141],
F_[6][0][141],
F_[6][1][141],
F_[6][2][141],
F_[7][0][141],
F_[7][1][141],
F_[7][2][141],
F_[8][0][141],
F_[8][1][141],
F_[8][2][141],
F_[9][0][141],
F_[9][1][141],
F_[9][2][141],
F_[10][0][141],
F_[10][1][141],
F_[10][2][141],
F_[11][0][141],
F_[11][1][141],
F_[11][2][141],
F_[12][0][141],
F_[12][1][141],
F_[12][2][141],
F_[13][0][141],
F_[13][1][141],
F_[13][2][141],
F_[14][0][141],
F_[14][1][141],
F_[14][2][141],
F_[15][0][141],
F_[15][1][141],
F_[15][2][141],
F_[0][0][142],
F_[0][1][142],
F_[0][2][142],
F_[1][0][142],
F_[1][1][142],
F_[1][2][142],
F_[2][0][142],
F_[2][1][142],
F_[2][2][142],
F_[3][0][142],
F_[3][1][142],
F_[3][2][142],
F_[4][0][142],
F_[4][1][142],
F_[4][2][142],
F_[5][0][142],
F_[5][1][142],
F_[5][2][142],
F_[6][0][142],
F_[6][1][142],
F_[6][2][142],
F_[7][0][142],
F_[7][1][142],
F_[7][2][142],
F_[8][0][142],
F_[8][1][142],
F_[8][2][142],
F_[9][0][142],
F_[9][1][142],
F_[9][2][142],
F_[10][0][142],
F_[10][1][142],
F_[10][2][142],
F_[11][0][142],
F_[11][1][142],
F_[11][2][142],
F_[12][0][142],
F_[12][1][142],
F_[12][2][142],
F_[13][0][142],
F_[13][1][142],
F_[13][2][142],
F_[14][0][142],
F_[14][1][142],
F_[14][2][142],
F_[15][0][142],
F_[15][1][142],
F_[15][2][142],
F_[0][0][143],
F_[0][1][143],
F_[0][2][143],
F_[1][0][143],
F_[1][1][143],
F_[1][2][143],
F_[2][0][143],
F_[2][1][143],
F_[2][2][143],
F_[3][0][143],
F_[3][1][143],
F_[3][2][143],
F_[4][0][143],
F_[4][1][143],
F_[4][2][143],
F_[5][0][143],
F_[5][1][143],
F_[5][2][143],
F_[6][0][143],
F_[6][1][143],
F_[6][2][143],
F_[7][0][143],
F_[7][1][143],
F_[7][2][143],
F_[8][0][143],
F_[8][1][143],
F_[8][2][143],
F_[9][0][143],
F_[9][1][143],
F_[9][2][143],
F_[10][0][143],
F_[10][1][143],
F_[10][2][143],
F_[11][0][143],
F_[11][1][143],
F_[11][2][143],
F_[12][0][143],
F_[12][1][143],
F_[12][2][143],
F_[13][0][143],
F_[13][1][143],
F_[13][2][143],
F_[14][0][143],
F_[14][1][143],
F_[14][2][143],
F_[15][0][143],
F_[15][1][143],
F_[15][2][143],
F_[0][0][144],
F_[0][1][144],
F_[0][2][144],
F_[1][0][144],
F_[1][1][144],
F_[1][2][144],
F_[2][0][144],
F_[2][1][144],
F_[2][2][144],
F_[3][0][144],
F_[3][1][144],
F_[3][2][144],
F_[4][0][144],
F_[4][1][144],
F_[4][2][144],
F_[5][0][144],
F_[5][1][144],
F_[5][2][144],
F_[6][0][144],
F_[6][1][144],
F_[6][2][144],
F_[7][0][144],
F_[7][1][144],
F_[7][2][144],
F_[8][0][144],
F_[8][1][144],
F_[8][2][144],
F_[9][0][144],
F_[9][1][144],
F_[9][2][144],
F_[10][0][144],
F_[10][1][144],
F_[10][2][144],
F_[11][0][144],
F_[11][1][144],
F_[11][2][144],
F_[12][0][144],
F_[12][1][144],
F_[12][2][144],
F_[13][0][144],
F_[13][1][144],
F_[13][2][144],
F_[14][0][144],
F_[14][1][144],
F_[14][2][144],
F_[15][0][144],
F_[15][1][144],
F_[15][2][144],
F_[0][0][145],
F_[0][1][145],
F_[0][2][145],
F_[1][0][145],
F_[1][1][145],
F_[1][2][145],
F_[2][0][145],
F_[2][1][145],
F_[2][2][145],
F_[3][0][145],
F_[3][1][145],
F_[3][2][145],
F_[4][0][145],
F_[4][1][145],
F_[4][2][145],
F_[5][0][145],
F_[5][1][145],
F_[5][2][145],
F_[6][0][145],
F_[6][1][145],
F_[6][2][145],
F_[7][0][145],
F_[7][1][145],
F_[7][2][145],
F_[8][0][145],
F_[8][1][145],
F_[8][2][145],
F_[9][0][145],
F_[9][1][145],
F_[9][2][145],
F_[10][0][145],
F_[10][1][145],
F_[10][2][145],
F_[11][0][145],
F_[11][1][145],
F_[11][2][145],
F_[12][0][145],
F_[12][1][145],
F_[12][2][145],
F_[13][0][145],
F_[13][1][145],
F_[13][2][145],
F_[14][0][145],
F_[14][1][145],
F_[14][2][145],
F_[15][0][145],
F_[15][1][145],
F_[15][2][145],
F_[0][0][146],
F_[0][1][146],
F_[0][2][146],
F_[1][0][146],
F_[1][1][146],
F_[1][2][146],
F_[2][0][146],
F_[2][1][146],
F_[2][2][146],
F_[3][0][146],
F_[3][1][146],
F_[3][2][146],
F_[4][0][146],
F_[4][1][146],
F_[4][2][146],
F_[5][0][146],
F_[5][1][146],
F_[5][2][146],
F_[6][0][146],
F_[6][1][146],
F_[6][2][146],
F_[7][0][146],
F_[7][1][146],
F_[7][2][146],
F_[8][0][146],
F_[8][1][146],
F_[8][2][146],
F_[9][0][146],
F_[9][1][146],
F_[9][2][146],
F_[10][0][146],
F_[10][1][146],
F_[10][2][146],
F_[11][0][146],
F_[11][1][146],
F_[11][2][146],
F_[12][0][146],
F_[12][1][146],
F_[12][2][146],
F_[13][0][146],
F_[13][1][146],
F_[13][2][146],
F_[14][0][146],
F_[14][1][146],
F_[14][2][146],
F_[15][0][146],
F_[15][1][146],
F_[15][2][146],
F_[0][0][147],
F_[0][1][147],
F_[0][2][147],
F_[1][0][147],
F_[1][1][147],
F_[1][2][147],
F_[2][0][147],
F_[2][1][147],
F_[2][2][147],
F_[3][0][147],
F_[3][1][147],
F_[3][2][147],
F_[4][0][147],
F_[4][1][147],
F_[4][2][147],
F_[5][0][147],
F_[5][1][147],
F_[5][2][147],
F_[6][0][147],
F_[6][1][147],
F_[6][2][147],
F_[7][0][147],
F_[7][1][147],
F_[7][2][147],
F_[8][0][147],
F_[8][1][147],
F_[8][2][147],
F_[9][0][147],
F_[9][1][147],
F_[9][2][147],
F_[10][0][147],
F_[10][1][147],
F_[10][2][147],
F_[11][0][147],
F_[11][1][147],
F_[11][2][147],
F_[12][0][147],
F_[12][1][147],
F_[12][2][147],
F_[13][0][147],
F_[13][1][147],
F_[13][2][147],
F_[14][0][147],
F_[14][1][147],
F_[14][2][147],
F_[15][0][147],
F_[15][1][147],
F_[15][2][147],
F_[0][0][148],
F_[0][1][148],
F_[0][2][148],
F_[1][0][148],
F_[1][1][148],
F_[1][2][148],
F_[2][0][148],
F_[2][1][148],
F_[2][2][148],
F_[3][0][148],
F_[3][1][148],
F_[3][2][148],
F_[4][0][148],
F_[4][1][148],
F_[4][2][148],
F_[5][0][148],
F_[5][1][148],
F_[5][2][148],
F_[6][0][148],
F_[6][1][148],
F_[6][2][148],
F_[7][0][148],
F_[7][1][148],
F_[7][2][148],
F_[8][0][148],
F_[8][1][148],
F_[8][2][148],
F_[9][0][148],
F_[9][1][148],
F_[9][2][148],
F_[10][0][148],
F_[10][1][148],
F_[10][2][148],
F_[11][0][148],
F_[11][1][148],
F_[11][2][148],
F_[12][0][148],
F_[12][1][148],
F_[12][2][148],
F_[13][0][148],
F_[13][1][148],
F_[13][2][148],
F_[14][0][148],
F_[14][1][148],
F_[14][2][148],
F_[15][0][148],
F_[15][1][148],
F_[15][2][148],
F_[0][0][149],
F_[0][1][149],
F_[0][2][149],
F_[1][0][149],
F_[1][1][149],
F_[1][2][149],
F_[2][0][149],
F_[2][1][149],
F_[2][2][149],
F_[3][0][149],
F_[3][1][149],
F_[3][2][149],
F_[4][0][149],
F_[4][1][149],
F_[4][2][149],
F_[5][0][149],
F_[5][1][149],
F_[5][2][149],
F_[6][0][149],
F_[6][1][149],
F_[6][2][149],
F_[7][0][149],
F_[7][1][149],
F_[7][2][149],
F_[8][0][149],
F_[8][1][149],
F_[8][2][149],
F_[9][0][149],
F_[9][1][149],
F_[9][2][149],
F_[10][0][149],
F_[10][1][149],
F_[10][2][149],
F_[11][0][149],
F_[11][1][149],
F_[11][2][149],
F_[12][0][149],
F_[12][1][149],
F_[12][2][149],
F_[13][0][149],
F_[13][1][149],
F_[13][2][149],
F_[14][0][149],
F_[14][1][149],
F_[14][2][149],
F_[15][0][149],
F_[15][1][149],
F_[15][2][149],
F_[0][0][150],
F_[0][1][150],
F_[0][2][150],
F_[1][0][150],
F_[1][1][150],
F_[1][2][150],
F_[2][0][150],
F_[2][1][150],
F_[2][2][150],
F_[3][0][150],
F_[3][1][150],
F_[3][2][150],
F_[4][0][150],
F_[4][1][150],
F_[4][2][150],
F_[5][0][150],
F_[5][1][150],
F_[5][2][150],
F_[6][0][150],
F_[6][1][150],
F_[6][2][150],
F_[7][0][150],
F_[7][1][150],
F_[7][2][150],
F_[8][0][150],
F_[8][1][150],
F_[8][2][150],
F_[9][0][150],
F_[9][1][150],
F_[9][2][150],
F_[10][0][150],
F_[10][1][150],
F_[10][2][150],
F_[11][0][150],
F_[11][1][150],
F_[11][2][150],
F_[12][0][150],
F_[12][1][150],
F_[12][2][150],
F_[13][0][150],
F_[13][1][150],
F_[13][2][150],
F_[14][0][150],
F_[14][1][150],
F_[14][2][150],
F_[15][0][150],
F_[15][1][150],
F_[15][2][150],
F_[0][0][151],
F_[0][1][151],
F_[0][2][151],
F_[1][0][151],
F_[1][1][151],
F_[1][2][151],
F_[2][0][151],
F_[2][1][151],
F_[2][2][151],
F_[3][0][151],
F_[3][1][151],
F_[3][2][151],
F_[4][0][151],
F_[4][1][151],
F_[4][2][151],
F_[5][0][151],
F_[5][1][151],
F_[5][2][151],
F_[6][0][151],
F_[6][1][151],
F_[6][2][151],
F_[7][0][151],
F_[7][1][151],
F_[7][2][151],
F_[8][0][151],
F_[8][1][151],
F_[8][2][151],
F_[9][0][151],
F_[9][1][151],
F_[9][2][151],
F_[10][0][151],
F_[10][1][151],
F_[10][2][151],
F_[11][0][151],
F_[11][1][151],
F_[11][2][151],
F_[12][0][151],
F_[12][1][151],
F_[12][2][151],
F_[13][0][151],
F_[13][1][151],
F_[13][2][151],
F_[14][0][151],
F_[14][1][151],
F_[14][2][151],
F_[15][0][151],
F_[15][1][151],
F_[15][2][151],
F_[0][0][152],
F_[0][1][152],
F_[0][2][152],
F_[1][0][152],
F_[1][1][152],
F_[1][2][152],
F_[2][0][152],
F_[2][1][152],
F_[2][2][152],
F_[3][0][152],
F_[3][1][152],
F_[3][2][152],
F_[4][0][152],
F_[4][1][152],
F_[4][2][152],
F_[5][0][152],
F_[5][1][152],
F_[5][2][152],
F_[6][0][152],
F_[6][1][152],
F_[6][2][152],
F_[7][0][152],
F_[7][1][152],
F_[7][2][152],
F_[8][0][152],
F_[8][1][152],
F_[8][2][152],
F_[9][0][152],
F_[9][1][152],
F_[9][2][152],
F_[10][0][152],
F_[10][1][152],
F_[10][2][152],
F_[11][0][152],
F_[11][1][152],
F_[11][2][152],
F_[12][0][152],
F_[12][1][152],
F_[12][2][152],
F_[13][0][152],
F_[13][1][152],
F_[13][2][152],
F_[14][0][152],
F_[14][1][152],
F_[14][2][152],
F_[15][0][152],
F_[15][1][152],
F_[15][2][152],
F_[0][0][153],
F_[0][1][153],
F_[0][2][153],
F_[1][0][153],
F_[1][1][153],
F_[1][2][153],
F_[2][0][153],
F_[2][1][153],
F_[2][2][153],
F_[3][0][153],
F_[3][1][153],
F_[3][2][153],
F_[4][0][153],
F_[4][1][153],
F_[4][2][153],
F_[5][0][153],
F_[5][1][153],
F_[5][2][153],
F_[6][0][153],
F_[6][1][153],
F_[6][2][153],
F_[7][0][153],
F_[7][1][153],
F_[7][2][153],
F_[8][0][153],
F_[8][1][153],
F_[8][2][153],
F_[9][0][153],
F_[9][1][153],
F_[9][2][153],
F_[10][0][153],
F_[10][1][153],
F_[10][2][153],
F_[11][0][153],
F_[11][1][153],
F_[11][2][153],
F_[12][0][153],
F_[12][1][153],
F_[12][2][153],
F_[13][0][153],
F_[13][1][153],
F_[13][2][153],
F_[14][0][153],
F_[14][1][153],
F_[14][2][153],
F_[15][0][153],
F_[15][1][153],
F_[15][2][153],
F_[0][0][154],
F_[0][1][154],
F_[0][2][154],
F_[1][0][154],
F_[1][1][154],
F_[1][2][154],
F_[2][0][154],
F_[2][1][154],
F_[2][2][154],
F_[3][0][154],
F_[3][1][154],
F_[3][2][154],
F_[4][0][154],
F_[4][1][154],
F_[4][2][154],
F_[5][0][154],
F_[5][1][154],
F_[5][2][154],
F_[6][0][154],
F_[6][1][154],
F_[6][2][154],
F_[7][0][154],
F_[7][1][154],
F_[7][2][154],
F_[8][0][154],
F_[8][1][154],
F_[8][2][154],
F_[9][0][154],
F_[9][1][154],
F_[9][2][154],
F_[10][0][154],
F_[10][1][154],
F_[10][2][154],
F_[11][0][154],
F_[11][1][154],
F_[11][2][154],
F_[12][0][154],
F_[12][1][154],
F_[12][2][154],
F_[13][0][154],
F_[13][1][154],
F_[13][2][154],
F_[14][0][154],
F_[14][1][154],
F_[14][2][154],
F_[15][0][154],
F_[15][1][154],
F_[15][2][154],
F_[0][0][155],
F_[0][1][155],
F_[0][2][155],
F_[1][0][155],
F_[1][1][155],
F_[1][2][155],
F_[2][0][155],
F_[2][1][155],
F_[2][2][155],
F_[3][0][155],
F_[3][1][155],
F_[3][2][155],
F_[4][0][155],
F_[4][1][155],
F_[4][2][155],
F_[5][0][155],
F_[5][1][155],
F_[5][2][155],
F_[6][0][155],
F_[6][1][155],
F_[6][2][155],
F_[7][0][155],
F_[7][1][155],
F_[7][2][155],
F_[8][0][155],
F_[8][1][155],
F_[8][2][155],
F_[9][0][155],
F_[9][1][155],
F_[9][2][155],
F_[10][0][155],
F_[10][1][155],
F_[10][2][155],
F_[11][0][155],
F_[11][1][155],
F_[11][2][155],
F_[12][0][155],
F_[12][1][155],
F_[12][2][155],
F_[13][0][155],
F_[13][1][155],
F_[13][2][155],
F_[14][0][155],
F_[14][1][155],
F_[14][2][155],
F_[15][0][155],
F_[15][1][155],
F_[15][2][155],
F_[0][0][156],
F_[0][1][156],
F_[0][2][156],
F_[1][0][156],
F_[1][1][156],
F_[1][2][156],
F_[2][0][156],
F_[2][1][156],
F_[2][2][156],
F_[3][0][156],
F_[3][1][156],
F_[3][2][156],
F_[4][0][156],
F_[4][1][156],
F_[4][2][156],
F_[5][0][156],
F_[5][1][156],
F_[5][2][156],
F_[6][0][156],
F_[6][1][156],
F_[6][2][156],
F_[7][0][156],
F_[7][1][156],
F_[7][2][156],
F_[8][0][156],
F_[8][1][156],
F_[8][2][156],
F_[9][0][156],
F_[9][1][156],
F_[9][2][156],
F_[10][0][156],
F_[10][1][156],
F_[10][2][156],
F_[11][0][156],
F_[11][1][156],
F_[11][2][156],
F_[12][0][156],
F_[12][1][156],
F_[12][2][156],
F_[13][0][156],
F_[13][1][156],
F_[13][2][156],
F_[14][0][156],
F_[14][1][156],
F_[14][2][156],
F_[15][0][156],
F_[15][1][156],
F_[15][2][156],
F_[0][0][157],
F_[0][1][157],
F_[0][2][157],
F_[1][0][157],
F_[1][1][157],
F_[1][2][157],
F_[2][0][157],
F_[2][1][157],
F_[2][2][157],
F_[3][0][157],
F_[3][1][157],
F_[3][2][157],
F_[4][0][157],
F_[4][1][157],
F_[4][2][157],
F_[5][0][157],
F_[5][1][157],
F_[5][2][157],
F_[6][0][157],
F_[6][1][157],
F_[6][2][157],
F_[7][0][157],
F_[7][1][157],
F_[7][2][157],
F_[8][0][157],
F_[8][1][157],
F_[8][2][157],
F_[9][0][157],
F_[9][1][157],
F_[9][2][157],
F_[10][0][157],
F_[10][1][157],
F_[10][2][157],
F_[11][0][157],
F_[11][1][157],
F_[11][2][157],
F_[12][0][157],
F_[12][1][157],
F_[12][2][157],
F_[13][0][157],
F_[13][1][157],
F_[13][2][157],
F_[14][0][157],
F_[14][1][157],
F_[14][2][157],
F_[15][0][157],
F_[15][1][157],
F_[15][2][157],
F_[0][0][158],
F_[0][1][158],
F_[0][2][158],
F_[1][0][158],
F_[1][1][158],
F_[1][2][158],
F_[2][0][158],
F_[2][1][158],
F_[2][2][158],
F_[3][0][158],
F_[3][1][158],
F_[3][2][158],
F_[4][0][158],
F_[4][1][158],
F_[4][2][158],
F_[5][0][158],
F_[5][1][158],
F_[5][2][158],
F_[6][0][158],
F_[6][1][158],
F_[6][2][158],
F_[7][0][158],
F_[7][1][158],
F_[7][2][158],
F_[8][0][158],
F_[8][1][158],
F_[8][2][158],
F_[9][0][158],
F_[9][1][158],
F_[9][2][158],
F_[10][0][158],
F_[10][1][158],
F_[10][2][158],
F_[11][0][158],
F_[11][1][158],
F_[11][2][158],
F_[12][0][158],
F_[12][1][158],
F_[12][2][158],
F_[13][0][158],
F_[13][1][158],
F_[13][2][158],
F_[14][0][158],
F_[14][1][158],
F_[14][2][158],
F_[15][0][158],
F_[15][1][158],
F_[15][2][158],
F_[0][0][159],
F_[0][1][159],
F_[0][2][159],
F_[1][0][159],
F_[1][1][159],
F_[1][2][159],
F_[2][0][159],
F_[2][1][159],
F_[2][2][159],
F_[3][0][159],
F_[3][1][159],
F_[3][2][159],
F_[4][0][159],
F_[4][1][159],
F_[4][2][159],
F_[5][0][159],
F_[5][1][159],
F_[5][2][159],
F_[6][0][159],
F_[6][1][159],
F_[6][2][159],
F_[7][0][159],
F_[7][1][159],
F_[7][2][159],
F_[8][0][159],
F_[8][1][159],
F_[8][2][159],
F_[9][0][159],
F_[9][1][159],
F_[9][2][159],
F_[10][0][159],
F_[10][1][159],
F_[10][2][159],
F_[11][0][159],
F_[11][1][159],
F_[11][2][159],
F_[12][0][159],
F_[12][1][159],
F_[12][2][159],
F_[13][0][159],
F_[13][1][159],
F_[13][2][159],
F_[14][0][159],
F_[14][1][159],
F_[14][2][159],
F_[15][0][159],
F_[15][1][159],
F_[15][2][159],
F_[0][0][160],
F_[0][1][160],
F_[0][2][160],
F_[1][0][160],
F_[1][1][160],
F_[1][2][160],
F_[2][0][160],
F_[2][1][160],
F_[2][2][160],
F_[3][0][160],
F_[3][1][160],
F_[3][2][160],
F_[4][0][160],
F_[4][1][160],
F_[4][2][160],
F_[5][0][160],
F_[5][1][160],
F_[5][2][160],
F_[6][0][160],
F_[6][1][160],
F_[6][2][160],
F_[7][0][160],
F_[7][1][160],
F_[7][2][160],
F_[8][0][160],
F_[8][1][160],
F_[8][2][160],
F_[9][0][160],
F_[9][1][160],
F_[9][2][160],
F_[10][0][160],
F_[10][1][160],
F_[10][2][160],
F_[11][0][160],
F_[11][1][160],
F_[11][2][160],
F_[12][0][160],
F_[12][1][160],
F_[12][2][160],
F_[13][0][160],
F_[13][1][160],
F_[13][2][160],
F_[14][0][160],
F_[14][1][160],
F_[14][2][160],
F_[15][0][160],
F_[15][1][160],
F_[15][2][160],
F_[0][0][161],
F_[0][1][161],
F_[0][2][161],
F_[1][0][161],
F_[1][1][161],
F_[1][2][161],
F_[2][0][161],
F_[2][1][161],
F_[2][2][161],
F_[3][0][161],
F_[3][1][161],
F_[3][2][161],
F_[4][0][161],
F_[4][1][161],
F_[4][2][161],
F_[5][0][161],
F_[5][1][161],
F_[5][2][161],
F_[6][0][161],
F_[6][1][161],
F_[6][2][161],
F_[7][0][161],
F_[7][1][161],
F_[7][2][161],
F_[8][0][161],
F_[8][1][161],
F_[8][2][161],
F_[9][0][161],
F_[9][1][161],
F_[9][2][161],
F_[10][0][161],
F_[10][1][161],
F_[10][2][161],
F_[11][0][161],
F_[11][1][161],
F_[11][2][161],
F_[12][0][161],
F_[12][1][161],
F_[12][2][161],
F_[13][0][161],
F_[13][1][161],
F_[13][2][161],
F_[14][0][161],
F_[14][1][161],
F_[14][2][161],
F_[15][0][161],
F_[15][1][161],
F_[15][2][161],
F_[0][0][162],
F_[0][1][162],
F_[0][2][162],
F_[1][0][162],
F_[1][1][162],
F_[1][2][162],
F_[2][0][162],
F_[2][1][162],
F_[2][2][162],
F_[3][0][162],
F_[3][1][162],
F_[3][2][162],
F_[4][0][162],
F_[4][1][162],
F_[4][2][162],
F_[5][0][162],
F_[5][1][162],
F_[5][2][162],
F_[6][0][162],
F_[6][1][162],
F_[6][2][162],
F_[7][0][162],
F_[7][1][162],
F_[7][2][162],
F_[8][0][162],
F_[8][1][162],
F_[8][2][162],
F_[9][0][162],
F_[9][1][162],
F_[9][2][162],
F_[10][0][162],
F_[10][1][162],
F_[10][2][162],
F_[11][0][162],
F_[11][1][162],
F_[11][2][162],
F_[12][0][162],
F_[12][1][162],
F_[12][2][162],
F_[13][0][162],
F_[13][1][162],
F_[13][2][162],
F_[14][0][162],
F_[14][1][162],
F_[14][2][162],
F_[15][0][162],
F_[15][1][162],
F_[15][2][162],
F_[0][0][163],
F_[0][1][163],
F_[0][2][163],
F_[1][0][163],
F_[1][1][163],
F_[1][2][163],
F_[2][0][163],
F_[2][1][163],
F_[2][2][163],
F_[3][0][163],
F_[3][1][163],
F_[3][2][163],
F_[4][0][163],
F_[4][1][163],
F_[4][2][163],
F_[5][0][163],
F_[5][1][163],
F_[5][2][163],
F_[6][0][163],
F_[6][1][163],
F_[6][2][163],
F_[7][0][163],
F_[7][1][163],
F_[7][2][163],
F_[8][0][163],
F_[8][1][163],
F_[8][2][163],
F_[9][0][163],
F_[9][1][163],
F_[9][2][163],
F_[10][0][163],
F_[10][1][163],
F_[10][2][163],
F_[11][0][163],
F_[11][1][163],
F_[11][2][163],
F_[12][0][163],
F_[12][1][163],
F_[12][2][163],
F_[13][0][163],
F_[13][1][163],
F_[13][2][163],
F_[14][0][163],
F_[14][1][163],
F_[14][2][163],
F_[15][0][163],
F_[15][1][163],
F_[15][2][163],
F_[0][0][164],
F_[0][1][164],
F_[0][2][164],
F_[1][0][164],
F_[1][1][164],
F_[1][2][164],
F_[2][0][164],
F_[2][1][164],
F_[2][2][164],
F_[3][0][164],
F_[3][1][164],
F_[3][2][164],
F_[4][0][164],
F_[4][1][164],
F_[4][2][164],
F_[5][0][164],
F_[5][1][164],
F_[5][2][164],
F_[6][0][164],
F_[6][1][164],
F_[6][2][164],
F_[7][0][164],
F_[7][1][164],
F_[7][2][164],
F_[8][0][164],
F_[8][1][164],
F_[8][2][164],
F_[9][0][164],
F_[9][1][164],
F_[9][2][164],
F_[10][0][164],
F_[10][1][164],
F_[10][2][164],
F_[11][0][164],
F_[11][1][164],
F_[11][2][164],
F_[12][0][164],
F_[12][1][164],
F_[12][2][164],
F_[13][0][164],
F_[13][1][164],
F_[13][2][164],
F_[14][0][164],
F_[14][1][164],
F_[14][2][164],
F_[15][0][164],
F_[15][1][164],
F_[15][2][164],
F_[0][0][165],
F_[0][1][165],
F_[0][2][165],
F_[1][0][165],
F_[1][1][165],
F_[1][2][165],
F_[2][0][165],
F_[2][1][165],
F_[2][2][165],
F_[3][0][165],
F_[3][1][165],
F_[3][2][165],
F_[4][0][165],
F_[4][1][165],
F_[4][2][165],
F_[5][0][165],
F_[5][1][165],
F_[5][2][165],
F_[6][0][165],
F_[6][1][165],
F_[6][2][165],
F_[7][0][165],
F_[7][1][165],
F_[7][2][165],
F_[8][0][165],
F_[8][1][165],
F_[8][2][165],
F_[9][0][165],
F_[9][1][165],
F_[9][2][165],
F_[10][0][165],
F_[10][1][165],
F_[10][2][165],
F_[11][0][165],
F_[11][1][165],
F_[11][2][165],
F_[12][0][165],
F_[12][1][165],
F_[12][2][165],
F_[13][0][165],
F_[13][1][165],
F_[13][2][165],
F_[14][0][165],
F_[14][1][165],
F_[14][2][165],
F_[15][0][165],
F_[15][1][165],
F_[15][2][165],
F_[0][0][166],
F_[0][1][166],
F_[0][2][166],
F_[1][0][166],
F_[1][1][166],
F_[1][2][166],
F_[2][0][166],
F_[2][1][166],
F_[2][2][166],
F_[3][0][166],
F_[3][1][166],
F_[3][2][166],
F_[4][0][166],
F_[4][1][166],
F_[4][2][166],
F_[5][0][166],
F_[5][1][166],
F_[5][2][166],
F_[6][0][166],
F_[6][1][166],
F_[6][2][166],
F_[7][0][166],
F_[7][1][166],
F_[7][2][166],
F_[8][0][166],
F_[8][1][166],
F_[8][2][166],
F_[9][0][166],
F_[9][1][166],
F_[9][2][166],
F_[10][0][166],
F_[10][1][166],
F_[10][2][166],
F_[11][0][166],
F_[11][1][166],
F_[11][2][166],
F_[12][0][166],
F_[12][1][166],
F_[12][2][166],
F_[13][0][166],
F_[13][1][166],
F_[13][2][166],
F_[14][0][166],
F_[14][1][166],
F_[14][2][166],
F_[15][0][166],
F_[15][1][166],
F_[15][2][166],
F_[0][0][167],
F_[0][1][167],
F_[0][2][167],
F_[1][0][167],
F_[1][1][167],
F_[1][2][167],
F_[2][0][167],
F_[2][1][167],
F_[2][2][167],
F_[3][0][167],
F_[3][1][167],
F_[3][2][167],
F_[4][0][167],
F_[4][1][167],
F_[4][2][167],
F_[5][0][167],
F_[5][1][167],
F_[5][2][167],
F_[6][0][167],
F_[6][1][167],
F_[6][2][167],
F_[7][0][167],
F_[7][1][167],
F_[7][2][167],
F_[8][0][167],
F_[8][1][167],
F_[8][2][167],
F_[9][0][167],
F_[9][1][167],
F_[9][2][167],
F_[10][0][167],
F_[10][1][167],
F_[10][2][167],
F_[11][0][167],
F_[11][1][167],
F_[11][2][167],
F_[12][0][167],
F_[12][1][167],
F_[12][2][167],
F_[13][0][167],
F_[13][1][167],
F_[13][2][167],
F_[14][0][167],
F_[14][1][167],
F_[14][2][167],
F_[15][0][167],
F_[15][1][167],
F_[15][2][167],
F_[0][0][168],
F_[0][1][168],
F_[0][2][168],
F_[1][0][168],
F_[1][1][168],
F_[1][2][168],
F_[2][0][168],
F_[2][1][168],
F_[2][2][168],
F_[3][0][168],
F_[3][1][168],
F_[3][2][168],
F_[4][0][168],
F_[4][1][168],
F_[4][2][168],
F_[5][0][168],
F_[5][1][168],
F_[5][2][168],
F_[6][0][168],
F_[6][1][168],
F_[6][2][168],
F_[7][0][168],
F_[7][1][168],
F_[7][2][168],
F_[8][0][168],
F_[8][1][168],
F_[8][2][168],
F_[9][0][168],
F_[9][1][168],
F_[9][2][168],
F_[10][0][168],
F_[10][1][168],
F_[10][2][168],
F_[11][0][168],
F_[11][1][168],
F_[11][2][168],
F_[12][0][168],
F_[12][1][168],
F_[12][2][168],
F_[13][0][168],
F_[13][1][168],
F_[13][2][168],
F_[14][0][168],
F_[14][1][168],
F_[14][2][168],
F_[15][0][168],
F_[15][1][168],
F_[15][2][168],
F_[0][0][169],
F_[0][1][169],
F_[0][2][169],
F_[1][0][169],
F_[1][1][169],
F_[1][2][169],
F_[2][0][169],
F_[2][1][169],
F_[2][2][169],
F_[3][0][169],
F_[3][1][169],
F_[3][2][169],
F_[4][0][169],
F_[4][1][169],
F_[4][2][169],
F_[5][0][169],
F_[5][1][169],
F_[5][2][169],
F_[6][0][169],
F_[6][1][169],
F_[6][2][169],
F_[7][0][169],
F_[7][1][169],
F_[7][2][169],
F_[8][0][169],
F_[8][1][169],
F_[8][2][169],
F_[9][0][169],
F_[9][1][169],
F_[9][2][169],
F_[10][0][169],
F_[10][1][169],
F_[10][2][169],
F_[11][0][169],
F_[11][1][169],
F_[11][2][169],
F_[12][0][169],
F_[12][1][169],
F_[12][2][169],
F_[13][0][169],
F_[13][1][169],
F_[13][2][169],
F_[14][0][169],
F_[14][1][169],
F_[14][2][169],
F_[15][0][169],
F_[15][1][169],
F_[15][2][169],
F_[0][0][170],
F_[0][1][170],
F_[0][2][170],
F_[1][0][170],
F_[1][1][170],
F_[1][2][170],
F_[2][0][170],
F_[2][1][170],
F_[2][2][170],
F_[3][0][170],
F_[3][1][170],
F_[3][2][170],
F_[4][0][170],
F_[4][1][170],
F_[4][2][170],
F_[5][0][170],
F_[5][1][170],
F_[5][2][170],
F_[6][0][170],
F_[6][1][170],
F_[6][2][170],
F_[7][0][170],
F_[7][1][170],
F_[7][2][170],
F_[8][0][170],
F_[8][1][170],
F_[8][2][170],
F_[9][0][170],
F_[9][1][170],
F_[9][2][170],
F_[10][0][170],
F_[10][1][170],
F_[10][2][170],
F_[11][0][170],
F_[11][1][170],
F_[11][2][170],
F_[12][0][170],
F_[12][1][170],
F_[12][2][170],
F_[13][0][170],
F_[13][1][170],
F_[13][2][170],
F_[14][0][170],
F_[14][1][170],
F_[14][2][170],
F_[15][0][170],
F_[15][1][170],
F_[15][2][170],
F_[0][0][171],
F_[0][1][171],
F_[0][2][171],
F_[1][0][171],
F_[1][1][171],
F_[1][2][171],
F_[2][0][171],
F_[2][1][171],
F_[2][2][171],
F_[3][0][171],
F_[3][1][171],
F_[3][2][171],
F_[4][0][171],
F_[4][1][171],
F_[4][2][171],
F_[5][0][171],
F_[5][1][171],
F_[5][2][171],
F_[6][0][171],
F_[6][1][171],
F_[6][2][171],
F_[7][0][171],
F_[7][1][171],
F_[7][2][171],
F_[8][0][171],
F_[8][1][171],
F_[8][2][171],
F_[9][0][171],
F_[9][1][171],
F_[9][2][171],
F_[10][0][171],
F_[10][1][171],
F_[10][2][171],
F_[11][0][171],
F_[11][1][171],
F_[11][2][171],
F_[12][0][171],
F_[12][1][171],
F_[12][2][171],
F_[13][0][171],
F_[13][1][171],
F_[13][2][171],
F_[14][0][171],
F_[14][1][171],
F_[14][2][171],
F_[15][0][171],
F_[15][1][171],
F_[15][2][171],
F_[0][0][172],
F_[0][1][172],
F_[0][2][172],
F_[1][0][172],
F_[1][1][172],
F_[1][2][172],
F_[2][0][172],
F_[2][1][172],
F_[2][2][172],
F_[3][0][172],
F_[3][1][172],
F_[3][2][172],
F_[4][0][172],
F_[4][1][172],
F_[4][2][172],
F_[5][0][172],
F_[5][1][172],
F_[5][2][172],
F_[6][0][172],
F_[6][1][172],
F_[6][2][172],
F_[7][0][172],
F_[7][1][172],
F_[7][2][172],
F_[8][0][172],
F_[8][1][172],
F_[8][2][172],
F_[9][0][172],
F_[9][1][172],
F_[9][2][172],
F_[10][0][172],
F_[10][1][172],
F_[10][2][172],
F_[11][0][172],
F_[11][1][172],
F_[11][2][172],
F_[12][0][172],
F_[12][1][172],
F_[12][2][172],
F_[13][0][172],
F_[13][1][172],
F_[13][2][172],
F_[14][0][172],
F_[14][1][172],
F_[14][2][172],
F_[15][0][172],
F_[15][1][172],
F_[15][2][172],
F_[0][0][173],
F_[0][1][173],
F_[0][2][173],
F_[1][0][173],
F_[1][1][173],
F_[1][2][173],
F_[2][0][173],
F_[2][1][173],
F_[2][2][173],
F_[3][0][173],
F_[3][1][173],
F_[3][2][173],
F_[4][0][173],
F_[4][1][173],
F_[4][2][173],
F_[5][0][173],
F_[5][1][173],
F_[5][2][173],
F_[6][0][173],
F_[6][1][173],
F_[6][2][173],
F_[7][0][173],
F_[7][1][173],
F_[7][2][173],
F_[8][0][173],
F_[8][1][173],
F_[8][2][173],
F_[9][0][173],
F_[9][1][173],
F_[9][2][173],
F_[10][0][173],
F_[10][1][173],
F_[10][2][173],
F_[11][0][173],
F_[11][1][173],
F_[11][2][173],
F_[12][0][173],
F_[12][1][173],
F_[12][2][173],
F_[13][0][173],
F_[13][1][173],
F_[13][2][173],
F_[14][0][173],
F_[14][1][173],
F_[14][2][173],
F_[15][0][173],
F_[15][1][173],
F_[15][2][173],
F_[0][0][174],
F_[0][1][174],
F_[0][2][174],
F_[1][0][174],
F_[1][1][174],
F_[1][2][174],
F_[2][0][174],
F_[2][1][174],
F_[2][2][174],
F_[3][0][174],
F_[3][1][174],
F_[3][2][174],
F_[4][0][174],
F_[4][1][174],
F_[4][2][174],
F_[5][0][174],
F_[5][1][174],
F_[5][2][174],
F_[6][0][174],
F_[6][1][174],
F_[6][2][174],
F_[7][0][174],
F_[7][1][174],
F_[7][2][174],
F_[8][0][174],
F_[8][1][174],
F_[8][2][174],
F_[9][0][174],
F_[9][1][174],
F_[9][2][174],
F_[10][0][174],
F_[10][1][174],
F_[10][2][174],
F_[11][0][174],
F_[11][1][174],
F_[11][2][174],
F_[12][0][174],
F_[12][1][174],
F_[12][2][174],
F_[13][0][174],
F_[13][1][174],
F_[13][2][174],
F_[14][0][174],
F_[14][1][174],
F_[14][2][174],
F_[15][0][174],
F_[15][1][174],
F_[15][2][174],
F_[0][0][175],
F_[0][1][175],
F_[0][2][175],
F_[1][0][175],
F_[1][1][175],
F_[1][2][175],
F_[2][0][175],
F_[2][1][175],
F_[2][2][175],
F_[3][0][175],
F_[3][1][175],
F_[3][2][175],
F_[4][0][175],
F_[4][1][175],
F_[4][2][175],
F_[5][0][175],
F_[5][1][175],
F_[5][2][175],
F_[6][0][175],
F_[6][1][175],
F_[6][2][175],
F_[7][0][175],
F_[7][1][175],
F_[7][2][175],
F_[8][0][175],
F_[8][1][175],
F_[8][2][175],
F_[9][0][175],
F_[9][1][175],
F_[9][2][175],
F_[10][0][175],
F_[10][1][175],
F_[10][2][175],
F_[11][0][175],
F_[11][1][175],
F_[11][2][175],
F_[12][0][175],
F_[12][1][175],
F_[12][2][175],
F_[13][0][175],
F_[13][1][175],
F_[13][2][175],
F_[14][0][175],
F_[14][1][175],
F_[14][2][175],
F_[15][0][175],
F_[15][1][175],
F_[15][2][175],
F_[0][0][176],
F_[0][1][176],
F_[0][2][176],
F_[1][0][176],
F_[1][1][176],
F_[1][2][176],
F_[2][0][176],
F_[2][1][176],
F_[2][2][176],
F_[3][0][176],
F_[3][1][176],
F_[3][2][176],
F_[4][0][176],
F_[4][1][176],
F_[4][2][176],
F_[5][0][176],
F_[5][1][176],
F_[5][2][176],
F_[6][0][176],
F_[6][1][176],
F_[6][2][176],
F_[7][0][176],
F_[7][1][176],
F_[7][2][176],
F_[8][0][176],
F_[8][1][176],
F_[8][2][176],
F_[9][0][176],
F_[9][1][176],
F_[9][2][176],
F_[10][0][176],
F_[10][1][176],
F_[10][2][176],
F_[11][0][176],
F_[11][1][176],
F_[11][2][176],
F_[12][0][176],
F_[12][1][176],
F_[12][2][176],
F_[13][0][176],
F_[13][1][176],
F_[13][2][176],
F_[14][0][176],
F_[14][1][176],
F_[14][2][176],
F_[15][0][176],
F_[15][1][176],
F_[15][2][176],
F_[0][0][177],
F_[0][1][177],
F_[0][2][177],
F_[1][0][177],
F_[1][1][177],
F_[1][2][177],
F_[2][0][177],
F_[2][1][177],
F_[2][2][177],
F_[3][0][177],
F_[3][1][177],
F_[3][2][177],
F_[4][0][177],
F_[4][1][177],
F_[4][2][177],
F_[5][0][177],
F_[5][1][177],
F_[5][2][177],
F_[6][0][177],
F_[6][1][177],
F_[6][2][177],
F_[7][0][177],
F_[7][1][177],
F_[7][2][177],
F_[8][0][177],
F_[8][1][177],
F_[8][2][177],
F_[9][0][177],
F_[9][1][177],
F_[9][2][177],
F_[10][0][177],
F_[10][1][177],
F_[10][2][177],
F_[11][0][177],
F_[11][1][177],
F_[11][2][177],
F_[12][0][177],
F_[12][1][177],
F_[12][2][177],
F_[13][0][177],
F_[13][1][177],
F_[13][2][177],
F_[14][0][177],
F_[14][1][177],
F_[14][2][177],
F_[15][0][177],
F_[15][1][177],
F_[15][2][177],
F_[0][0][178],
F_[0][1][178],
F_[0][2][178],
F_[1][0][178],
F_[1][1][178],
F_[1][2][178],
F_[2][0][178],
F_[2][1][178],
F_[2][2][178],
F_[3][0][178],
F_[3][1][178],
F_[3][2][178],
F_[4][0][178],
F_[4][1][178],
F_[4][2][178],
F_[5][0][178],
F_[5][1][178],
F_[5][2][178],
F_[6][0][178],
F_[6][1][178],
F_[6][2][178],
F_[7][0][178],
F_[7][1][178],
F_[7][2][178],
F_[8][0][178],
F_[8][1][178],
F_[8][2][178],
F_[9][0][178],
F_[9][1][178],
F_[9][2][178],
F_[10][0][178],
F_[10][1][178],
F_[10][2][178],
F_[11][0][178],
F_[11][1][178],
F_[11][2][178],
F_[12][0][178],
F_[12][1][178],
F_[12][2][178],
F_[13][0][178],
F_[13][1][178],
F_[13][2][178],
F_[14][0][178],
F_[14][1][178],
F_[14][2][178],
F_[15][0][178],
F_[15][1][178],
F_[15][2][178],
F_[0][0][179],
F_[0][1][179],
F_[0][2][179],
F_[1][0][179],
F_[1][1][179],
F_[1][2][179],
F_[2][0][179],
F_[2][1][179],
F_[2][2][179],
F_[3][0][179],
F_[3][1][179],
F_[3][2][179],
F_[4][0][179],
F_[4][1][179],
F_[4][2][179],
F_[5][0][179],
F_[5][1][179],
F_[5][2][179],
F_[6][0][179],
F_[6][1][179],
F_[6][2][179],
F_[7][0][179],
F_[7][1][179],
F_[7][2][179],
F_[8][0][179],
F_[8][1][179],
F_[8][2][179],
F_[9][0][179],
F_[9][1][179],
F_[9][2][179],
F_[10][0][179],
F_[10][1][179],
F_[10][2][179],
F_[11][0][179],
F_[11][1][179],
F_[11][2][179],
F_[12][0][179],
F_[12][1][179],
F_[12][2][179],
F_[13][0][179],
F_[13][1][179],
F_[13][2][179],
F_[14][0][179],
F_[14][1][179],
F_[14][2][179],
F_[15][0][179],
F_[15][1][179],
F_[15][2][179],
F_[0][0][180],
F_[0][1][180],
F_[0][2][180],
F_[1][0][180],
F_[1][1][180],
F_[1][2][180],
F_[2][0][180],
F_[2][1][180],
F_[2][2][180],
F_[3][0][180],
F_[3][1][180],
F_[3][2][180],
F_[4][0][180],
F_[4][1][180],
F_[4][2][180],
F_[5][0][180],
F_[5][1][180],
F_[5][2][180],
F_[6][0][180],
F_[6][1][180],
F_[6][2][180],
F_[7][0][180],
F_[7][1][180],
F_[7][2][180],
F_[8][0][180],
F_[8][1][180],
F_[8][2][180],
F_[9][0][180],
F_[9][1][180],
F_[9][2][180],
F_[10][0][180],
F_[10][1][180],
F_[10][2][180],
F_[11][0][180],
F_[11][1][180],
F_[11][2][180],
F_[12][0][180],
F_[12][1][180],
F_[12][2][180],
F_[13][0][180],
F_[13][1][180],
F_[13][2][180],
F_[14][0][180],
F_[14][1][180],
F_[14][2][180],
F_[15][0][180],
F_[15][1][180],
F_[15][2][180],
F_[0][0][181],
F_[0][1][181],
F_[0][2][181],
F_[1][0][181],
F_[1][1][181],
F_[1][2][181],
F_[2][0][181],
F_[2][1][181],
F_[2][2][181],
F_[3][0][181],
F_[3][1][181],
F_[3][2][181],
F_[4][0][181],
F_[4][1][181],
F_[4][2][181],
F_[5][0][181],
F_[5][1][181],
F_[5][2][181],
F_[6][0][181],
F_[6][1][181],
F_[6][2][181],
F_[7][0][181],
F_[7][1][181],
F_[7][2][181],
F_[8][0][181],
F_[8][1][181],
F_[8][2][181],
F_[9][0][181],
F_[9][1][181],
F_[9][2][181],
F_[10][0][181],
F_[10][1][181],
F_[10][2][181],
F_[11][0][181],
F_[11][1][181],
F_[11][2][181],
F_[12][0][181],
F_[12][1][181],
F_[12][2][181],
F_[13][0][181],
F_[13][1][181],
F_[13][2][181],
F_[14][0][181],
F_[14][1][181],
F_[14][2][181],
F_[15][0][181],
F_[15][1][181],
F_[15][2][181],
F_[0][0][182],
F_[0][1][182],
F_[0][2][182],
F_[1][0][182],
F_[1][1][182],
F_[1][2][182],
F_[2][0][182],
F_[2][1][182],
F_[2][2][182],
F_[3][0][182],
F_[3][1][182],
F_[3][2][182],
F_[4][0][182],
F_[4][1][182],
F_[4][2][182],
F_[5][0][182],
F_[5][1][182],
F_[5][2][182],
F_[6][0][182],
F_[6][1][182],
F_[6][2][182],
F_[7][0][182],
F_[7][1][182],
F_[7][2][182],
F_[8][0][182],
F_[8][1][182],
F_[8][2][182],
F_[9][0][182],
F_[9][1][182],
F_[9][2][182],
F_[10][0][182],
F_[10][1][182],
F_[10][2][182],
F_[11][0][182],
F_[11][1][182],
F_[11][2][182],
F_[12][0][182],
F_[12][1][182],
F_[12][2][182],
F_[13][0][182],
F_[13][1][182],
F_[13][2][182],
F_[14][0][182],
F_[14][1][182],
F_[14][2][182],
F_[15][0][182],
F_[15][1][182],
F_[15][2][182],
F_[0][0][183],
F_[0][1][183],
F_[0][2][183],
F_[1][0][183],
F_[1][1][183],
F_[1][2][183],
F_[2][0][183],
F_[2][1][183],
F_[2][2][183],
F_[3][0][183],
F_[3][1][183],
F_[3][2][183],
F_[4][0][183],
F_[4][1][183],
F_[4][2][183],
F_[5][0][183],
F_[5][1][183],
F_[5][2][183],
F_[6][0][183],
F_[6][1][183],
F_[6][2][183],
F_[7][0][183],
F_[7][1][183],
F_[7][2][183],
F_[8][0][183],
F_[8][1][183],
F_[8][2][183],
F_[9][0][183],
F_[9][1][183],
F_[9][2][183],
F_[10][0][183],
F_[10][1][183],
F_[10][2][183],
F_[11][0][183],
F_[11][1][183],
F_[11][2][183],
F_[12][0][183],
F_[12][1][183],
F_[12][2][183],
F_[13][0][183],
F_[13][1][183],
F_[13][2][183],
F_[14][0][183],
F_[14][1][183],
F_[14][2][183],
F_[15][0][183],
F_[15][1][183],
F_[15][2][183],
F_[0][0][184],
F_[0][1][184],
F_[0][2][184],
F_[1][0][184],
F_[1][1][184],
F_[1][2][184],
F_[2][0][184],
F_[2][1][184],
F_[2][2][184],
F_[3][0][184],
F_[3][1][184],
F_[3][2][184],
F_[4][0][184],
F_[4][1][184],
F_[4][2][184],
F_[5][0][184],
F_[5][1][184],
F_[5][2][184],
F_[6][0][184],
F_[6][1][184],
F_[6][2][184],
F_[7][0][184],
F_[7][1][184],
F_[7][2][184],
F_[8][0][184],
F_[8][1][184],
F_[8][2][184],
F_[9][0][184],
F_[9][1][184],
F_[9][2][184],
F_[10][0][184],
F_[10][1][184],
F_[10][2][184],
F_[11][0][184],
F_[11][1][184],
F_[11][2][184],
F_[12][0][184],
F_[12][1][184],
F_[12][2][184],
F_[13][0][184],
F_[13][1][184],
F_[13][2][184],
F_[14][0][184],
F_[14][1][184],
F_[14][2][184],
F_[15][0][184],
F_[15][1][184],
F_[15][2][184],
F_[0][0][185],
F_[0][1][185],
F_[0][2][185],
F_[1][0][185],
F_[1][1][185],
F_[1][2][185],
F_[2][0][185],
F_[2][1][185],
F_[2][2][185],
F_[3][0][185],
F_[3][1][185],
F_[3][2][185],
F_[4][0][185],
F_[4][1][185],
F_[4][2][185],
F_[5][0][185],
F_[5][1][185],
F_[5][2][185],
F_[6][0][185],
F_[6][1][185],
F_[6][2][185],
F_[7][0][185],
F_[7][1][185],
F_[7][2][185],
F_[8][0][185],
F_[8][1][185],
F_[8][2][185],
F_[9][0][185],
F_[9][1][185],
F_[9][2][185],
F_[10][0][185],
F_[10][1][185],
F_[10][2][185],
F_[11][0][185],
F_[11][1][185],
F_[11][2][185],
F_[12][0][185],
F_[12][1][185],
F_[12][2][185],
F_[13][0][185],
F_[13][1][185],
F_[13][2][185],
F_[14][0][185],
F_[14][1][185],
F_[14][2][185],
F_[15][0][185],
F_[15][1][185],
F_[15][2][185],
F_[0][0][186],
F_[0][1][186],
F_[0][2][186],
F_[1][0][186],
F_[1][1][186],
F_[1][2][186],
F_[2][0][186],
F_[2][1][186],
F_[2][2][186],
F_[3][0][186],
F_[3][1][186],
F_[3][2][186],
F_[4][0][186],
F_[4][1][186],
F_[4][2][186],
F_[5][0][186],
F_[5][1][186],
F_[5][2][186],
F_[6][0][186],
F_[6][1][186],
F_[6][2][186],
F_[7][0][186],
F_[7][1][186],
F_[7][2][186],
F_[8][0][186],
F_[8][1][186],
F_[8][2][186],
F_[9][0][186],
F_[9][1][186],
F_[9][2][186],
F_[10][0][186],
F_[10][1][186],
F_[10][2][186],
F_[11][0][186],
F_[11][1][186],
F_[11][2][186],
F_[12][0][186],
F_[12][1][186],
F_[12][2][186],
F_[13][0][186],
F_[13][1][186],
F_[13][2][186],
F_[14][0][186],
F_[14][1][186],
F_[14][2][186],
F_[15][0][186],
F_[15][1][186],
F_[15][2][186],
F_[0][0][187],
F_[0][1][187],
F_[0][2][187],
F_[1][0][187],
F_[1][1][187],
F_[1][2][187],
F_[2][0][187],
F_[2][1][187],
F_[2][2][187],
F_[3][0][187],
F_[3][1][187],
F_[3][2][187],
F_[4][0][187],
F_[4][1][187],
F_[4][2][187],
F_[5][0][187],
F_[5][1][187],
F_[5][2][187],
F_[6][0][187],
F_[6][1][187],
F_[6][2][187],
F_[7][0][187],
F_[7][1][187],
F_[7][2][187],
F_[8][0][187],
F_[8][1][187],
F_[8][2][187],
F_[9][0][187],
F_[9][1][187],
F_[9][2][187],
F_[10][0][187],
F_[10][1][187],
F_[10][2][187],
F_[11][0][187],
F_[11][1][187],
F_[11][2][187],
F_[12][0][187],
F_[12][1][187],
F_[12][2][187],
F_[13][0][187],
F_[13][1][187],
F_[13][2][187],
F_[14][0][187],
F_[14][1][187],
F_[14][2][187],
F_[15][0][187],
F_[15][1][187],
F_[15][2][187],
F_[0][0][188],
F_[0][1][188],
F_[0][2][188],
F_[1][0][188],
F_[1][1][188],
F_[1][2][188],
F_[2][0][188],
F_[2][1][188],
F_[2][2][188],
F_[3][0][188],
F_[3][1][188],
F_[3][2][188],
F_[4][0][188],
F_[4][1][188],
F_[4][2][188],
F_[5][0][188],
F_[5][1][188],
F_[5][2][188],
F_[6][0][188],
F_[6][1][188],
F_[6][2][188],
F_[7][0][188],
F_[7][1][188],
F_[7][2][188],
F_[8][0][188],
F_[8][1][188],
F_[8][2][188],
F_[9][0][188],
F_[9][1][188],
F_[9][2][188],
F_[10][0][188],
F_[10][1][188],
F_[10][2][188],
F_[11][0][188],
F_[11][1][188],
F_[11][2][188],
F_[12][0][188],
F_[12][1][188],
F_[12][2][188],
F_[13][0][188],
F_[13][1][188],
F_[13][2][188],
F_[14][0][188],
F_[14][1][188],
F_[14][2][188],
F_[15][0][188],
F_[15][1][188],
F_[15][2][188],
F_[0][0][189],
F_[0][1][189],
F_[0][2][189],
F_[1][0][189],
F_[1][1][189],
F_[1][2][189],
F_[2][0][189],
F_[2][1][189],
F_[2][2][189],
F_[3][0][189],
F_[3][1][189],
F_[3][2][189],
F_[4][0][189],
F_[4][1][189],
F_[4][2][189],
F_[5][0][189],
F_[5][1][189],
F_[5][2][189],
F_[6][0][189],
F_[6][1][189],
F_[6][2][189],
F_[7][0][189],
F_[7][1][189],
F_[7][2][189],
F_[8][0][189],
F_[8][1][189],
F_[8][2][189],
F_[9][0][189],
F_[9][1][189],
F_[9][2][189],
F_[10][0][189],
F_[10][1][189],
F_[10][2][189],
F_[11][0][189],
F_[11][1][189],
F_[11][2][189],
F_[12][0][189],
F_[12][1][189],
F_[12][2][189],
F_[13][0][189],
F_[13][1][189],
F_[13][2][189],
F_[14][0][189],
F_[14][1][189],
F_[14][2][189],
F_[15][0][189],
F_[15][1][189],
F_[15][2][189],
F_[0][0][190],
F_[0][1][190],
F_[0][2][190],
F_[1][0][190],
F_[1][1][190],
F_[1][2][190],
F_[2][0][190],
F_[2][1][190],
F_[2][2][190],
F_[3][0][190],
F_[3][1][190],
F_[3][2][190],
F_[4][0][190],
F_[4][1][190],
F_[4][2][190],
F_[5][0][190],
F_[5][1][190],
F_[5][2][190],
F_[6][0][190],
F_[6][1][190],
F_[6][2][190],
F_[7][0][190],
F_[7][1][190],
F_[7][2][190],
F_[8][0][190],
F_[8][1][190],
F_[8][2][190],
F_[9][0][190],
F_[9][1][190],
F_[9][2][190],
F_[10][0][190],
F_[10][1][190],
F_[10][2][190],
F_[11][0][190],
F_[11][1][190],
F_[11][2][190],
F_[12][0][190],
F_[12][1][190],
F_[12][2][190],
F_[13][0][190],
F_[13][1][190],
F_[13][2][190],
F_[14][0][190],
F_[14][1][190],
F_[14][2][190],
F_[15][0][190],
F_[15][1][190],
F_[15][2][190],
F_[0][0][191],
F_[0][1][191],
F_[0][2][191],
F_[1][0][191],
F_[1][1][191],
F_[1][2][191],
F_[2][0][191],
F_[2][1][191],
F_[2][2][191],
F_[3][0][191],
F_[3][1][191],
F_[3][2][191],
F_[4][0][191],
F_[4][1][191],
F_[4][2][191],
F_[5][0][191],
F_[5][1][191],
F_[5][2][191],
F_[6][0][191],
F_[6][1][191],
F_[6][2][191],
F_[7][0][191],
F_[7][1][191],
F_[7][2][191],
F_[8][0][191],
F_[8][1][191],
F_[8][2][191],
F_[9][0][191],
F_[9][1][191],
F_[9][2][191],
F_[10][0][191],
F_[10][1][191],
F_[10][2][191],
F_[11][0][191],
F_[11][1][191],
F_[11][2][191],
F_[12][0][191],
F_[12][1][191],
F_[12][2][191],
F_[13][0][191],
F_[13][1][191],
F_[13][2][191],
F_[14][0][191],
F_[14][1][191],
F_[14][2][191],
F_[15][0][191],
F_[15][1][191],
F_[15][2][191],
F_[0][0][192],
F_[0][1][192],
F_[0][2][192],
F_[1][0][192],
F_[1][1][192],
F_[1][2][192],
F_[2][0][192],
F_[2][1][192],
F_[2][2][192],
F_[3][0][192],
F_[3][1][192],
F_[3][2][192],
F_[4][0][192],
F_[4][1][192],
F_[4][2][192],
F_[5][0][192],
F_[5][1][192],
F_[5][2][192],
F_[6][0][192],
F_[6][1][192],
F_[6][2][192],
F_[7][0][192],
F_[7][1][192],
F_[7][2][192],
F_[8][0][192],
F_[8][1][192],
F_[8][2][192],
F_[9][0][192],
F_[9][1][192],
F_[9][2][192],
F_[10][0][192],
F_[10][1][192],
F_[10][2][192],
F_[11][0][192],
F_[11][1][192],
F_[11][2][192],
F_[12][0][192],
F_[12][1][192],
F_[12][2][192],
F_[13][0][192],
F_[13][1][192],
F_[13][2][192],
F_[14][0][192],
F_[14][1][192],
F_[14][2][192],
F_[15][0][192],
F_[15][1][192],
F_[15][2][192],
F_[0][0][193],
F_[0][1][193],
F_[0][2][193],
F_[1][0][193],
F_[1][1][193],
F_[1][2][193],
F_[2][0][193],
F_[2][1][193],
F_[2][2][193],
F_[3][0][193],
F_[3][1][193],
F_[3][2][193],
F_[4][0][193],
F_[4][1][193],
F_[4][2][193],
F_[5][0][193],
F_[5][1][193],
F_[5][2][193],
F_[6][0][193],
F_[6][1][193],
F_[6][2][193],
F_[7][0][193],
F_[7][1][193],
F_[7][2][193],
F_[8][0][193],
F_[8][1][193],
F_[8][2][193],
F_[9][0][193],
F_[9][1][193],
F_[9][2][193],
F_[10][0][193],
F_[10][1][193],
F_[10][2][193],
F_[11][0][193],
F_[11][1][193],
F_[11][2][193],
F_[12][0][193],
F_[12][1][193],
F_[12][2][193],
F_[13][0][193],
F_[13][1][193],
F_[13][2][193],
F_[14][0][193],
F_[14][1][193],
F_[14][2][193],
F_[15][0][193],
F_[15][1][193],
F_[15][2][193],
F_[0][0][194],
F_[0][1][194],
F_[0][2][194],
F_[1][0][194],
F_[1][1][194],
F_[1][2][194],
F_[2][0][194],
F_[2][1][194],
F_[2][2][194],
F_[3][0][194],
F_[3][1][194],
F_[3][2][194],
F_[4][0][194],
F_[4][1][194],
F_[4][2][194],
F_[5][0][194],
F_[5][1][194],
F_[5][2][194],
F_[6][0][194],
F_[6][1][194],
F_[6][2][194],
F_[7][0][194],
F_[7][1][194],
F_[7][2][194],
F_[8][0][194],
F_[8][1][194],
F_[8][2][194],
F_[9][0][194],
F_[9][1][194],
F_[9][2][194],
F_[10][0][194],
F_[10][1][194],
F_[10][2][194],
F_[11][0][194],
F_[11][1][194],
F_[11][2][194],
F_[12][0][194],
F_[12][1][194],
F_[12][2][194],
F_[13][0][194],
F_[13][1][194],
F_[13][2][194],
F_[14][0][194],
F_[14][1][194],
F_[14][2][194],
F_[15][0][194],
F_[15][1][194],
F_[15][2][194],
F_[0][0][195],
F_[0][1][195],
F_[0][2][195],
F_[1][0][195],
F_[1][1][195],
F_[1][2][195],
F_[2][0][195],
F_[2][1][195],
F_[2][2][195],
F_[3][0][195],
F_[3][1][195],
F_[3][2][195],
F_[4][0][195],
F_[4][1][195],
F_[4][2][195],
F_[5][0][195],
F_[5][1][195],
F_[5][2][195],
F_[6][0][195],
F_[6][1][195],
F_[6][2][195],
F_[7][0][195],
F_[7][1][195],
F_[7][2][195],
F_[8][0][195],
F_[8][1][195],
F_[8][2][195],
F_[9][0][195],
F_[9][1][195],
F_[9][2][195],
F_[10][0][195],
F_[10][1][195],
F_[10][2][195],
F_[11][0][195],
F_[11][1][195],
F_[11][2][195],
F_[12][0][195],
F_[12][1][195],
F_[12][2][195],
F_[13][0][195],
F_[13][1][195],
F_[13][2][195],
F_[14][0][195],
F_[14][1][195],
F_[14][2][195],
F_[15][0][195],
F_[15][1][195],
F_[15][2][195],
F_[0][0][196],
F_[0][1][196],
F_[0][2][196],
F_[1][0][196],
F_[1][1][196],
F_[1][2][196],
F_[2][0][196],
F_[2][1][196],
F_[2][2][196],
F_[3][0][196],
F_[3][1][196],
F_[3][2][196],
F_[4][0][196],
F_[4][1][196],
F_[4][2][196],
F_[5][0][196],
F_[5][1][196],
F_[5][2][196],
F_[6][0][196],
F_[6][1][196],
F_[6][2][196],
F_[7][0][196],
F_[7][1][196],
F_[7][2][196],
F_[8][0][196],
F_[8][1][196],
F_[8][2][196],
F_[9][0][196],
F_[9][1][196],
F_[9][2][196],
F_[10][0][196],
F_[10][1][196],
F_[10][2][196],
F_[11][0][196],
F_[11][1][196],
F_[11][2][196],
F_[12][0][196],
F_[12][1][196],
F_[12][2][196],
F_[13][0][196],
F_[13][1][196],
F_[13][2][196],
F_[14][0][196],
F_[14][1][196],
F_[14][2][196],
F_[15][0][196],
F_[15][1][196],
F_[15][2][196],
F_[0][0][197],
F_[0][1][197],
F_[0][2][197],
F_[1][0][197],
F_[1][1][197],
F_[1][2][197],
F_[2][0][197],
F_[2][1][197],
F_[2][2][197],
F_[3][0][197],
F_[3][1][197],
F_[3][2][197],
F_[4][0][197],
F_[4][1][197],
F_[4][2][197],
F_[5][0][197],
F_[5][1][197],
F_[5][2][197],
F_[6][0][197],
F_[6][1][197],
F_[6][2][197],
F_[7][0][197],
F_[7][1][197],
F_[7][2][197],
F_[8][0][197],
F_[8][1][197],
F_[8][2][197],
F_[9][0][197],
F_[9][1][197],
F_[9][2][197],
F_[10][0][197],
F_[10][1][197],
F_[10][2][197],
F_[11][0][197],
F_[11][1][197],
F_[11][2][197],
F_[12][0][197],
F_[12][1][197],
F_[12][2][197],
F_[13][0][197],
F_[13][1][197],
F_[13][2][197],
F_[14][0][197],
F_[14][1][197],
F_[14][2][197],
F_[15][0][197],
F_[15][1][197],
F_[15][2][197],
F_[0][0][198],
F_[0][1][198],
F_[0][2][198],
F_[1][0][198],
F_[1][1][198],
F_[1][2][198],
F_[2][0][198],
F_[2][1][198],
F_[2][2][198],
F_[3][0][198],
F_[3][1][198],
F_[3][2][198],
F_[4][0][198],
F_[4][1][198],
F_[4][2][198],
F_[5][0][198],
F_[5][1][198],
F_[5][2][198],
F_[6][0][198],
F_[6][1][198],
F_[6][2][198],
F_[7][0][198],
F_[7][1][198],
F_[7][2][198],
F_[8][0][198],
F_[8][1][198],
F_[8][2][198],
F_[9][0][198],
F_[9][1][198],
F_[9][2][198],
F_[10][0][198],
F_[10][1][198],
F_[10][2][198],
F_[11][0][198],
F_[11][1][198],
F_[11][2][198],
F_[12][0][198],
F_[12][1][198],
F_[12][2][198],
F_[13][0][198],
F_[13][1][198],
F_[13][2][198],
F_[14][0][198],
F_[14][1][198],
F_[14][2][198],
F_[15][0][198],
F_[15][1][198],
F_[15][2][198],
F_[0][0][199],
F_[0][1][199],
F_[0][2][199],
F_[1][0][199],
F_[1][1][199],
F_[1][2][199],
F_[2][0][199],
F_[2][1][199],
F_[2][2][199],
F_[3][0][199],
F_[3][1][199],
F_[3][2][199],
F_[4][0][199],
F_[4][1][199],
F_[4][2][199],
F_[5][0][199],
F_[5][1][199],
F_[5][2][199],
F_[6][0][199],
F_[6][1][199],
F_[6][2][199],
F_[7][0][199],
F_[7][1][199],
F_[7][2][199],
F_[8][0][199],
F_[8][1][199],
F_[8][2][199],
F_[9][0][199],
F_[9][1][199],
F_[9][2][199],
F_[10][0][199],
F_[10][1][199],
F_[10][2][199],
F_[11][0][199],
F_[11][1][199],
F_[11][2][199],
F_[12][0][199],
F_[12][1][199],
F_[12][2][199],
F_[13][0][199],
F_[13][1][199],
F_[13][2][199],
F_[14][0][199],
F_[14][1][199],
F_[14][2][199],
F_[15][0][199],
F_[15][1][199],
F_[15][2][199],
F_[0][0][200],
F_[0][1][200],
F_[0][2][200],
F_[1][0][200],
F_[1][1][200],
F_[1][2][200],
F_[2][0][200],
F_[2][1][200],
F_[2][2][200],
F_[3][0][200],
F_[3][1][200],
F_[3][2][200],
F_[4][0][200],
F_[4][1][200],
F_[4][2][200],
F_[5][0][200],
F_[5][1][200],
F_[5][2][200],
F_[6][0][200],
F_[6][1][200],
F_[6][2][200],
F_[7][0][200],
F_[7][1][200],
F_[7][2][200],
F_[8][0][200],
F_[8][1][200],
F_[8][2][200],
F_[9][0][200],
F_[9][1][200],
F_[9][2][200],
F_[10][0][200],
F_[10][1][200],
F_[10][2][200],
F_[11][0][200],
F_[11][1][200],
F_[11][2][200],
F_[12][0][200],
F_[12][1][200],
F_[12][2][200],
F_[13][0][200],
F_[13][1][200],
F_[13][2][200],
F_[14][0][200],
F_[14][1][200],
F_[14][2][200],
F_[15][0][200],
F_[15][1][200],
F_[15][2][200],
F_[0][0][201],
F_[0][1][201],
F_[0][2][201],
F_[1][0][201],
F_[1][1][201],
F_[1][2][201],
F_[2][0][201],
F_[2][1][201],
F_[2][2][201],
F_[3][0][201],
F_[3][1][201],
F_[3][2][201],
F_[4][0][201],
F_[4][1][201],
F_[4][2][201],
F_[5][0][201],
F_[5][1][201],
F_[5][2][201],
F_[6][0][201],
F_[6][1][201],
F_[6][2][201],
F_[7][0][201],
F_[7][1][201],
F_[7][2][201],
F_[8][0][201],
F_[8][1][201],
F_[8][2][201],
F_[9][0][201],
F_[9][1][201],
F_[9][2][201],
F_[10][0][201],
F_[10][1][201],
F_[10][2][201],
F_[11][0][201],
F_[11][1][201],
F_[11][2][201],
F_[12][0][201],
F_[12][1][201],
F_[12][2][201],
F_[13][0][201],
F_[13][1][201],
F_[13][2][201],
F_[14][0][201],
F_[14][1][201],
F_[14][2][201],
F_[15][0][201],
F_[15][1][201],
F_[15][2][201],
F_[0][0][202],
F_[0][1][202],
F_[0][2][202],
F_[1][0][202],
F_[1][1][202],
F_[1][2][202],
F_[2][0][202],
F_[2][1][202],
F_[2][2][202],
F_[3][0][202],
F_[3][1][202],
F_[3][2][202],
F_[4][0][202],
F_[4][1][202],
F_[4][2][202],
F_[5][0][202],
F_[5][1][202],
F_[5][2][202],
F_[6][0][202],
F_[6][1][202],
F_[6][2][202],
F_[7][0][202],
F_[7][1][202],
F_[7][2][202],
F_[8][0][202],
F_[8][1][202],
F_[8][2][202],
F_[9][0][202],
F_[9][1][202],
F_[9][2][202],
F_[10][0][202],
F_[10][1][202],
F_[10][2][202],
F_[11][0][202],
F_[11][1][202],
F_[11][2][202],
F_[12][0][202],
F_[12][1][202],
F_[12][2][202],
F_[13][0][202],
F_[13][1][202],
F_[13][2][202],
F_[14][0][202],
F_[14][1][202],
F_[14][2][202],
F_[15][0][202],
F_[15][1][202],
F_[15][2][202],
F_[0][0][203],
F_[0][1][203],
F_[0][2][203],
F_[1][0][203],
F_[1][1][203],
F_[1][2][203],
F_[2][0][203],
F_[2][1][203],
F_[2][2][203],
F_[3][0][203],
F_[3][1][203],
F_[3][2][203],
F_[4][0][203],
F_[4][1][203],
F_[4][2][203],
F_[5][0][203],
F_[5][1][203],
F_[5][2][203],
F_[6][0][203],
F_[6][1][203],
F_[6][2][203],
F_[7][0][203],
F_[7][1][203],
F_[7][2][203],
F_[8][0][203],
F_[8][1][203],
F_[8][2][203],
F_[9][0][203],
F_[9][1][203],
F_[9][2][203],
F_[10][0][203],
F_[10][1][203],
F_[10][2][203],
F_[11][0][203],
F_[11][1][203],
F_[11][2][203],
F_[12][0][203],
F_[12][1][203],
F_[12][2][203],
F_[13][0][203],
F_[13][1][203],
F_[13][2][203],
F_[14][0][203],
F_[14][1][203],
F_[14][2][203],
F_[15][0][203],
F_[15][1][203],
F_[15][2][203],
F_[0][0][204],
F_[0][1][204],
F_[0][2][204],
F_[1][0][204],
F_[1][1][204],
F_[1][2][204],
F_[2][0][204],
F_[2][1][204],
F_[2][2][204],
F_[3][0][204],
F_[3][1][204],
F_[3][2][204],
F_[4][0][204],
F_[4][1][204],
F_[4][2][204],
F_[5][0][204],
F_[5][1][204],
F_[5][2][204],
F_[6][0][204],
F_[6][1][204],
F_[6][2][204],
F_[7][0][204],
F_[7][1][204],
F_[7][2][204],
F_[8][0][204],
F_[8][1][204],
F_[8][2][204],
F_[9][0][204],
F_[9][1][204],
F_[9][2][204],
F_[10][0][204],
F_[10][1][204],
F_[10][2][204],
F_[11][0][204],
F_[11][1][204],
F_[11][2][204],
F_[12][0][204],
F_[12][1][204],
F_[12][2][204],
F_[13][0][204],
F_[13][1][204],
F_[13][2][204],
F_[14][0][204],
F_[14][1][204],
F_[14][2][204],
F_[15][0][204],
F_[15][1][204],
F_[15][2][204],
F_[0][0][205],
F_[0][1][205],
F_[0][2][205],
F_[1][0][205],
F_[1][1][205],
F_[1][2][205],
F_[2][0][205],
F_[2][1][205],
F_[2][2][205],
F_[3][0][205],
F_[3][1][205],
F_[3][2][205],
F_[4][0][205],
F_[4][1][205],
F_[4][2][205],
F_[5][0][205],
F_[5][1][205],
F_[5][2][205],
F_[6][0][205],
F_[6][1][205],
F_[6][2][205],
F_[7][0][205],
F_[7][1][205],
F_[7][2][205],
F_[8][0][205],
F_[8][1][205],
F_[8][2][205],
F_[9][0][205],
F_[9][1][205],
F_[9][2][205],
F_[10][0][205],
F_[10][1][205],
F_[10][2][205],
F_[11][0][205],
F_[11][1][205],
F_[11][2][205],
F_[12][0][205],
F_[12][1][205],
F_[12][2][205],
F_[13][0][205],
F_[13][1][205],
F_[13][2][205],
F_[14][0][205],
F_[14][1][205],
F_[14][2][205],
F_[15][0][205],
F_[15][1][205],
F_[15][2][205],
F_[0][0][206],
F_[0][1][206],
F_[0][2][206],
F_[1][0][206],
F_[1][1][206],
F_[1][2][206],
F_[2][0][206],
F_[2][1][206],
F_[2][2][206],
F_[3][0][206],
F_[3][1][206],
F_[3][2][206],
F_[4][0][206],
F_[4][1][206],
F_[4][2][206],
F_[5][0][206],
F_[5][1][206],
F_[5][2][206],
F_[6][0][206],
F_[6][1][206],
F_[6][2][206],
F_[7][0][206],
F_[7][1][206],
F_[7][2][206],
F_[8][0][206],
F_[8][1][206],
F_[8][2][206],
F_[9][0][206],
F_[9][1][206],
F_[9][2][206],
F_[10][0][206],
F_[10][1][206],
F_[10][2][206],
F_[11][0][206],
F_[11][1][206],
F_[11][2][206],
F_[12][0][206],
F_[12][1][206],
F_[12][2][206],
F_[13][0][206],
F_[13][1][206],
F_[13][2][206],
F_[14][0][206],
F_[14][1][206],
F_[14][2][206],
F_[15][0][206],
F_[15][1][206],
F_[15][2][206],
F_[0][0][207],
F_[0][1][207],
F_[0][2][207],
F_[1][0][207],
F_[1][1][207],
F_[1][2][207],
F_[2][0][207],
F_[2][1][207],
F_[2][2][207],
F_[3][0][207],
F_[3][1][207],
F_[3][2][207],
F_[4][0][207],
F_[4][1][207],
F_[4][2][207],
F_[5][0][207],
F_[5][1][207],
F_[5][2][207],
F_[6][0][207],
F_[6][1][207],
F_[6][2][207],
F_[7][0][207],
F_[7][1][207],
F_[7][2][207],
F_[8][0][207],
F_[8][1][207],
F_[8][2][207],
F_[9][0][207],
F_[9][1][207],
F_[9][2][207],
F_[10][0][207],
F_[10][1][207],
F_[10][2][207],
F_[11][0][207],
F_[11][1][207],
F_[11][2][207],
F_[12][0][207],
F_[12][1][207],
F_[12][2][207],
F_[13][0][207],
F_[13][1][207],
F_[13][2][207],
F_[14][0][207],
F_[14][1][207],
F_[14][2][207],
F_[15][0][207],
F_[15][1][207],
F_[15][2][207],
F_[0][0][208],
F_[0][1][208],
F_[0][2][208],
F_[1][0][208],
F_[1][1][208],
F_[1][2][208],
F_[2][0][208],
F_[2][1][208],
F_[2][2][208],
F_[3][0][208],
F_[3][1][208],
F_[3][2][208],
F_[4][0][208],
F_[4][1][208],
F_[4][2][208],
F_[5][0][208],
F_[5][1][208],
F_[5][2][208],
F_[6][0][208],
F_[6][1][208],
F_[6][2][208],
F_[7][0][208],
F_[7][1][208],
F_[7][2][208],
F_[8][0][208],
F_[8][1][208],
F_[8][2][208],
F_[9][0][208],
F_[9][1][208],
F_[9][2][208],
F_[10][0][208],
F_[10][1][208],
F_[10][2][208],
F_[11][0][208],
F_[11][1][208],
F_[11][2][208],
F_[12][0][208],
F_[12][1][208],
F_[12][2][208],
F_[13][0][208],
F_[13][1][208],
F_[13][2][208],
F_[14][0][208],
F_[14][1][208],
F_[14][2][208],
F_[15][0][208],
F_[15][1][208],
F_[15][2][208],
F_[0][0][209],
F_[0][1][209],
F_[0][2][209],
F_[1][0][209],
F_[1][1][209],
F_[1][2][209],
F_[2][0][209],
F_[2][1][209],
F_[2][2][209],
F_[3][0][209],
F_[3][1][209],
F_[3][2][209],
F_[4][0][209],
F_[4][1][209],
F_[4][2][209],
F_[5][0][209],
F_[5][1][209],
F_[5][2][209],
F_[6][0][209],
F_[6][1][209],
F_[6][2][209],
F_[7][0][209],
F_[7][1][209],
F_[7][2][209],
F_[8][0][209],
F_[8][1][209],
F_[8][2][209],
F_[9][0][209],
F_[9][1][209],
F_[9][2][209],
F_[10][0][209],
F_[10][1][209],
F_[10][2][209],
F_[11][0][209],
F_[11][1][209],
F_[11][2][209],
F_[12][0][209],
F_[12][1][209],
F_[12][2][209],
F_[13][0][209],
F_[13][1][209],
F_[13][2][209],
F_[14][0][209],
F_[14][1][209],
F_[14][2][209],
F_[15][0][209],
F_[15][1][209],
F_[15][2][209],
F_[0][0][210],
F_[0][1][210],
F_[0][2][210],
F_[1][0][210],
F_[1][1][210],
F_[1][2][210],
F_[2][0][210],
F_[2][1][210],
F_[2][2][210],
F_[3][0][210],
F_[3][1][210],
F_[3][2][210],
F_[4][0][210],
F_[4][1][210],
F_[4][2][210],
F_[5][0][210],
F_[5][1][210],
F_[5][2][210],
F_[6][0][210],
F_[6][1][210],
F_[6][2][210],
F_[7][0][210],
F_[7][1][210],
F_[7][2][210],
F_[8][0][210],
F_[8][1][210],
F_[8][2][210],
F_[9][0][210],
F_[9][1][210],
F_[9][2][210],
F_[10][0][210],
F_[10][1][210],
F_[10][2][210],
F_[11][0][210],
F_[11][1][210],
F_[11][2][210],
F_[12][0][210],
F_[12][1][210],
F_[12][2][210],
F_[13][0][210],
F_[13][1][210],
F_[13][2][210],
F_[14][0][210],
F_[14][1][210],
F_[14][2][210],
F_[15][0][210],
F_[15][1][210],
F_[15][2][210],
F_[0][0][211],
F_[0][1][211],
F_[0][2][211],
F_[1][0][211],
F_[1][1][211],
F_[1][2][211],
F_[2][0][211],
F_[2][1][211],
F_[2][2][211],
F_[3][0][211],
F_[3][1][211],
F_[3][2][211],
F_[4][0][211],
F_[4][1][211],
F_[4][2][211],
F_[5][0][211],
F_[5][1][211],
F_[5][2][211],
F_[6][0][211],
F_[6][1][211],
F_[6][2][211],
F_[7][0][211],
F_[7][1][211],
F_[7][2][211],
F_[8][0][211],
F_[8][1][211],
F_[8][2][211],
F_[9][0][211],
F_[9][1][211],
F_[9][2][211],
F_[10][0][211],
F_[10][1][211],
F_[10][2][211],
F_[11][0][211],
F_[11][1][211],
F_[11][2][211],
F_[12][0][211],
F_[12][1][211],
F_[12][2][211],
F_[13][0][211],
F_[13][1][211],
F_[13][2][211],
F_[14][0][211],
F_[14][1][211],
F_[14][2][211],
F_[15][0][211],
F_[15][1][211],
F_[15][2][211],
F_[0][0][212],
F_[0][1][212],
F_[0][2][212],
F_[1][0][212],
F_[1][1][212],
F_[1][2][212],
F_[2][0][212],
F_[2][1][212],
F_[2][2][212],
F_[3][0][212],
F_[3][1][212],
F_[3][2][212],
F_[4][0][212],
F_[4][1][212],
F_[4][2][212],
F_[5][0][212],
F_[5][1][212],
F_[5][2][212],
F_[6][0][212],
F_[6][1][212],
F_[6][2][212],
F_[7][0][212],
F_[7][1][212],
F_[7][2][212],
F_[8][0][212],
F_[8][1][212],
F_[8][2][212],
F_[9][0][212],
F_[9][1][212],
F_[9][2][212],
F_[10][0][212],
F_[10][1][212],
F_[10][2][212],
F_[11][0][212],
F_[11][1][212],
F_[11][2][212],
F_[12][0][212],
F_[12][1][212],
F_[12][2][212],
F_[13][0][212],
F_[13][1][212],
F_[13][2][212],
F_[14][0][212],
F_[14][1][212],
F_[14][2][212],
F_[15][0][212],
F_[15][1][212],
F_[15][2][212],
F_[0][0][213],
F_[0][1][213],
F_[0][2][213],
F_[1][0][213],
F_[1][1][213],
F_[1][2][213],
F_[2][0][213],
F_[2][1][213],
F_[2][2][213],
F_[3][0][213],
F_[3][1][213],
F_[3][2][213],
F_[4][0][213],
F_[4][1][213],
F_[4][2][213],
F_[5][0][213],
F_[5][1][213],
F_[5][2][213],
F_[6][0][213],
F_[6][1][213],
F_[6][2][213],
F_[7][0][213],
F_[7][1][213],
F_[7][2][213],
F_[8][0][213],
F_[8][1][213],
F_[8][2][213],
F_[9][0][213],
F_[9][1][213],
F_[9][2][213],
F_[10][0][213],
F_[10][1][213],
F_[10][2][213],
F_[11][0][213],
F_[11][1][213],
F_[11][2][213],
F_[12][0][213],
F_[12][1][213],
F_[12][2][213],
F_[13][0][213],
F_[13][1][213],
F_[13][2][213],
F_[14][0][213],
F_[14][1][213],
F_[14][2][213],
F_[15][0][213],
F_[15][1][213],
F_[15][2][213],
F_[0][0][214],
F_[0][1][214],
F_[0][2][214],
F_[1][0][214],
F_[1][1][214],
F_[1][2][214],
F_[2][0][214],
F_[2][1][214],
F_[2][2][214],
F_[3][0][214],
F_[3][1][214],
F_[3][2][214],
F_[4][0][214],
F_[4][1][214],
F_[4][2][214],
F_[5][0][214],
F_[5][1][214],
F_[5][2][214],
F_[6][0][214],
F_[6][1][214],
F_[6][2][214],
F_[7][0][214],
F_[7][1][214],
F_[7][2][214],
F_[8][0][214],
F_[8][1][214],
F_[8][2][214],
F_[9][0][214],
F_[9][1][214],
F_[9][2][214],
F_[10][0][214],
F_[10][1][214],
F_[10][2][214],
F_[11][0][214],
F_[11][1][214],
F_[11][2][214],
F_[12][0][214],
F_[12][1][214],
F_[12][2][214],
F_[13][0][214],
F_[13][1][214],
F_[13][2][214],
F_[14][0][214],
F_[14][1][214],
F_[14][2][214],
F_[15][0][214],
F_[15][1][214],
F_[15][2][214],
F_[0][0][215],
F_[0][1][215],
F_[0][2][215],
F_[1][0][215],
F_[1][1][215],
F_[1][2][215],
F_[2][0][215],
F_[2][1][215],
F_[2][2][215],
F_[3][0][215],
F_[3][1][215],
F_[3][2][215],
F_[4][0][215],
F_[4][1][215],
F_[4][2][215],
F_[5][0][215],
F_[5][1][215],
F_[5][2][215],
F_[6][0][215],
F_[6][1][215],
F_[6][2][215],
F_[7][0][215],
F_[7][1][215],
F_[7][2][215],
F_[8][0][215],
F_[8][1][215],
F_[8][2][215],
F_[9][0][215],
F_[9][1][215],
F_[9][2][215],
F_[10][0][215],
F_[10][1][215],
F_[10][2][215],
F_[11][0][215],
F_[11][1][215],
F_[11][2][215],
F_[12][0][215],
F_[12][1][215],
F_[12][2][215],
F_[13][0][215],
F_[13][1][215],
F_[13][2][215],
F_[14][0][215],
F_[14][1][215],
F_[14][2][215],
F_[15][0][215],
F_[15][1][215],
F_[15][2][215],
F_[0][0][216],
F_[0][1][216],
F_[0][2][216],
F_[1][0][216],
F_[1][1][216],
F_[1][2][216],
F_[2][0][216],
F_[2][1][216],
F_[2][2][216],
F_[3][0][216],
F_[3][1][216],
F_[3][2][216],
F_[4][0][216],
F_[4][1][216],
F_[4][2][216],
F_[5][0][216],
F_[5][1][216],
F_[5][2][216],
F_[6][0][216],
F_[6][1][216],
F_[6][2][216],
F_[7][0][216],
F_[7][1][216],
F_[7][2][216],
F_[8][0][216],
F_[8][1][216],
F_[8][2][216],
F_[9][0][216],
F_[9][1][216],
F_[9][2][216],
F_[10][0][216],
F_[10][1][216],
F_[10][2][216],
F_[11][0][216],
F_[11][1][216],
F_[11][2][216],
F_[12][0][216],
F_[12][1][216],
F_[12][2][216],
F_[13][0][216],
F_[13][1][216],
F_[13][2][216],
F_[14][0][216],
F_[14][1][216],
F_[14][2][216],
F_[15][0][216],
F_[15][1][216],
F_[15][2][216],
F_[0][0][217],
F_[0][1][217],
F_[0][2][217],
F_[1][0][217],
F_[1][1][217],
F_[1][2][217],
F_[2][0][217],
F_[2][1][217],
F_[2][2][217],
F_[3][0][217],
F_[3][1][217],
F_[3][2][217],
F_[4][0][217],
F_[4][1][217],
F_[4][2][217],
F_[5][0][217],
F_[5][1][217],
F_[5][2][217],
F_[6][0][217],
F_[6][1][217],
F_[6][2][217],
F_[7][0][217],
F_[7][1][217],
F_[7][2][217],
F_[8][0][217],
F_[8][1][217],
F_[8][2][217],
F_[9][0][217],
F_[9][1][217],
F_[9][2][217],
F_[10][0][217],
F_[10][1][217],
F_[10][2][217],
F_[11][0][217],
F_[11][1][217],
F_[11][2][217],
F_[12][0][217],
F_[12][1][217],
F_[12][2][217],
F_[13][0][217],
F_[13][1][217],
F_[13][2][217],
F_[14][0][217],
F_[14][1][217],
F_[14][2][217],
F_[15][0][217],
F_[15][1][217],
F_[15][2][217],
F_[0][0][218],
F_[0][1][218],
F_[0][2][218],
F_[1][0][218],
F_[1][1][218],
F_[1][2][218],
F_[2][0][218],
F_[2][1][218],
F_[2][2][218],
F_[3][0][218],
F_[3][1][218],
F_[3][2][218],
F_[4][0][218],
F_[4][1][218],
F_[4][2][218],
F_[5][0][218],
F_[5][1][218],
F_[5][2][218],
F_[6][0][218],
F_[6][1][218],
F_[6][2][218],
F_[7][0][218],
F_[7][1][218],
F_[7][2][218],
F_[8][0][218],
F_[8][1][218],
F_[8][2][218],
F_[9][0][218],
F_[9][1][218],
F_[9][2][218],
F_[10][0][218],
F_[10][1][218],
F_[10][2][218],
F_[11][0][218],
F_[11][1][218],
F_[11][2][218],
F_[12][0][218],
F_[12][1][218],
F_[12][2][218],
F_[13][0][218],
F_[13][1][218],
F_[13][2][218],
F_[14][0][218],
F_[14][1][218],
F_[14][2][218],
F_[15][0][218],
F_[15][1][218],
F_[15][2][218],
F_[0][0][219],
F_[0][1][219],
F_[0][2][219],
F_[1][0][219],
F_[1][1][219],
F_[1][2][219],
F_[2][0][219],
F_[2][1][219],
F_[2][2][219],
F_[3][0][219],
F_[3][1][219],
F_[3][2][219],
F_[4][0][219],
F_[4][1][219],
F_[4][2][219],
F_[5][0][219],
F_[5][1][219],
F_[5][2][219],
F_[6][0][219],
F_[6][1][219],
F_[6][2][219],
F_[7][0][219],
F_[7][1][219],
F_[7][2][219],
F_[8][0][219],
F_[8][1][219],
F_[8][2][219],
F_[9][0][219],
F_[9][1][219],
F_[9][2][219],
F_[10][0][219],
F_[10][1][219],
F_[10][2][219],
F_[11][0][219],
F_[11][1][219],
F_[11][2][219],
F_[12][0][219],
F_[12][1][219],
F_[12][2][219],
F_[13][0][219],
F_[13][1][219],
F_[13][2][219],
F_[14][0][219],
F_[14][1][219],
F_[14][2][219],
F_[15][0][219],
F_[15][1][219],
F_[15][2][219],
F_[0][0][220],
F_[0][1][220],
F_[0][2][220],
F_[1][0][220],
F_[1][1][220],
F_[1][2][220],
F_[2][0][220],
F_[2][1][220],
F_[2][2][220],
F_[3][0][220],
F_[3][1][220],
F_[3][2][220],
F_[4][0][220],
F_[4][1][220],
F_[4][2][220],
F_[5][0][220],
F_[5][1][220],
F_[5][2][220],
F_[6][0][220],
F_[6][1][220],
F_[6][2][220],
F_[7][0][220],
F_[7][1][220],
F_[7][2][220],
F_[8][0][220],
F_[8][1][220],
F_[8][2][220],
F_[9][0][220],
F_[9][1][220],
F_[9][2][220],
F_[10][0][220],
F_[10][1][220],
F_[10][2][220],
F_[11][0][220],
F_[11][1][220],
F_[11][2][220],
F_[12][0][220],
F_[12][1][220],
F_[12][2][220],
F_[13][0][220],
F_[13][1][220],
F_[13][2][220],
F_[14][0][220],
F_[14][1][220],
F_[14][2][220],
F_[15][0][220],
F_[15][1][220],
F_[15][2][220],
F_[0][0][221],
F_[0][1][221],
F_[0][2][221],
F_[1][0][221],
F_[1][1][221],
F_[1][2][221],
F_[2][0][221],
F_[2][1][221],
F_[2][2][221],
F_[3][0][221],
F_[3][1][221],
F_[3][2][221],
F_[4][0][221],
F_[4][1][221],
F_[4][2][221],
F_[5][0][221],
F_[5][1][221],
F_[5][2][221],
F_[6][0][221],
F_[6][1][221],
F_[6][2][221],
F_[7][0][221],
F_[7][1][221],
F_[7][2][221],
F_[8][0][221],
F_[8][1][221],
F_[8][2][221],
F_[9][0][221],
F_[9][1][221],
F_[9][2][221],
F_[10][0][221],
F_[10][1][221],
F_[10][2][221],
F_[11][0][221],
F_[11][1][221],
F_[11][2][221],
F_[12][0][221],
F_[12][1][221],
F_[12][2][221],
F_[13][0][221],
F_[13][1][221],
F_[13][2][221],
F_[14][0][221],
F_[14][1][221],
F_[14][2][221],
F_[15][0][221],
F_[15][1][221],
F_[15][2][221],
F_[0][0][222],
F_[0][1][222],
F_[0][2][222],
F_[1][0][222],
F_[1][1][222],
F_[1][2][222],
F_[2][0][222],
F_[2][1][222],
F_[2][2][222],
F_[3][0][222],
F_[3][1][222],
F_[3][2][222],
F_[4][0][222],
F_[4][1][222],
F_[4][2][222],
F_[5][0][222],
F_[5][1][222],
F_[5][2][222],
F_[6][0][222],
F_[6][1][222],
F_[6][2][222],
F_[7][0][222],
F_[7][1][222],
F_[7][2][222],
F_[8][0][222],
F_[8][1][222],
F_[8][2][222],
F_[9][0][222],
F_[9][1][222],
F_[9][2][222],
F_[10][0][222],
F_[10][1][222],
F_[10][2][222],
F_[11][0][222],
F_[11][1][222],
F_[11][2][222],
F_[12][0][222],
F_[12][1][222],
F_[12][2][222],
F_[13][0][222],
F_[13][1][222],
F_[13][2][222],
F_[14][0][222],
F_[14][1][222],
F_[14][2][222],
F_[15][0][222],
F_[15][1][222],
F_[15][2][222],
F_[0][0][223],
F_[0][1][223],
F_[0][2][223],
F_[1][0][223],
F_[1][1][223],
F_[1][2][223],
F_[2][0][223],
F_[2][1][223],
F_[2][2][223],
F_[3][0][223],
F_[3][1][223],
F_[3][2][223],
F_[4][0][223],
F_[4][1][223],
F_[4][2][223],
F_[5][0][223],
F_[5][1][223],
F_[5][2][223],
F_[6][0][223],
F_[6][1][223],
F_[6][2][223],
F_[7][0][223],
F_[7][1][223],
F_[7][2][223],
F_[8][0][223],
F_[8][1][223],
F_[8][2][223],
F_[9][0][223],
F_[9][1][223],
F_[9][2][223],
F_[10][0][223],
F_[10][1][223],
F_[10][2][223],
F_[11][0][223],
F_[11][1][223],
F_[11][2][223],
F_[12][0][223],
F_[12][1][223],
F_[12][2][223],
F_[13][0][223],
F_[13][1][223],
F_[13][2][223],
F_[14][0][223],
F_[14][1][223],
F_[14][2][223],
F_[15][0][223],
F_[15][1][223],
F_[15][2][223],
F_[0][0][224],
F_[0][1][224],
F_[0][2][224],
F_[1][0][224],
F_[1][1][224],
F_[1][2][224],
F_[2][0][224],
F_[2][1][224],
F_[2][2][224],
F_[3][0][224],
F_[3][1][224],
F_[3][2][224],
F_[4][0][224],
F_[4][1][224],
F_[4][2][224],
F_[5][0][224],
F_[5][1][224],
F_[5][2][224],
F_[6][0][224],
F_[6][1][224],
F_[6][2][224],
F_[7][0][224],
F_[7][1][224],
F_[7][2][224],
F_[8][0][224],
F_[8][1][224],
F_[8][2][224],
F_[9][0][224],
F_[9][1][224],
F_[9][2][224],
F_[10][0][224],
F_[10][1][224],
F_[10][2][224],
F_[11][0][224],
F_[11][1][224],
F_[11][2][224],
F_[12][0][224],
F_[12][1][224],
F_[12][2][224],
F_[13][0][224],
F_[13][1][224],
F_[13][2][224],
F_[14][0][224],
F_[14][1][224],
F_[14][2][224],
F_[15][0][224],
F_[15][1][224],
F_[15][2][224],
F_[0][0][225],
F_[0][1][225],
F_[0][2][225],
F_[1][0][225],
F_[1][1][225],
F_[1][2][225],
F_[2][0][225],
F_[2][1][225],
F_[2][2][225],
F_[3][0][225],
F_[3][1][225],
F_[3][2][225],
F_[4][0][225],
F_[4][1][225],
F_[4][2][225],
F_[5][0][225],
F_[5][1][225],
F_[5][2][225],
F_[6][0][225],
F_[6][1][225],
F_[6][2][225],
F_[7][0][225],
F_[7][1][225],
F_[7][2][225],
F_[8][0][225],
F_[8][1][225],
F_[8][2][225],
F_[9][0][225],
F_[9][1][225],
F_[9][2][225],
F_[10][0][225],
F_[10][1][225],
F_[10][2][225],
F_[11][0][225],
F_[11][1][225],
F_[11][2][225],
F_[12][0][225],
F_[12][1][225],
F_[12][2][225],
F_[13][0][225],
F_[13][1][225],
F_[13][2][225],
F_[14][0][225],
F_[14][1][225],
F_[14][2][225],
F_[15][0][225],
F_[15][1][225],
F_[15][2][225],
F_[0][0][226],
F_[0][1][226],
F_[0][2][226],
F_[1][0][226],
F_[1][1][226],
F_[1][2][226],
F_[2][0][226],
F_[2][1][226],
F_[2][2][226],
F_[3][0][226],
F_[3][1][226],
F_[3][2][226],
F_[4][0][226],
F_[4][1][226],
F_[4][2][226],
F_[5][0][226],
F_[5][1][226],
F_[5][2][226],
F_[6][0][226],
F_[6][1][226],
F_[6][2][226],
F_[7][0][226],
F_[7][1][226],
F_[7][2][226],
F_[8][0][226],
F_[8][1][226],
F_[8][2][226],
F_[9][0][226],
F_[9][1][226],
F_[9][2][226],
F_[10][0][226],
F_[10][1][226],
F_[10][2][226],
F_[11][0][226],
F_[11][1][226],
F_[11][2][226],
F_[12][0][226],
F_[12][1][226],
F_[12][2][226],
F_[13][0][226],
F_[13][1][226],
F_[13][2][226],
F_[14][0][226],
F_[14][1][226],
F_[14][2][226],
F_[15][0][226],
F_[15][1][226],
F_[15][2][226],
F_[0][0][227],
F_[0][1][227],
F_[0][2][227],
F_[1][0][227],
F_[1][1][227],
F_[1][2][227],
F_[2][0][227],
F_[2][1][227],
F_[2][2][227],
F_[3][0][227],
F_[3][1][227],
F_[3][2][227],
F_[4][0][227],
F_[4][1][227],
F_[4][2][227],
F_[5][0][227],
F_[5][1][227],
F_[5][2][227],
F_[6][0][227],
F_[6][1][227],
F_[6][2][227],
F_[7][0][227],
F_[7][1][227],
F_[7][2][227],
F_[8][0][227],
F_[8][1][227],
F_[8][2][227],
F_[9][0][227],
F_[9][1][227],
F_[9][2][227],
F_[10][0][227],
F_[10][1][227],
F_[10][2][227],
F_[11][0][227],
F_[11][1][227],
F_[11][2][227],
F_[12][0][227],
F_[12][1][227],
F_[12][2][227],
F_[13][0][227],
F_[13][1][227],
F_[13][2][227],
F_[14][0][227],
F_[14][1][227],
F_[14][2][227],
F_[15][0][227],
F_[15][1][227],
F_[15][2][227],
F_[0][0][228],
F_[0][1][228],
F_[0][2][228],
F_[1][0][228],
F_[1][1][228],
F_[1][2][228],
F_[2][0][228],
F_[2][1][228],
F_[2][2][228],
F_[3][0][228],
F_[3][1][228],
F_[3][2][228],
F_[4][0][228],
F_[4][1][228],
F_[4][2][228],
F_[5][0][228],
F_[5][1][228],
F_[5][2][228],
F_[6][0][228],
F_[6][1][228],
F_[6][2][228],
F_[7][0][228],
F_[7][1][228],
F_[7][2][228],
F_[8][0][228],
F_[8][1][228],
F_[8][2][228],
F_[9][0][228],
F_[9][1][228],
F_[9][2][228],
F_[10][0][228],
F_[10][1][228],
F_[10][2][228],
F_[11][0][228],
F_[11][1][228],
F_[11][2][228],
F_[12][0][228],
F_[12][1][228],
F_[12][2][228],
F_[13][0][228],
F_[13][1][228],
F_[13][2][228],
F_[14][0][228],
F_[14][1][228],
F_[14][2][228],
F_[15][0][228],
F_[15][1][228],
F_[15][2][228],
F_[0][0][229],
F_[0][1][229],
F_[0][2][229],
F_[1][0][229],
F_[1][1][229],
F_[1][2][229],
F_[2][0][229],
F_[2][1][229],
F_[2][2][229],
F_[3][0][229],
F_[3][1][229],
F_[3][2][229],
F_[4][0][229],
F_[4][1][229],
F_[4][2][229],
F_[5][0][229],
F_[5][1][229],
F_[5][2][229],
F_[6][0][229],
F_[6][1][229],
F_[6][2][229],
F_[7][0][229],
F_[7][1][229],
F_[7][2][229],
F_[8][0][229],
F_[8][1][229],
F_[8][2][229],
F_[9][0][229],
F_[9][1][229],
F_[9][2][229],
F_[10][0][229],
F_[10][1][229],
F_[10][2][229],
F_[11][0][229],
F_[11][1][229],
F_[11][2][229],
F_[12][0][229],
F_[12][1][229],
F_[12][2][229],
F_[13][0][229],
F_[13][1][229],
F_[13][2][229],
F_[14][0][229],
F_[14][1][229],
F_[14][2][229],
F_[15][0][229],
F_[15][1][229],
F_[15][2][229],
F_[0][0][230],
F_[0][1][230],
F_[0][2][230],
F_[1][0][230],
F_[1][1][230],
F_[1][2][230],
F_[2][0][230],
F_[2][1][230],
F_[2][2][230],
F_[3][0][230],
F_[3][1][230],
F_[3][2][230],
F_[4][0][230],
F_[4][1][230],
F_[4][2][230],
F_[5][0][230],
F_[5][1][230],
F_[5][2][230],
F_[6][0][230],
F_[6][1][230],
F_[6][2][230],
F_[7][0][230],
F_[7][1][230],
F_[7][2][230],
F_[8][0][230],
F_[8][1][230],
F_[8][2][230],
F_[9][0][230],
F_[9][1][230],
F_[9][2][230],
F_[10][0][230],
F_[10][1][230],
F_[10][2][230],
F_[11][0][230],
F_[11][1][230],
F_[11][2][230],
F_[12][0][230],
F_[12][1][230],
F_[12][2][230],
F_[13][0][230],
F_[13][1][230],
F_[13][2][230],
F_[14][0][230],
F_[14][1][230],
F_[14][2][230],
F_[15][0][230],
F_[15][1][230],
F_[15][2][230],
F_[0][0][231],
F_[0][1][231],
F_[0][2][231],
F_[1][0][231],
F_[1][1][231],
F_[1][2][231],
F_[2][0][231],
F_[2][1][231],
F_[2][2][231],
F_[3][0][231],
F_[3][1][231],
F_[3][2][231],
F_[4][0][231],
F_[4][1][231],
F_[4][2][231],
F_[5][0][231],
F_[5][1][231],
F_[5][2][231],
F_[6][0][231],
F_[6][1][231],
F_[6][2][231],
F_[7][0][231],
F_[7][1][231],
F_[7][2][231],
F_[8][0][231],
F_[8][1][231],
F_[8][2][231],
F_[9][0][231],
F_[9][1][231],
F_[9][2][231],
F_[10][0][231],
F_[10][1][231],
F_[10][2][231],
F_[11][0][231],
F_[11][1][231],
F_[11][2][231],
F_[12][0][231],
F_[12][1][231],
F_[12][2][231],
F_[13][0][231],
F_[13][1][231],
F_[13][2][231],
F_[14][0][231],
F_[14][1][231],
F_[14][2][231],
F_[15][0][231],
F_[15][1][231],
F_[15][2][231],
F_[0][0][232],
F_[0][1][232],
F_[0][2][232],
F_[1][0][232],
F_[1][1][232],
F_[1][2][232],
F_[2][0][232],
F_[2][1][232],
F_[2][2][232],
F_[3][0][232],
F_[3][1][232],
F_[3][2][232],
F_[4][0][232],
F_[4][1][232],
F_[4][2][232],
F_[5][0][232],
F_[5][1][232],
F_[5][2][232],
F_[6][0][232],
F_[6][1][232],
F_[6][2][232],
F_[7][0][232],
F_[7][1][232],
F_[7][2][232],
F_[8][0][232],
F_[8][1][232],
F_[8][2][232],
F_[9][0][232],
F_[9][1][232],
F_[9][2][232],
F_[10][0][232],
F_[10][1][232],
F_[10][2][232],
F_[11][0][232],
F_[11][1][232],
F_[11][2][232],
F_[12][0][232],
F_[12][1][232],
F_[12][2][232],
F_[13][0][232],
F_[13][1][232],
F_[13][2][232],
F_[14][0][232],
F_[14][1][232],
F_[14][2][232],
F_[15][0][232],
F_[15][1][232],
F_[15][2][232],
F_[0][0][233],
F_[0][1][233],
F_[0][2][233],
F_[1][0][233],
F_[1][1][233],
F_[1][2][233],
F_[2][0][233],
F_[2][1][233],
F_[2][2][233],
F_[3][0][233],
F_[3][1][233],
F_[3][2][233],
F_[4][0][233],
F_[4][1][233],
F_[4][2][233],
F_[5][0][233],
F_[5][1][233],
F_[5][2][233],
F_[6][0][233],
F_[6][1][233],
F_[6][2][233],
F_[7][0][233],
F_[7][1][233],
F_[7][2][233],
F_[8][0][233],
F_[8][1][233],
F_[8][2][233],
F_[9][0][233],
F_[9][1][233],
F_[9][2][233],
F_[10][0][233],
F_[10][1][233],
F_[10][2][233],
F_[11][0][233],
F_[11][1][233],
F_[11][2][233],
F_[12][0][233],
F_[12][1][233],
F_[12][2][233],
F_[13][0][233],
F_[13][1][233],
F_[13][2][233],
F_[14][0][233],
F_[14][1][233],
F_[14][2][233],
F_[15][0][233],
F_[15][1][233],
F_[15][2][233],
F_[0][0][234],
F_[0][1][234],
F_[0][2][234],
F_[1][0][234],
F_[1][1][234],
F_[1][2][234],
F_[2][0][234],
F_[2][1][234],
F_[2][2][234],
F_[3][0][234],
F_[3][1][234],
F_[3][2][234],
F_[4][0][234],
F_[4][1][234],
F_[4][2][234],
F_[5][0][234],
F_[5][1][234],
F_[5][2][234],
F_[6][0][234],
F_[6][1][234],
F_[6][2][234],
F_[7][0][234],
F_[7][1][234],
F_[7][2][234],
F_[8][0][234],
F_[8][1][234],
F_[8][2][234],
F_[9][0][234],
F_[9][1][234],
F_[9][2][234],
F_[10][0][234],
F_[10][1][234],
F_[10][2][234],
F_[11][0][234],
F_[11][1][234],
F_[11][2][234],
F_[12][0][234],
F_[12][1][234],
F_[12][2][234],
F_[13][0][234],
F_[13][1][234],
F_[13][2][234],
F_[14][0][234],
F_[14][1][234],
F_[14][2][234],
F_[15][0][234],
F_[15][1][234],
F_[15][2][234],
F_[0][0][235],
F_[0][1][235],
F_[0][2][235],
F_[1][0][235],
F_[1][1][235],
F_[1][2][235],
F_[2][0][235],
F_[2][1][235],
F_[2][2][235],
F_[3][0][235],
F_[3][1][235],
F_[3][2][235],
F_[4][0][235],
F_[4][1][235],
F_[4][2][235],
F_[5][0][235],
F_[5][1][235],
F_[5][2][235],
F_[6][0][235],
F_[6][1][235],
F_[6][2][235],
F_[7][0][235],
F_[7][1][235],
F_[7][2][235],
F_[8][0][235],
F_[8][1][235],
F_[8][2][235],
F_[9][0][235],
F_[9][1][235],
F_[9][2][235],
F_[10][0][235],
F_[10][1][235],
F_[10][2][235],
F_[11][0][235],
F_[11][1][235],
F_[11][2][235],
F_[12][0][235],
F_[12][1][235],
F_[12][2][235],
F_[13][0][235],
F_[13][1][235],
F_[13][2][235],
F_[14][0][235],
F_[14][1][235],
F_[14][2][235],
F_[15][0][235],
F_[15][1][235],
F_[15][2][235],
F_[0][0][236],
F_[0][1][236],
F_[0][2][236],
F_[1][0][236],
F_[1][1][236],
F_[1][2][236],
F_[2][0][236],
F_[2][1][236],
F_[2][2][236],
F_[3][0][236],
F_[3][1][236],
F_[3][2][236],
F_[4][0][236],
F_[4][1][236],
F_[4][2][236],
F_[5][0][236],
F_[5][1][236],
F_[5][2][236],
F_[6][0][236],
F_[6][1][236],
F_[6][2][236],
F_[7][0][236],
F_[7][1][236],
F_[7][2][236],
F_[8][0][236],
F_[8][1][236],
F_[8][2][236],
F_[9][0][236],
F_[9][1][236],
F_[9][2][236],
F_[10][0][236],
F_[10][1][236],
F_[10][2][236],
F_[11][0][236],
F_[11][1][236],
F_[11][2][236],
F_[12][0][236],
F_[12][1][236],
F_[12][2][236],
F_[13][0][236],
F_[13][1][236],
F_[13][2][236],
F_[14][0][236],
F_[14][1][236],
F_[14][2][236],
F_[15][0][236],
F_[15][1][236],
F_[15][2][236],
F_[0][0][237],
F_[0][1][237],
F_[0][2][237],
F_[1][0][237],
F_[1][1][237],
F_[1][2][237],
F_[2][0][237],
F_[2][1][237],
F_[2][2][237],
F_[3][0][237],
F_[3][1][237],
F_[3][2][237],
F_[4][0][237],
F_[4][1][237],
F_[4][2][237],
F_[5][0][237],
F_[5][1][237],
F_[5][2][237],
F_[6][0][237],
F_[6][1][237],
F_[6][2][237],
F_[7][0][237],
F_[7][1][237],
F_[7][2][237],
F_[8][0][237],
F_[8][1][237],
F_[8][2][237],
F_[9][0][237],
F_[9][1][237],
F_[9][2][237],
F_[10][0][237],
F_[10][1][237],
F_[10][2][237],
F_[11][0][237],
F_[11][1][237],
F_[11][2][237],
F_[12][0][237],
F_[12][1][237],
F_[12][2][237],
F_[13][0][237],
F_[13][1][237],
F_[13][2][237],
F_[14][0][237],
F_[14][1][237],
F_[14][2][237],
F_[15][0][237],
F_[15][1][237],
F_[15][2][237],
F_[0][0][238],
F_[0][1][238],
F_[0][2][238],
F_[1][0][238],
F_[1][1][238],
F_[1][2][238],
F_[2][0][238],
F_[2][1][238],
F_[2][2][238],
F_[3][0][238],
F_[3][1][238],
F_[3][2][238],
F_[4][0][238],
F_[4][1][238],
F_[4][2][238],
F_[5][0][238],
F_[5][1][238],
F_[5][2][238],
F_[6][0][238],
F_[6][1][238],
F_[6][2][238],
F_[7][0][238],
F_[7][1][238],
F_[7][2][238],
F_[8][0][238],
F_[8][1][238],
F_[8][2][238],
F_[9][0][238],
F_[9][1][238],
F_[9][2][238],
F_[10][0][238],
F_[10][1][238],
F_[10][2][238],
F_[11][0][238],
F_[11][1][238],
F_[11][2][238],
F_[12][0][238],
F_[12][1][238],
F_[12][2][238],
F_[13][0][238],
F_[13][1][238],
F_[13][2][238],
F_[14][0][238],
F_[14][1][238],
F_[14][2][238],
F_[15][0][238],
F_[15][1][238],
F_[15][2][238],
F_[0][0][239],
F_[0][1][239],
F_[0][2][239],
F_[1][0][239],
F_[1][1][239],
F_[1][2][239],
F_[2][0][239],
F_[2][1][239],
F_[2][2][239],
F_[3][0][239],
F_[3][1][239],
F_[3][2][239],
F_[4][0][239],
F_[4][1][239],
F_[4][2][239],
F_[5][0][239],
F_[5][1][239],
F_[5][2][239],
F_[6][0][239],
F_[6][1][239],
F_[6][2][239],
F_[7][0][239],
F_[7][1][239],
F_[7][2][239],
F_[8][0][239],
F_[8][1][239],
F_[8][2][239],
F_[9][0][239],
F_[9][1][239],
F_[9][2][239],
F_[10][0][239],
F_[10][1][239],
F_[10][2][239],
F_[11][0][239],
F_[11][1][239],
F_[11][2][239],
F_[12][0][239],
F_[12][1][239],
F_[12][2][239],
F_[13][0][239],
F_[13][1][239],
F_[13][2][239],
F_[14][0][239],
F_[14][1][239],
F_[14][2][239],
F_[15][0][239],
F_[15][1][239],
F_[15][2][239],
F_[0][0][240],
F_[0][1][240],
F_[0][2][240],
F_[1][0][240],
F_[1][1][240],
F_[1][2][240],
F_[2][0][240],
F_[2][1][240],
F_[2][2][240],
F_[3][0][240],
F_[3][1][240],
F_[3][2][240],
F_[4][0][240],
F_[4][1][240],
F_[4][2][240],
F_[5][0][240],
F_[5][1][240],
F_[5][2][240],
F_[6][0][240],
F_[6][1][240],
F_[6][2][240],
F_[7][0][240],
F_[7][1][240],
F_[7][2][240],
F_[8][0][240],
F_[8][1][240],
F_[8][2][240],
F_[9][0][240],
F_[9][1][240],
F_[9][2][240],
F_[10][0][240],
F_[10][1][240],
F_[10][2][240],
F_[11][0][240],
F_[11][1][240],
F_[11][2][240],
F_[12][0][240],
F_[12][1][240],
F_[12][2][240],
F_[13][0][240],
F_[13][1][240],
F_[13][2][240],
F_[14][0][240],
F_[14][1][240],
F_[14][2][240],
F_[15][0][240],
F_[15][1][240],
F_[15][2][240],
F_[0][0][241],
F_[0][1][241],
F_[0][2][241],
F_[1][0][241],
F_[1][1][241],
F_[1][2][241],
F_[2][0][241],
F_[2][1][241],
F_[2][2][241],
F_[3][0][241],
F_[3][1][241],
F_[3][2][241],
F_[4][0][241],
F_[4][1][241],
F_[4][2][241],
F_[5][0][241],
F_[5][1][241],
F_[5][2][241],
F_[6][0][241],
F_[6][1][241],
F_[6][2][241],
F_[7][0][241],
F_[7][1][241],
F_[7][2][241],
F_[8][0][241],
F_[8][1][241],
F_[8][2][241],
F_[9][0][241],
F_[9][1][241],
F_[9][2][241],
F_[10][0][241],
F_[10][1][241],
F_[10][2][241],
F_[11][0][241],
F_[11][1][241],
F_[11][2][241],
F_[12][0][241],
F_[12][1][241],
F_[12][2][241],
F_[13][0][241],
F_[13][1][241],
F_[13][2][241],
F_[14][0][241],
F_[14][1][241],
F_[14][2][241],
F_[15][0][241],
F_[15][1][241],
F_[15][2][241],
F_[0][0][242],
F_[0][1][242],
F_[0][2][242],
F_[1][0][242],
F_[1][1][242],
F_[1][2][242],
F_[2][0][242],
F_[2][1][242],
F_[2][2][242],
F_[3][0][242],
F_[3][1][242],
F_[3][2][242],
F_[4][0][242],
F_[4][1][242],
F_[4][2][242],
F_[5][0][242],
F_[5][1][242],
F_[5][2][242],
F_[6][0][242],
F_[6][1][242],
F_[6][2][242],
F_[7][0][242],
F_[7][1][242],
F_[7][2][242],
F_[8][0][242],
F_[8][1][242],
F_[8][2][242],
F_[9][0][242],
F_[9][1][242],
F_[9][2][242],
F_[10][0][242],
F_[10][1][242],
F_[10][2][242],
F_[11][0][242],
F_[11][1][242],
F_[11][2][242],
F_[12][0][242],
F_[12][1][242],
F_[12][2][242],
F_[13][0][242],
F_[13][1][242],
F_[13][2][242],
F_[14][0][242],
F_[14][1][242],
F_[14][2][242],
F_[15][0][242],
F_[15][1][242],
F_[15][2][242],
F_[0][0][243],
F_[0][1][243],
F_[0][2][243],
F_[1][0][243],
F_[1][1][243],
F_[1][2][243],
F_[2][0][243],
F_[2][1][243],
F_[2][2][243],
F_[3][0][243],
F_[3][1][243],
F_[3][2][243],
F_[4][0][243],
F_[4][1][243],
F_[4][2][243],
F_[5][0][243],
F_[5][1][243],
F_[5][2][243],
F_[6][0][243],
F_[6][1][243],
F_[6][2][243],
F_[7][0][243],
F_[7][1][243],
F_[7][2][243],
F_[8][0][243],
F_[8][1][243],
F_[8][2][243],
F_[9][0][243],
F_[9][1][243],
F_[9][2][243],
F_[10][0][243],
F_[10][1][243],
F_[10][2][243],
F_[11][0][243],
F_[11][1][243],
F_[11][2][243],
F_[12][0][243],
F_[12][1][243],
F_[12][2][243],
F_[13][0][243],
F_[13][1][243],
F_[13][2][243],
F_[14][0][243],
F_[14][1][243],
F_[14][2][243],
F_[15][0][243],
F_[15][1][243],
F_[15][2][243],
F_[0][0][244],
F_[0][1][244],
F_[0][2][244],
F_[1][0][244],
F_[1][1][244],
F_[1][2][244],
F_[2][0][244],
F_[2][1][244],
F_[2][2][244],
F_[3][0][244],
F_[3][1][244],
F_[3][2][244],
F_[4][0][244],
F_[4][1][244],
F_[4][2][244],
F_[5][0][244],
F_[5][1][244],
F_[5][2][244],
F_[6][0][244],
F_[6][1][244],
F_[6][2][244],
F_[7][0][244],
F_[7][1][244],
F_[7][2][244],
F_[8][0][244],
F_[8][1][244],
F_[8][2][244],
F_[9][0][244],
F_[9][1][244],
F_[9][2][244],
F_[10][0][244],
F_[10][1][244],
F_[10][2][244],
F_[11][0][244],
F_[11][1][244],
F_[11][2][244],
F_[12][0][244],
F_[12][1][244],
F_[12][2][244],
F_[13][0][244],
F_[13][1][244],
F_[13][2][244],
F_[14][0][244],
F_[14][1][244],
F_[14][2][244],
F_[15][0][244],
F_[15][1][244],
F_[15][2][244],
F_[0][0][245],
F_[0][1][245],
F_[0][2][245],
F_[1][0][245],
F_[1][1][245],
F_[1][2][245],
F_[2][0][245],
F_[2][1][245],
F_[2][2][245],
F_[3][0][245],
F_[3][1][245],
F_[3][2][245],
F_[4][0][245],
F_[4][1][245],
F_[4][2][245],
F_[5][0][245],
F_[5][1][245],
F_[5][2][245],
F_[6][0][245],
F_[6][1][245],
F_[6][2][245],
F_[7][0][245],
F_[7][1][245],
F_[7][2][245],
F_[8][0][245],
F_[8][1][245],
F_[8][2][245],
F_[9][0][245],
F_[9][1][245],
F_[9][2][245],
F_[10][0][245],
F_[10][1][245],
F_[10][2][245],
F_[11][0][245],
F_[11][1][245],
F_[11][2][245],
F_[12][0][245],
F_[12][1][245],
F_[12][2][245],
F_[13][0][245],
F_[13][1][245],
F_[13][2][245],
F_[14][0][245],
F_[14][1][245],
F_[14][2][245],
F_[15][0][245],
F_[15][1][245],
F_[15][2][245],
F_[0][0][246],
F_[0][1][246],
F_[0][2][246],
F_[1][0][246],
F_[1][1][246],
F_[1][2][246],
F_[2][0][246],
F_[2][1][246],
F_[2][2][246],
F_[3][0][246],
F_[3][1][246],
F_[3][2][246],
F_[4][0][246],
F_[4][1][246],
F_[4][2][246],
F_[5][0][246],
F_[5][1][246],
F_[5][2][246],
F_[6][0][246],
F_[6][1][246],
F_[6][2][246],
F_[7][0][246],
F_[7][1][246],
F_[7][2][246],
F_[8][0][246],
F_[8][1][246],
F_[8][2][246],
F_[9][0][246],
F_[9][1][246],
F_[9][2][246],
F_[10][0][246],
F_[10][1][246],
F_[10][2][246],
F_[11][0][246],
F_[11][1][246],
F_[11][2][246],
F_[12][0][246],
F_[12][1][246],
F_[12][2][246],
F_[13][0][246],
F_[13][1][246],
F_[13][2][246],
F_[14][0][246],
F_[14][1][246],
F_[14][2][246],
F_[15][0][246],
F_[15][1][246],
F_[15][2][246],
F_[0][0][247],
F_[0][1][247],
F_[0][2][247],
F_[1][0][247],
F_[1][1][247],
F_[1][2][247],
F_[2][0][247],
F_[2][1][247],
F_[2][2][247],
F_[3][0][247],
F_[3][1][247],
F_[3][2][247],
F_[4][0][247],
F_[4][1][247],
F_[4][2][247],
F_[5][0][247],
F_[5][1][247],
F_[5][2][247],
F_[6][0][247],
F_[6][1][247],
F_[6][2][247],
F_[7][0][247],
F_[7][1][247],
F_[7][2][247],
F_[8][0][247],
F_[8][1][247],
F_[8][2][247],
F_[9][0][247],
F_[9][1][247],
F_[9][2][247],
F_[10][0][247],
F_[10][1][247],
F_[10][2][247],
F_[11][0][247],
F_[11][1][247],
F_[11][2][247],
F_[12][0][247],
F_[12][1][247],
F_[12][2][247],
F_[13][0][247],
F_[13][1][247],
F_[13][2][247],
F_[14][0][247],
F_[14][1][247],
F_[14][2][247],
F_[15][0][247],
F_[15][1][247],
F_[15][2][247],
F_[0][0][248],
F_[0][1][248],
F_[0][2][248],
F_[1][0][248],
F_[1][1][248],
F_[1][2][248],
F_[2][0][248],
F_[2][1][248],
F_[2][2][248],
F_[3][0][248],
F_[3][1][248],
F_[3][2][248],
F_[4][0][248],
F_[4][1][248],
F_[4][2][248],
F_[5][0][248],
F_[5][1][248],
F_[5][2][248],
F_[6][0][248],
F_[6][1][248],
F_[6][2][248],
F_[7][0][248],
F_[7][1][248],
F_[7][2][248],
F_[8][0][248],
F_[8][1][248],
F_[8][2][248],
F_[9][0][248],
F_[9][1][248],
F_[9][2][248],
F_[10][0][248],
F_[10][1][248],
F_[10][2][248],
F_[11][0][248],
F_[11][1][248],
F_[11][2][248],
F_[12][0][248],
F_[12][1][248],
F_[12][2][248],
F_[13][0][248],
F_[13][1][248],
F_[13][2][248],
F_[14][0][248],
F_[14][1][248],
F_[14][2][248],
F_[15][0][248],
F_[15][1][248],
F_[15][2][248],
F_[0][0][249],
F_[0][1][249],
F_[0][2][249],
F_[1][0][249],
F_[1][1][249],
F_[1][2][249],
F_[2][0][249],
F_[2][1][249],
F_[2][2][249],
F_[3][0][249],
F_[3][1][249],
F_[3][2][249],
F_[4][0][249],
F_[4][1][249],
F_[4][2][249],
F_[5][0][249],
F_[5][1][249],
F_[5][2][249],
F_[6][0][249],
F_[6][1][249],
F_[6][2][249],
F_[7][0][249],
F_[7][1][249],
F_[7][2][249],
F_[8][0][249],
F_[8][1][249],
F_[8][2][249],
F_[9][0][249],
F_[9][1][249],
F_[9][2][249],
F_[10][0][249],
F_[10][1][249],
F_[10][2][249],
F_[11][0][249],
F_[11][1][249],
F_[11][2][249],
F_[12][0][249],
F_[12][1][249],
F_[12][2][249],
F_[13][0][249],
F_[13][1][249],
F_[13][2][249],
F_[14][0][249],
F_[14][1][249],
F_[14][2][249],
F_[15][0][249],
F_[15][1][249],
F_[15][2][249],
F_[0][0][250],
F_[0][1][250],
F_[0][2][250],
F_[1][0][250],
F_[1][1][250],
F_[1][2][250],
F_[2][0][250],
F_[2][1][250],
F_[2][2][250],
F_[3][0][250],
F_[3][1][250],
F_[3][2][250],
F_[4][0][250],
F_[4][1][250],
F_[4][2][250],
F_[5][0][250],
F_[5][1][250],
F_[5][2][250],
F_[6][0][250],
F_[6][1][250],
F_[6][2][250],
F_[7][0][250],
F_[7][1][250],
F_[7][2][250],
F_[8][0][250],
F_[8][1][250],
F_[8][2][250],
F_[9][0][250],
F_[9][1][250],
F_[9][2][250],
F_[10][0][250],
F_[10][1][250],
F_[10][2][250],
F_[11][0][250],
F_[11][1][250],
F_[11][2][250],
F_[12][0][250],
F_[12][1][250],
F_[12][2][250],
F_[13][0][250],
F_[13][1][250],
F_[13][2][250],
F_[14][0][250],
F_[14][1][250],
F_[14][2][250],
F_[15][0][250],
F_[15][1][250],
F_[15][2][250],
F_[0][0][251],
F_[0][1][251],
F_[0][2][251],
F_[1][0][251],
F_[1][1][251],
F_[1][2][251],
F_[2][0][251],
F_[2][1][251],
F_[2][2][251],
F_[3][0][251],
F_[3][1][251],
F_[3][2][251],
F_[4][0][251],
F_[4][1][251],
F_[4][2][251],
F_[5][0][251],
F_[5][1][251],
F_[5][2][251],
F_[6][0][251],
F_[6][1][251],
F_[6][2][251],
F_[7][0][251],
F_[7][1][251],
F_[7][2][251],
F_[8][0][251],
F_[8][1][251],
F_[8][2][251],
F_[9][0][251],
F_[9][1][251],
F_[9][2][251],
F_[10][0][251],
F_[10][1][251],
F_[10][2][251],
F_[11][0][251],
F_[11][1][251],
F_[11][2][251],
F_[12][0][251],
F_[12][1][251],
F_[12][2][251],
F_[13][0][251],
F_[13][1][251],
F_[13][2][251],
F_[14][0][251],
F_[14][1][251],
F_[14][2][251],
F_[15][0][251],
F_[15][1][251],
F_[15][2][251],
F_[0][0][252],
F_[0][1][252],
F_[0][2][252],
F_[1][0][252],
F_[1][1][252],
F_[1][2][252],
F_[2][0][252],
F_[2][1][252],
F_[2][2][252],
F_[3][0][252],
F_[3][1][252],
F_[3][2][252],
F_[4][0][252],
F_[4][1][252],
F_[4][2][252],
F_[5][0][252],
F_[5][1][252],
F_[5][2][252],
F_[6][0][252],
F_[6][1][252],
F_[6][2][252],
F_[7][0][252],
F_[7][1][252],
F_[7][2][252],
F_[8][0][252],
F_[8][1][252],
F_[8][2][252],
F_[9][0][252],
F_[9][1][252],
F_[9][2][252],
F_[10][0][252],
F_[10][1][252],
F_[10][2][252],
F_[11][0][252],
F_[11][1][252],
F_[11][2][252],
F_[12][0][252],
F_[12][1][252],
F_[12][2][252],
F_[13][0][252],
F_[13][1][252],
F_[13][2][252],
F_[14][0][252],
F_[14][1][252],
F_[14][2][252],
F_[15][0][252],
F_[15][1][252],
F_[15][2][252],
F_[0][0][253],
F_[0][1][253],
F_[0][2][253],
F_[1][0][253],
F_[1][1][253],
F_[1][2][253],
F_[2][0][253],
F_[2][1][253],
F_[2][2][253],
F_[3][0][253],
F_[3][1][253],
F_[3][2][253],
F_[4][0][253],
F_[4][1][253],
F_[4][2][253],
F_[5][0][253],
F_[5][1][253],
F_[5][2][253],
F_[6][0][253],
F_[6][1][253],
F_[6][2][253],
F_[7][0][253],
F_[7][1][253],
F_[7][2][253],
F_[8][0][253],
F_[8][1][253],
F_[8][2][253],
F_[9][0][253],
F_[9][1][253],
F_[9][2][253],
F_[10][0][253],
F_[10][1][253],
F_[10][2][253],
F_[11][0][253],
F_[11][1][253],
F_[11][2][253],
F_[12][0][253],
F_[12][1][253],
F_[12][2][253],
F_[13][0][253],
F_[13][1][253],
F_[13][2][253],
F_[14][0][253],
F_[14][1][253],
F_[14][2][253],
F_[15][0][253],
F_[15][1][253],
F_[15][2][253],
F_[0][0][254],
F_[0][1][254],
F_[0][2][254],
F_[1][0][254],
F_[1][1][254],
F_[1][2][254],
F_[2][0][254],
F_[2][1][254],
F_[2][2][254],
F_[3][0][254],
F_[3][1][254],
F_[3][2][254],
F_[4][0][254],
F_[4][1][254],
F_[4][2][254],
F_[5][0][254],
F_[5][1][254],
F_[5][2][254],
F_[6][0][254],
F_[6][1][254],
F_[6][2][254],
F_[7][0][254],
F_[7][1][254],
F_[7][2][254],
F_[8][0][254],
F_[8][1][254],
F_[8][2][254],
F_[9][0][254],
F_[9][1][254],
F_[9][2][254],
F_[10][0][254],
F_[10][1][254],
F_[10][2][254],
F_[11][0][254],
F_[11][1][254],
F_[11][2][254],
F_[12][0][254],
F_[12][1][254],
F_[12][2][254],
F_[13][0][254],
F_[13][1][254],
F_[13][2][254],
F_[14][0][254],
F_[14][1][254],
F_[14][2][254],
F_[15][0][254],
F_[15][1][254],
F_[15][2][254],
F_[0][0][255],
F_[0][1][255],
F_[0][2][255],
F_[1][0][255],
F_[1][1][255],
F_[1][2][255],
F_[2][0][255],
F_[2][1][255],
F_[2][2][255],
F_[3][0][255],
F_[3][1][255],
F_[3][2][255],
F_[4][0][255],
F_[4][1][255],
F_[4][2][255],
F_[5][0][255],
F_[5][1][255],
F_[5][2][255],
F_[6][0][255],
F_[6][1][255],
F_[6][2][255],
F_[7][0][255],
F_[7][1][255],
F_[7][2][255],
F_[8][0][255],
F_[8][1][255],
F_[8][2][255],
F_[9][0][255],
F_[9][1][255],
F_[9][2][255],
F_[10][0][255],
F_[10][1][255],
F_[10][2][255],
F_[11][0][255],
F_[11][1][255],
F_[11][2][255],
F_[12][0][255],
F_[12][1][255],
F_[12][2][255],
F_[13][0][255],
F_[13][1][255],
F_[13][2][255],
F_[14][0][255],
F_[14][1][255],
F_[14][2][255],
F_[15][0][255],
F_[15][1][255],
F_[15][2][255],

   col_row[ 0 ][0],
   col_row[ 0 ][1],
   col_row[ 0 ][2],
   col_row[ 1 ][0],
   col_row[ 1 ][1],
   col_row[ 1 ][2],
   col_row[ 2 ][0],
   col_row[ 2 ][1],
   col_row[ 2 ][2],
   col_row[ 3 ][0],
   col_row[ 3 ][1],
   col_row[ 3 ][2],
   col_row[ 4 ][0],
   col_row[ 4 ][1],
   col_row[ 4 ][2],
   col_row[ 5 ][0],
   col_row[ 5 ][1],
   col_row[ 5 ][2],
   col_row[ 6 ][0],
   col_row[ 6 ][1],
   col_row[ 6 ][2],
   col_row[ 7 ][0],
   col_row[ 7 ][1],
   col_row[ 7 ][2],
   col_row[ 8 ][0],
   col_row[ 8 ][1],
   col_row[ 8 ][2],
   col_row[ 9 ][0],
   col_row[ 9 ][1],
   col_row[ 9 ][2],
   col_row[ 10 ][0],
   col_row[ 10 ][1],
   col_row[ 10 ][2],
   col_row[ 11 ][0],
   col_row[ 11 ][1],
   col_row[ 11 ][2],
   col_row[ 12 ][0],
   col_row[ 12 ][1],
   col_row[ 12 ][2],
   col_row[ 13 ][0],
   col_row[ 13 ][1],
   col_row[ 13 ][2],
   col_row[ 14 ][0],
   col_row[ 14 ][1],
   col_row[ 14 ][2],
   col_row[ 15 ][0],
   col_row[ 15 ][1],
   col_row[ 15 ][2],
   col_row[ 16 ][0],
   col_row[ 16 ][1],
   col_row[ 16 ][2],
   col_row[ 17 ][0],
   col_row[ 17 ][1],
   col_row[ 17 ][2],
   col_row[ 18 ][0],
   col_row[ 18 ][1],
   col_row[ 18 ][2],
   col_row[ 19 ][0],
   col_row[ 19 ][1],
   col_row[ 19 ][2],
   col_row[ 20 ][0],
   col_row[ 20 ][1],
   col_row[ 20 ][2],
   col_row[ 21 ][0],
   col_row[ 21 ][1],
   col_row[ 21 ][2],
   col_row[ 22 ][0],
   col_row[ 22 ][1],
   col_row[ 22 ][2],
   col_row[ 23 ][0],
   col_row[ 23 ][1],
   col_row[ 23 ][2],
   col_row[ 24 ][0],
   col_row[ 24 ][1],
   col_row[ 24 ][2],
   col_row[ 25 ][0],
   col_row[ 25 ][1],
   col_row[ 25 ][2],
   col_row[ 26 ][0],
   col_row[ 26 ][1],
   col_row[ 26 ][2],
   col_row[ 27 ][0],
   col_row[ 27 ][1],
   col_row[ 27 ][2],
   col_row[ 28 ][0],
   col_row[ 28 ][1],
   col_row[ 28 ][2],
   col_row[ 29 ][0],
   col_row[ 29 ][1],
   col_row[ 29 ][2],
   col_row[ 30 ][0],
   col_row[ 30 ][1],
   col_row[ 30 ][2],
   col_row[ 31 ][0],
   col_row[ 31 ][1],
   col_row[ 31 ][2],
   col_row[ 32 ][0],
   col_row[ 32 ][1],
   col_row[ 32 ][2],
   col_row[ 33 ][0],
   col_row[ 33 ][1],
   col_row[ 33 ][2],
   col_row[ 34 ][0],
   col_row[ 34 ][1],
   col_row[ 34 ][2],
   col_row[ 35 ][0],
   col_row[ 35 ][1],
   col_row[ 35 ][2],
   col_row[ 36 ][0],
   col_row[ 36 ][1],
   col_row[ 36 ][2],
   col_row[ 37 ][0],
   col_row[ 37 ][1],
   col_row[ 37 ][2],
   col_row[ 38 ][0],
   col_row[ 38 ][1],
   col_row[ 38 ][2],
   col_row[ 39 ][0],
   col_row[ 39 ][1],
   col_row[ 39 ][2],
   col_row[ 40 ][0],
   col_row[ 40 ][1],
   col_row[ 40 ][2],
   col_row[ 41 ][0],
   col_row[ 41 ][1],
   col_row[ 41 ][2],
   col_row[ 42 ][0],
   col_row[ 42 ][1],
   col_row[ 42 ][2],
   col_row[ 43 ][0],
   col_row[ 43 ][1],
   col_row[ 43 ][2],
   col_row[ 44 ][0],
   col_row[ 44 ][1],
   col_row[ 44 ][2],
   col_row[ 45 ][0],
   col_row[ 45 ][1],
   col_row[ 45 ][2],
   col_row[ 46 ][0],
   col_row[ 46 ][1],
   col_row[ 46 ][2],
   col_row[ 47 ][0],
   col_row[ 47 ][1],
   col_row[ 47 ][2],
   col_row[ 48 ][0],
   col_row[ 48 ][1],
   col_row[ 48 ][2],
   col_row[ 49 ][0],
   col_row[ 49 ][1],
   col_row[ 49 ][2],
   col_row[ 50 ][0],
   col_row[ 50 ][1],
   col_row[ 50 ][2],
   col_row[ 51 ][0],
   col_row[ 51 ][1],
   col_row[ 51 ][2],
   col_row[ 52 ][0],
   col_row[ 52 ][1],
   col_row[ 52 ][2],
   col_row[ 53 ][0],
   col_row[ 53 ][1],
   col_row[ 53 ][2],
   col_row[ 54 ][0],
   col_row[ 54 ][1],
   col_row[ 54 ][2],
   col_row[ 55 ][0],
   col_row[ 55 ][1],
   col_row[ 55 ][2],
   col_row[ 56 ][0],
   col_row[ 56 ][1],
   col_row[ 56 ][2],
   col_row[ 57 ][0],
   col_row[ 57 ][1],
   col_row[ 57 ][2],
   col_row[ 58 ][0],
   col_row[ 58 ][1],
   col_row[ 58 ][2],
   col_row[ 59 ][0],
   col_row[ 59 ][1],
   col_row[ 59 ][2],
   col_row[ 60 ][0],
   col_row[ 60 ][1],
   col_row[ 60 ][2],
   col_row[ 61 ][0],
   col_row[ 61 ][1],
   col_row[ 61 ][2],
   col_row[ 62 ][0],
   col_row[ 62 ][1],
   col_row[ 62 ][2],
   col_row[ 63 ][0],
   col_row[ 63 ][1],
   col_row[ 63 ][2],
   col_row[ 64 ][0],
   col_row[ 64 ][1],
   col_row[ 64 ][2],
   col_row[ 65 ][0],
   col_row[ 65 ][1],
   col_row[ 65 ][2],
   col_row[ 66 ][0],
   col_row[ 66 ][1],
   col_row[ 66 ][2],
   col_row[ 67 ][0],
   col_row[ 67 ][1],
   col_row[ 67 ][2],
   col_row[ 68 ][0],
   col_row[ 68 ][1],
   col_row[ 68 ][2],
   col_row[ 69 ][0],
   col_row[ 69 ][1],
   col_row[ 69 ][2],
   col_row[ 70 ][0],
   col_row[ 70 ][1],
   col_row[ 70 ][2],
   col_row[ 71 ][0],
   col_row[ 71 ][1],
   col_row[ 71 ][2],
   col_row[ 72 ][0],
   col_row[ 72 ][1],
   col_row[ 72 ][2],
   col_row[ 73 ][0],
   col_row[ 73 ][1],
   col_row[ 73 ][2],
   col_row[ 74 ][0],
   col_row[ 74 ][1],
   col_row[ 74 ][2],
   col_row[ 75 ][0],
   col_row[ 75 ][1],
   col_row[ 75 ][2],
   col_row[ 76 ][0],
   col_row[ 76 ][1],
   col_row[ 76 ][2],
   col_row[ 77 ][0],
   col_row[ 77 ][1],
   col_row[ 77 ][2],
   col_row[ 78 ][0],
   col_row[ 78 ][1],
   col_row[ 78 ][2],
   col_row[ 79 ][0],
   col_row[ 79 ][1],
   col_row[ 79 ][2],
   col_row[ 80 ][0],
   col_row[ 80 ][1],
   col_row[ 80 ][2],
   col_row[ 81 ][0],
   col_row[ 81 ][1],
   col_row[ 81 ][2],
   col_row[ 82 ][0],
   col_row[ 82 ][1],
   col_row[ 82 ][2],
   col_row[ 83 ][0],
   col_row[ 83 ][1],
   col_row[ 83 ][2],
   col_row[ 84 ][0],
   col_row[ 84 ][1],
   col_row[ 84 ][2],
   col_row[ 85 ][0],
   col_row[ 85 ][1],
   col_row[ 85 ][2],
   col_row[ 86 ][0],
   col_row[ 86 ][1],
   col_row[ 86 ][2],
   col_row[ 87 ][0],
   col_row[ 87 ][1],
   col_row[ 87 ][2],
   col_row[ 88 ][0],
   col_row[ 88 ][1],
   col_row[ 88 ][2],
   col_row[ 89 ][0],
   col_row[ 89 ][1],
   col_row[ 89 ][2],
   col_row[ 90 ][0],
   col_row[ 90 ][1],
   col_row[ 90 ][2],
   col_row[ 91 ][0],
   col_row[ 91 ][1],
   col_row[ 91 ][2],
   col_row[ 92 ][0],
   col_row[ 92 ][1],
   col_row[ 92 ][2],
   col_row[ 93 ][0],
   col_row[ 93 ][1],
   col_row[ 93 ][2],
   col_row[ 94 ][0],
   col_row[ 94 ][1],
   col_row[ 94 ][2],
   col_row[ 95 ][0],
   col_row[ 95 ][1],
   col_row[ 95 ][2],
   col_row[ 96 ][0],
   col_row[ 96 ][1],
   col_row[ 96 ][2],
   col_row[ 97 ][0],
   col_row[ 97 ][1],
   col_row[ 97 ][2],
   col_row[ 98 ][0],
   col_row[ 98 ][1],
   col_row[ 98 ][2],
   col_row[ 99 ][0],
   col_row[ 99 ][1],
   col_row[ 99 ][2],
   col_row[ 100 ][0],
   col_row[ 100 ][1],
   col_row[ 100 ][2],
   col_row[ 101 ][0],
   col_row[ 101 ][1],
   col_row[ 101 ][2],
   col_row[ 102 ][0],
   col_row[ 102 ][1],
   col_row[ 102 ][2],
   col_row[ 103 ][0],
   col_row[ 103 ][1],
   col_row[ 103 ][2],
   col_row[ 104 ][0],
   col_row[ 104 ][1],
   col_row[ 104 ][2],
   col_row[ 105 ][0],
   col_row[ 105 ][1],
   col_row[ 105 ][2],
   col_row[ 106 ][0],
   col_row[ 106 ][1],
   col_row[ 106 ][2],
   col_row[ 107 ][0],
   col_row[ 107 ][1],
   col_row[ 107 ][2],
   col_row[ 108 ][0],
   col_row[ 108 ][1],
   col_row[ 108 ][2],
   col_row[ 109 ][0],
   col_row[ 109 ][1],
   col_row[ 109 ][2],
   col_row[ 110 ][0],
   col_row[ 110 ][1],
   col_row[ 110 ][2],
   col_row[ 111 ][0],
   col_row[ 111 ][1],
   col_row[ 111 ][2],
   col_row[ 112 ][0],
   col_row[ 112 ][1],
   col_row[ 112 ][2],
   col_row[ 113 ][0],
   col_row[ 113 ][1],
   col_row[ 113 ][2],
   col_row[ 114 ][0],
   col_row[ 114 ][1],
   col_row[ 114 ][2],
   col_row[ 115 ][0],
   col_row[ 115 ][1],
   col_row[ 115 ][2],
   col_row[ 116 ][0],
   col_row[ 116 ][1],
   col_row[ 116 ][2],
   col_row[ 117 ][0],
   col_row[ 117 ][1],
   col_row[ 117 ][2],
   col_row[ 118 ][0],
   col_row[ 118 ][1],
   col_row[ 118 ][2],
   col_row[ 119 ][0],
   col_row[ 119 ][1],
   col_row[ 119 ][2],
   col_row[ 120 ][0],
   col_row[ 120 ][1],
   col_row[ 120 ][2],
   col_row[ 121 ][0],
   col_row[ 121 ][1],
   col_row[ 121 ][2],
   col_row[ 122 ][0],
   col_row[ 122 ][1],
   col_row[ 122 ][2],
   col_row[ 123 ][0],
   col_row[ 123 ][1],
   col_row[ 123 ][2],
   col_row[ 124 ][0],
   col_row[ 124 ][1],
   col_row[ 124 ][2],
   col_row[ 125 ][0],
   col_row[ 125 ][1],
   col_row[ 125 ][2],
   col_row[ 126 ][0],
   col_row[ 126 ][1],
   col_row[ 126 ][2],
   col_row[ 127 ][0],
   col_row[ 127 ][1],
   col_row[ 127 ][2],
   col_row[ 128 ][0],
   col_row[ 128 ][1],
   col_row[ 128 ][2],
   col_row[ 129 ][0],
   col_row[ 129 ][1],
   col_row[ 129 ][2],
   col_row[ 130 ][0],
   col_row[ 130 ][1],
   col_row[ 130 ][2],
   col_row[ 131 ][0],
   col_row[ 131 ][1],
   col_row[ 131 ][2],
   col_row[ 132 ][0],
   col_row[ 132 ][1],
   col_row[ 132 ][2],
   col_row[ 133 ][0],
   col_row[ 133 ][1],
   col_row[ 133 ][2],
   col_row[ 134 ][0],
   col_row[ 134 ][1],
   col_row[ 134 ][2],
   col_row[ 135 ][0],
   col_row[ 135 ][1],
   col_row[ 135 ][2],
   col_row[ 136 ][0],
   col_row[ 136 ][1],
   col_row[ 136 ][2],
   col_row[ 137 ][0],
   col_row[ 137 ][1],
   col_row[ 137 ][2],
   col_row[ 138 ][0],
   col_row[ 138 ][1],
   col_row[ 138 ][2],
   col_row[ 139 ][0],
   col_row[ 139 ][1],
   col_row[ 139 ][2],
   col_row[ 140 ][0],
   col_row[ 140 ][1],
   col_row[ 140 ][2],
   col_row[ 141 ][0],
   col_row[ 141 ][1],
   col_row[ 141 ][2],
   col_row[ 142 ][0],
   col_row[ 142 ][1],
   col_row[ 142 ][2],
   col_row[ 143 ][0],
   col_row[ 143 ][1],
   col_row[ 143 ][2],
   col_row[ 144 ][0],
   col_row[ 144 ][1],
   col_row[ 144 ][2],
   col_row[ 145 ][0],
   col_row[ 145 ][1],
   col_row[ 145 ][2],
   col_row[ 146 ][0],
   col_row[ 146 ][1],
   col_row[ 146 ][2],
   col_row[ 147 ][0],
   col_row[ 147 ][1],
   col_row[ 147 ][2],
   col_row[ 148 ][0],
   col_row[ 148 ][1],
   col_row[ 148 ][2],
   col_row[ 149 ][0],
   col_row[ 149 ][1],
   col_row[ 149 ][2],
   col_row[ 150 ][0],
   col_row[ 150 ][1],
   col_row[ 150 ][2],
   col_row[ 151 ][0],
   col_row[ 151 ][1],
   col_row[ 151 ][2],
   col_row[ 152 ][0],
   col_row[ 152 ][1],
   col_row[ 152 ][2],
   col_row[ 153 ][0],
   col_row[ 153 ][1],
   col_row[ 153 ][2],
   col_row[ 154 ][0],
   col_row[ 154 ][1],
   col_row[ 154 ][2],
   col_row[ 155 ][0],
   col_row[ 155 ][1],
   col_row[ 155 ][2],
   col_row[ 156 ][0],
   col_row[ 156 ][1],
   col_row[ 156 ][2],
   col_row[ 157 ][0],
   col_row[ 157 ][1],
   col_row[ 157 ][2],
   col_row[ 158 ][0],
   col_row[ 158 ][1],
   col_row[ 158 ][2],
   col_row[ 159 ][0],
   col_row[ 159 ][1],
   col_row[ 159 ][2],
   col_row[ 160 ][0],
   col_row[ 160 ][1],
   col_row[ 160 ][2],
   col_row[ 161 ][0],
   col_row[ 161 ][1],
   col_row[ 161 ][2],
   col_row[ 162 ][0],
   col_row[ 162 ][1],
   col_row[ 162 ][2],
   col_row[ 163 ][0],
   col_row[ 163 ][1],
   col_row[ 163 ][2],
   col_row[ 164 ][0],
   col_row[ 164 ][1],
   col_row[ 164 ][2],
   col_row[ 165 ][0],
   col_row[ 165 ][1],
   col_row[ 165 ][2],
   col_row[ 166 ][0],
   col_row[ 166 ][1],
   col_row[ 166 ][2],
   col_row[ 167 ][0],
   col_row[ 167 ][1],
   col_row[ 167 ][2],
   col_row[ 168 ][0],
   col_row[ 168 ][1],
   col_row[ 168 ][2],
   col_row[ 169 ][0],
   col_row[ 169 ][1],
   col_row[ 169 ][2],
   col_row[ 170 ][0],
   col_row[ 170 ][1],
   col_row[ 170 ][2],
   col_row[ 171 ][0],
   col_row[ 171 ][1],
   col_row[ 171 ][2],
   col_row[ 172 ][0],
   col_row[ 172 ][1],
   col_row[ 172 ][2],
   col_row[ 173 ][0],
   col_row[ 173 ][1],
   col_row[ 173 ][2],
   col_row[ 174 ][0],
   col_row[ 174 ][1],
   col_row[ 174 ][2],
   col_row[ 175 ][0],
   col_row[ 175 ][1],
   col_row[ 175 ][2],
   col_row[ 176 ][0],
   col_row[ 176 ][1],
   col_row[ 176 ][2],
   col_row[ 177 ][0],
   col_row[ 177 ][1],
   col_row[ 177 ][2],
   col_row[ 178 ][0],
   col_row[ 178 ][1],
   col_row[ 178 ][2],
   col_row[ 179 ][0],
   col_row[ 179 ][1],
   col_row[ 179 ][2],
   col_row[ 180 ][0],
   col_row[ 180 ][1],
   col_row[ 180 ][2],
   col_row[ 181 ][0],
   col_row[ 181 ][1],
   col_row[ 181 ][2],
   col_row[ 182 ][0],
   col_row[ 182 ][1],
   col_row[ 182 ][2],
   col_row[ 183 ][0],
   col_row[ 183 ][1],
   col_row[ 183 ][2],
   col_row[ 184 ][0],
   col_row[ 184 ][1],
   col_row[ 184 ][2],
   col_row[ 185 ][0],
   col_row[ 185 ][1],
   col_row[ 185 ][2],
   col_row[ 186 ][0],
   col_row[ 186 ][1],
   col_row[ 186 ][2],
   col_row[ 187 ][0],
   col_row[ 187 ][1],
   col_row[ 187 ][2],
   col_row[ 188 ][0],
   col_row[ 188 ][1],
   col_row[ 188 ][2],
   col_row[ 189 ][0],
   col_row[ 189 ][1],
   col_row[ 189 ][2],
   col_row[ 190 ][0],
   col_row[ 190 ][1],
   col_row[ 190 ][2],
   col_row[ 191 ][0],
   col_row[ 191 ][1],
   col_row[ 191 ][2],
   col_row[ 192 ][0],
   col_row[ 192 ][1],
   col_row[ 192 ][2],
   col_row[ 193 ][0],
   col_row[ 193 ][1],
   col_row[ 193 ][2],
   col_row[ 194 ][0],
   col_row[ 194 ][1],
   col_row[ 194 ][2],
   col_row[ 195 ][0],
   col_row[ 195 ][1],
   col_row[ 195 ][2],
   col_row[ 196 ][0],
   col_row[ 196 ][1],
   col_row[ 196 ][2],
   col_row[ 197 ][0],
   col_row[ 197 ][1],
   col_row[ 197 ][2],
   col_row[ 198 ][0],
   col_row[ 198 ][1],
   col_row[ 198 ][2],
   col_row[ 199 ][0],
   col_row[ 199 ][1],
   col_row[ 199 ][2],
   col_row[ 200 ][0],
   col_row[ 200 ][1],
   col_row[ 200 ][2],
   col_row[ 201 ][0],
   col_row[ 201 ][1],
   col_row[ 201 ][2],
   col_row[ 202 ][0],
   col_row[ 202 ][1],
   col_row[ 202 ][2],
   col_row[ 203 ][0],
   col_row[ 203 ][1],
   col_row[ 203 ][2],
   col_row[ 204 ][0],
   col_row[ 204 ][1],
   col_row[ 204 ][2],
   col_row[ 205 ][0],
   col_row[ 205 ][1],
   col_row[ 205 ][2],
   col_row[ 206 ][0],
   col_row[ 206 ][1],
   col_row[ 206 ][2],
   col_row[ 207 ][0],
   col_row[ 207 ][1],
   col_row[ 207 ][2],
   col_row[ 208 ][0],
   col_row[ 208 ][1],
   col_row[ 208 ][2],
   col_row[ 209 ][0],
   col_row[ 209 ][1],
   col_row[ 209 ][2],
   col_row[ 210 ][0],
   col_row[ 210 ][1],
   col_row[ 210 ][2],
   col_row[ 211 ][0],
   col_row[ 211 ][1],
   col_row[ 211 ][2],
   col_row[ 212 ][0],
   col_row[ 212 ][1],
   col_row[ 212 ][2],
   col_row[ 213 ][0],
   col_row[ 213 ][1],
   col_row[ 213 ][2],
   col_row[ 214 ][0],
   col_row[ 214 ][1],
   col_row[ 214 ][2],
   col_row[ 215 ][0],
   col_row[ 215 ][1],
   col_row[ 215 ][2],
   col_row[ 216 ][0],
   col_row[ 216 ][1],
   col_row[ 216 ][2],
   col_row[ 217 ][0],
   col_row[ 217 ][1],
   col_row[ 217 ][2],
   col_row[ 218 ][0],
   col_row[ 218 ][1],
   col_row[ 218 ][2],
   col_row[ 219 ][0],
   col_row[ 219 ][1],
   col_row[ 219 ][2],
   col_row[ 220 ][0],
   col_row[ 220 ][1],
   col_row[ 220 ][2],
   col_row[ 221 ][0],
   col_row[ 221 ][1],
   col_row[ 221 ][2],
   col_row[ 222 ][0],
   col_row[ 222 ][1],
   col_row[ 222 ][2],
   col_row[ 223 ][0],
   col_row[ 223 ][1],
   col_row[ 223 ][2],
   col_row[ 224 ][0],
   col_row[ 224 ][1],
   col_row[ 224 ][2],
   col_row[ 225 ][0],
   col_row[ 225 ][1],
   col_row[ 225 ][2],
   col_row[ 226 ][0],
   col_row[ 226 ][1],
   col_row[ 226 ][2],
   col_row[ 227 ][0],
   col_row[ 227 ][1],
   col_row[ 227 ][2],
   col_row[ 228 ][0],
   col_row[ 228 ][1],
   col_row[ 228 ][2],
   col_row[ 229 ][0],
   col_row[ 229 ][1],
   col_row[ 229 ][2],
   col_row[ 230 ][0],
   col_row[ 230 ][1],
   col_row[ 230 ][2],
   col_row[ 231 ][0],
   col_row[ 231 ][1],
   col_row[ 231 ][2],
   col_row[ 232 ][0],
   col_row[ 232 ][1],
   col_row[ 232 ][2],
   col_row[ 233 ][0],
   col_row[ 233 ][1],
   col_row[ 233 ][2],
   col_row[ 234 ][0],
   col_row[ 234 ][1],
   col_row[ 234 ][2],
   col_row[ 235 ][0],
   col_row[ 235 ][1],
   col_row[ 235 ][2],
   col_row[ 236 ][0],
   col_row[ 236 ][1],
   col_row[ 236 ][2],
   col_row[ 237 ][0],
   col_row[ 237 ][1],
   col_row[ 237 ][2],
   col_row[ 238 ][0],
   col_row[ 238 ][1],
   col_row[ 238 ][2],
   col_row[ 239 ][0],
   col_row[ 239 ][1],
   col_row[ 239 ][2],
   col_row[ 240 ][0],
   col_row[ 240 ][1],
   col_row[ 240 ][2],
   col_row[ 241 ][0],
   col_row[ 241 ][1],
   col_row[ 241 ][2],
   col_row[ 242 ][0],
   col_row[ 242 ][1],
   col_row[ 242 ][2],
   col_row[ 243 ][0],
   col_row[ 243 ][1],
   col_row[ 243 ][2],
   col_row[ 244 ][0],
   col_row[ 244 ][1],
   col_row[ 244 ][2],
   col_row[ 245 ][0],
   col_row[ 245 ][1],
   col_row[ 245 ][2],
   col_row[ 246 ][0],
   col_row[ 246 ][1],
   col_row[ 246 ][2],
   col_row[ 247 ][0],
   col_row[ 247 ][1],
   col_row[ 247 ][2],
   col_row[ 248 ][0],
   col_row[ 248 ][1],
   col_row[ 248 ][2],
   col_row[ 249 ][0],
   col_row[ 249 ][1],
   col_row[ 249 ][2],
   col_row[ 250 ][0],
   col_row[ 250 ][1],
   col_row[ 250 ][2],
   col_row[ 251 ][0],
   col_row[ 251 ][1],
   col_row[ 251 ][2],
   col_row[ 252 ][0],
   col_row[ 252 ][1],
   col_row[ 252 ][2],
   col_row[ 253 ][0],
   col_row[ 253 ][1],
   col_row[ 253 ][2],
   col_row[ 254 ][0],
   col_row[ 254 ][1],
   col_row[ 254 ][2],
   col_row[ 255 ][0],
   col_row[ 255 ][1],
   col_row[ 255 ][2],H[0][0],
   H[0][1],
   H[0][256],
   H[1][1],
   H[1][2],
   H[1][257],
   H[2][2],
   H[2][3],
   H[2][258],
   H[3][3],
   H[3][4],
   H[3][259],
   H[4][4],
   H[4][5],
   H[4][260],
   H[5][5],
   H[5][6],
   H[5][261],
   H[6][6],
   H[6][7],
   H[6][262],
   H[7][7],
   H[7][8],
   H[7][263],
   H[8][8],
   H[8][9],
   H[8][264],
   H[9][9],
   H[9][10],
   H[9][265],
   H[10][10],
   H[10][11],
   H[10][266],
   H[11][11],
   H[11][12],
   H[11][267],
   H[12][12],
   H[12][13],
   H[12][268],
   H[13][13],
   H[13][14],
   H[13][269],
   H[14][14],
   H[14][15],
   H[14][270],
   H[15][15],
   H[15][16],
   H[15][271],
   H[16][16],
   H[16][17],
   H[16][272],
   H[17][17],
   H[17][18],
   H[17][273],
   H[18][18],
   H[18][19],
   H[18][274],
   H[19][19],
   H[19][20],
   H[19][275],
   H[20][20],
   H[20][21],
   H[20][276],
   H[21][21],
   H[21][22],
   H[21][277],
   H[22][22],
   H[22][23],
   H[22][278],
   H[23][23],
   H[23][24],
   H[23][279],
   H[24][24],
   H[24][25],
   H[24][280],
   H[25][25],
   H[25][26],
   H[25][281],
   H[26][26],
   H[26][27],
   H[26][282],
   H[27][27],
   H[27][28],
   H[27][283],
   H[28][28],
   H[28][29],
   H[28][284],
   H[29][29],
   H[29][30],
   H[29][285],
   H[30][30],
   H[30][31],
   H[30][286],
   H[31][31],
   H[31][32],
   H[31][287],
   H[32][32],
   H[32][33],
   H[32][288],
   H[33][33],
   H[33][34],
   H[33][289],
   H[34][34],
   H[34][35],
   H[34][290],
   H[35][35],
   H[35][36],
   H[35][291],
   H[36][36],
   H[36][37],
   H[36][292],
   H[37][37],
   H[37][38],
   H[37][293],
   H[38][38],
   H[38][39],
   H[38][294],
   H[39][39],
   H[39][40],
   H[39][295],
   H[40][40],
   H[40][41],
   H[40][296],
   H[41][41],
   H[41][42],
   H[41][297],
   H[42][42],
   H[42][43],
   H[42][298],
   H[43][43],
   H[43][44],
   H[43][299],
   H[44][44],
   H[44][45],
   H[44][300],
   H[45][45],
   H[45][46],
   H[45][301],
   H[46][46],
   H[46][47],
   H[46][302],
   H[47][47],
   H[47][48],
   H[47][303],
   H[48][48],
   H[48][49],
   H[48][304],
   H[49][49],
   H[49][50],
   H[49][305],
   H[50][50],
   H[50][51],
   H[50][306],
   H[51][51],
   H[51][52],
   H[51][307],
   H[52][52],
   H[52][53],
   H[52][308],
   H[53][53],
   H[53][54],
   H[53][309],
   H[54][54],
   H[54][55],
   H[54][310],
   H[55][55],
   H[55][56],
   H[55][311],
   H[56][56],
   H[56][57],
   H[56][312],
   H[57][57],
   H[57][58],
   H[57][313],
   H[58][58],
   H[58][59],
   H[58][314],
   H[59][59],
   H[59][60],
   H[59][315],
   H[60][60],
   H[60][61],
   H[60][316],
   H[61][61],
   H[61][62],
   H[61][317],
   H[62][62],
   H[62][63],
   H[62][318],
   H[63][63],
   H[63][64],
   H[63][319],
   H[64][64],
   H[64][65],
   H[64][320],
   H[65][65],
   H[65][66],
   H[65][321],
   H[66][66],
   H[66][67],
   H[66][322],
   H[67][67],
   H[67][68],
   H[67][323],
   H[68][68],
   H[68][69],
   H[68][324],
   H[69][69],
   H[69][70],
   H[69][325],
   H[70][70],
   H[70][71],
   H[70][326],
   H[71][71],
   H[71][72],
   H[71][327],
   H[72][72],
   H[72][73],
   H[72][328],
   H[73][73],
   H[73][74],
   H[73][329],
   H[74][74],
   H[74][75],
   H[74][330],
   H[75][75],
   H[75][76],
   H[75][331],
   H[76][76],
   H[76][77],
   H[76][332],
   H[77][77],
   H[77][78],
   H[77][333],
   H[78][78],
   H[78][79],
   H[78][334],
   H[79][79],
   H[79][80],
   H[79][335],
   H[80][80],
   H[80][81],
   H[80][336],
   H[81][81],
   H[81][82],
   H[81][337],
   H[82][82],
   H[82][83],
   H[82][338],
   H[83][83],
   H[83][84],
   H[83][339],
   H[84][84],
   H[84][85],
   H[84][340],
   H[85][85],
   H[85][86],
   H[85][341],
   H[86][86],
   H[86][87],
   H[86][342],
   H[87][87],
   H[87][88],
   H[87][343],
   H[88][88],
   H[88][89],
   H[88][344],
   H[89][89],
   H[89][90],
   H[89][345],
   H[90][90],
   H[90][91],
   H[90][346],
   H[91][91],
   H[91][92],
   H[91][347],
   H[92][92],
   H[92][93],
   H[92][348],
   H[93][93],
   H[93][94],
   H[93][349],
   H[94][94],
   H[94][95],
   H[94][350],
   H[95][95],
   H[95][96],
   H[95][351],
   H[96][96],
   H[96][97],
   H[96][352],
   H[97][97],
   H[97][98],
   H[97][353],
   H[98][98],
   H[98][99],
   H[98][354],
   H[99][99],
   H[99][100],
   H[99][355],
   H[100][100],
   H[100][101],
   H[100][356],
   H[101][101],
   H[101][102],
   H[101][357],
   H[102][102],
   H[102][103],
   H[102][358],
   H[103][103],
   H[103][104],
   H[103][359],
   H[104][104],
   H[104][105],
   H[104][360],
   H[105][105],
   H[105][106],
   H[105][361],
   H[106][106],
   H[106][107],
   H[106][362],
   H[107][107],
   H[107][108],
   H[107][363],
   H[108][108],
   H[108][109],
   H[108][364],
   H[109][109],
   H[109][110],
   H[109][365],
   H[110][110],
   H[110][111],
   H[110][366],
   H[111][111],
   H[111][112],
   H[111][367],
   H[112][112],
   H[112][113],
   H[112][368],
   H[113][113],
   H[113][114],
   H[113][369],
   H[114][114],
   H[114][115],
   H[114][370],
   H[115][115],
   H[115][116],
   H[115][371],
   H[116][116],
   H[116][117],
   H[116][372],
   H[117][117],
   H[117][118],
   H[117][373],
   H[118][118],
   H[118][119],
   H[118][374],
   H[119][119],
   H[119][120],
   H[119][375],
   H[120][120],
   H[120][121],
   H[120][376],
   H[121][121],
   H[121][122],
   H[121][377],
   H[122][122],
   H[122][123],
   H[122][378],
   H[123][123],
   H[123][124],
   H[123][379],
   H[124][124],
   H[124][125],
   H[124][380],
   H[125][125],
   H[125][126],
   H[125][381],
   H[126][126],
   H[126][127],
   H[126][382],
   H[127][0],
   H[127][127],
   H[127][383],
   H[128][128],
   H[128][129],
   H[128][334],
   H[129][129],
   H[129][130],
   H[129][268],
   H[130][130],
   H[130][131],
   H[130][359],
   H[131][131],
   H[131][132],
   H[131][342],
   H[132][132],
   H[132][133],
   H[132][257],
   H[133][133],
   H[133][134],
   H[133][320],
   H[134][134],
   H[134][135],
   H[134][297],
   H[135][135],
   H[135][136],
   H[135][264],
   H[136][136],
   H[136][137],
   H[136][326],
   H[137][137],
   H[137][138],
   H[137][355],
   H[138][138],
   H[138][139],
   H[138][289],
   H[139][139],
   H[139][140],
   H[139][314],
   H[140][140],
   H[140][141],
   H[140][336],
   H[141][141],
   H[141][142],
   H[141][256],
   H[142][142],
   H[142][143],
   H[142][277],
   H[143][143],
   H[143][144],
   H[143][350],
   H[144][144],
   H[144][145],
   H[144][307],
   H[145][145],
   H[145][146],
   H[145][266],
   H[146][146],
   H[146][147],
   H[146][363],
   H[147][147],
   H[147][148],
   H[147][300],
   H[148][148],
   H[148][149],
   H[148][259],
   H[149][149],
   H[149][150],
   H[149][325],
   H[150][150],
   H[150][151],
   H[150][293],
   H[151][151],
   H[151][152],
   H[151][367],
   H[152][152],
   H[152][153],
   H[152][269],
   H[153][153],
   H[153][154],
   H[153][278],
   H[154][154],
   H[154][155],
   H[154][339],
   H[155][155],
   H[155][156],
   H[155][322],
   H[156][156],
   H[156][157],
   H[156][261],
   H[157][157],
   H[157][158],
   H[157][356],
   H[158][158],
   H[158][159],
   H[158][305],
   H[159][159],
   H[159][160],
   H[159][272],
   H[160][160],
   H[160][161],
   H[160][371],
   H[161][161],
   H[161][162],
   H[161][344],
   H[162][162],
   H[162][163],
   H[162][315],
   H[163][163],
   H[163][164],
   H[163][294],
   H[164][164],
   H[164][165],
   H[164][351],
   H[165][165],
   H[165][166],
   H[165][262],
   H[166][166],
   H[166][167],
   H[166][378],
   H[167][167],
   H[167][168],
   H[167][288],
   H[168][168],
   H[168][169],
   H[168][330],
   H[169][169],
   H[169][170],
   H[169][343],
   H[170][170],
   H[170][171],
   H[170][279],
   H[171][171],
   H[171][172],
   H[171][374],
   H[172][172],
   H[172][173],
   H[172][265],
   H[173][173],
   H[173][174],
   H[173][337],
   H[174][174],
   H[174][175],
   H[174][285],
   H[175][175],
   H[175][176],
   H[175][302],
   H[176][176],
   H[176][177],
   H[176][353],
   H[177][177],
   H[177][178],
   H[177][270],
   H[178][178],
   H[178][179],
   H[178][319],
   H[179][179],
   H[179][180],
   H[179][376],
   H[180][180],
   H[180][181],
   H[180][345],
   H[181][181],
   H[181][182],
   H[181][308],
   H[182][182],
   H[182][183],
   H[182][338],
   H[183][183],
   H[183][184],
   H[183][327],
   H[184][184],
   H[184][185],
   H[184][273],
   H[185][185],
   H[185][186],
   H[185][381],
   H[186][186],
   H[186][187],
   H[186][299],
   H[187][187],
   H[187][188],
   H[187][280],
   H[188][188],
   H[188][189],
   H[188][357],
   H[189][189],
   H[189][190],
   H[189][292],
   H[190][190],
   H[190][191],
   H[190][311],
   H[191][191],
   H[191][192],
   H[191][341],
   H[192][192],
   H[192][193],
   H[192][349],
   H[193][193],
   H[193][194],
   H[193][370],
   H[194][194],
   H[194][195],
   H[194][321],
   H[195][195],
   H[195][196],
   H[195][282],
   H[196][196],
   H[196][197],
   H[196][335],
   H[197][197],
   H[197][198],
   H[197][306],
   H[198][198],
   H[198][199],
   H[198][295],
   H[199][199],
   H[199][200],
   H[199][373],
   H[200][200],
   H[200][201],
   H[200][287],
   H[201][201],
   H[201][202],
   H[201][364],
   H[202][202],
   H[202][203],
   H[202][340],
   H[203][203],
   H[203][204],
   H[203][318],
   H[204][204],
   H[204][205],
   H[204][382],
   H[205][205],
   H[205][206],
   H[205][304],
   H[206][206],
   H[206][207],
   H[206][360],
   H[207][207],
   H[207][208],
   H[207][375],
   H[208][208],
   H[208][209],
   H[208][313],
   H[209][209],
   H[209][210],
   H[209][298],
   H[210][210],
   H[210][211],
   H[210][368],
   H[211][211],
   H[211][212],
   H[211][286],
   H[212][212],
   H[212][213],
   H[212][323],
   H[213][213],
   H[213][214],
   H[213][383],
   H[214][214],
   H[214][215],
   H[214][309],
   H[215][215],
   H[215][216],
   H[215][331],
   H[216][216],
   H[216][217],
   H[216][348],
   H[217][217],
   H[217][218],
   H[217][296],
   H[218][218],
   H[218][219],
   H[218][377],
   H[219][219],
   H[219][220],
   H[219][284],
   H[220][220],
   H[220][221],
   H[220][358],
   H[221][221],
   H[221][222],
   H[221][328],
   H[222][222],
   H[222][223],
   H[222][372],
   H[223][223],
   H[223][224],
   H[223][276],
   H[224][224],
   H[224][225],
   H[224][301],
   H[225][225],
   H[225][226],
   H[225][316],
   H[226][226],
   H[226][227],
   H[226][332],
   H[227][227],
   H[227][228],
   H[227][380],
   H[228][228],
   H[228][229],
   H[228][291],
   H[229][229],
   H[229][230],
   H[229][362],
   H[230][230],
   H[230][231],
   H[230][283],
   H[231][231],
   H[231][232],
   H[231][274],
   H[232][232],
   H[232][233],
   H[232][346],
   H[233][233],
   H[233][234],
   H[233][354],
   H[234][234],
   H[234][235],
   H[234][333],
   H[235][235],
   H[235][236],
   H[235][369],
   H[236][236],
   H[236][237],
   H[236][263],
   H[237][237],
   H[237][238],
   H[237][361],
   H[238][238],
   H[238][239],
   H[238][271],
   H[239][239],
   H[239][240],
   H[239][310],
   H[240][240],
   H[240][241],
   H[240][379],
   H[241][241],
   H[241][242],
   H[241][366],
   H[242][242],
   H[242][243],
   H[242][281],
   H[243][243],
   H[243][244],
   H[243][260],
   H[244][244],
   H[244][245],
   H[244][317],
   H[245][245],
   H[245][246],
   H[245][347],
   H[246][246],
   H[246][247],
   H[246][267],
   H[247][247],
   H[247][248],
   H[247][290],
   H[248][248],
   H[248][249],
   H[248][303],
   H[249][249],
   H[249][250],
   H[249][365],
   H[250][250],
   H[250][251],
   H[250][329],
   H[251][251],
   H[251][252],
   H[251][258],
   H[252][252],
   H[252][253],
   H[252][352],
   H[253][253],
   H[253][254],
   H[253][312],
   H[254][254],
   H[254][255],
   H[254][275],
   H[255][128],
   H[255][255],
   H[255][324],



addrA_[0],
addrA_[1],
addrA_[2],
addrA_[3],
addrA_[4],
addrA_[5],
addrA_[6],
addrA_[7],
addrA_[8],
addrA_[9],
addrA_[10],
addrA_[11],
addrA_[12],
addrA_[13],
addrA_[14],
addrA_[15],
addrA_[16],
addrA_[17],
addrA_[18],
addrA_[19],
addrA_[20],
addrA_[21],
addrA_[22],
addrA_[23],
addrA_[24],
addrA_[25],
addrA_[26],
addrA_[27],
addrA_[28],
addrA_[29],
addrA_[30],
addrA_[31],
addrA_[32],
addrA_[33],
addrA_[34],
addrA_[35],
addrA_[36],
addrA_[37],
addrA_[38],
addrA_[39],
addrA_[40],
addrA_[41],
addrA_[42],
addrA_[43],
addrA_[44],
addrA_[45],
addrA_[46],
addrA_[47],
addrA_[48],
addrA_[49],
addrA_[50],
addrA_[51],
addrA_[52],
addrA_[53],
addrA_[54],
addrA_[55],
addrA_[56],
addrA_[57],
addrA_[58],
addrA_[59],
addrA_[60],
addrA_[61],
addrA_[62],
addrA_[63],
addrA_[64],
addrA_[65],
addrA_[66],
addrA_[67],
addrA_[68],
addrA_[69],
addrA_[70],
addrA_[71],
addrA_[72],
addrA_[73],
addrA_[74],
addrA_[75],
addrA_[76],
addrA_[77],
addrA_[78],
addrA_[79],
addrA_[80],
addrA_[81],
addrA_[82],
addrA_[83],
addrA_[84],
addrA_[85],
addrA_[86],
addrA_[87],
addrA_[88],
addrA_[89],
addrA_[90],
addrA_[91],
addrA_[92],
addrA_[93],
addrA_[94],
addrA_[95],
addrA_[96],
addrA_[97],
addrA_[98],
addrA_[99],
addrA_[100],
addrA_[101],
addrA_[102],
addrA_[103],
addrA_[104],
addrA_[105],
addrA_[106],
addrA_[107],
addrA_[108],
addrA_[109],
addrA_[110],
addrA_[111],
addrA_[112],
addrA_[113],
addrA_[114],
addrA_[115],
addrA_[116],
addrA_[117],
addrA_[118],
addrA_[119],
addrA_[120],
addrA_[121],
addrA_[122],
addrA_[123],
addrA_[124],
addrA_[125],
addrA_[126],
addrA_[127],
addrA_[128],
addrA_[129],
addrA_[130],
addrA_[131],
addrA_[132],
addrA_[133],
addrA_[134],
addrA_[135],
addrA_[136],
addrA_[137],
addrA_[138],
addrA_[139],
addrA_[140],
addrA_[141],
addrA_[142],
addrA_[143],
addrA_[144],
addrA_[145],
addrA_[146],
addrA_[147],
addrA_[148],
addrA_[149],
addrA_[150],
addrA_[151],
addrA_[152],
addrA_[153],
addrA_[154],
addrA_[155],
addrA_[156],
addrA_[157],
addrA_[158],
addrA_[159],
addrA_[160],
addrA_[161],
addrA_[162],
addrA_[163],
addrA_[164],
addrA_[165],
addrA_[166],
addrA_[167],
addrA_[168],
addrA_[169],
addrA_[170],
addrA_[171],
addrA_[172],
addrA_[173],
addrA_[174],
addrA_[175],
addrA_[176],
addrA_[177],
addrA_[178],
addrA_[179],
addrA_[180],
addrA_[181],
addrA_[182],
addrA_[183],
addrA_[184],
addrA_[185],
addrA_[186],
addrA_[187],
addrA_[188],
addrA_[189],
addrA_[190],
addrA_[191],
addrA_[192],
addrA_[193],
addrA_[194],
addrA_[195],
addrA_[196],
addrA_[197],
addrA_[198],
addrA_[199],
addrA_[200],
addrA_[201],
addrA_[202],
addrA_[203],
addrA_[204],
addrA_[205],
addrA_[206],
addrA_[207],
addrA_[208],
addrA_[209],
addrA_[210],
addrA_[211],
addrA_[212],
addrA_[213],
addrA_[214],
addrA_[215],
addrA_[216],
addrA_[217],
addrA_[218],
addrA_[219],
addrA_[220],
addrA_[221],
addrA_[222],
addrA_[223],
addrA_[224],
addrA_[225],
addrA_[226],
addrA_[227],
addrA_[228],
addrA_[229],
addrA_[230],
addrA_[231],
addrA_[232],
addrA_[233],
addrA_[234],
addrA_[235],
addrA_[236],
addrA_[237],
addrA_[238],
addrA_[239],
addrA_[240],
addrA_[241],
addrA_[242],
addrA_[243],
addrA_[244],
addrA_[245],
addrA_[246],
addrA_[247],
addrA_[248],
addrA_[249],
addrA_[250],
addrA_[251],
addrA_[252],
addrA_[253],
addrA_[254],
addrA_[255],
addrA_[256],
addrA_[257],
addrA_[258],
addrA_[259],
addrA_[260],
addrA_[261],
addrA_[262],
addrA_[263],
addrA_[264],
addrA_[265],
addrA_[266],
addrA_[267],
addrA_[268],
addrA_[269],
addrA_[270],
addrA_[271],
addrA_[272],
addrA_[273],
addrA_[274],
addrA_[275],
addrA_[276],
addrA_[277],
addrA_[278],
addrA_[279],
addrA_[280],
addrA_[281],
addrA_[282],
addrA_[283],
addrA_[284],
addrA_[285],
addrA_[286],
addrA_[287],
addrA_[288],
addrA_[289],
addrA_[290],
addrA_[291],
addrA_[292],
addrA_[293],
addrA_[294],
addrA_[295],
addrA_[296],
addrA_[297],
addrA_[298],
addrA_[299],
addrA_[300],
addrA_[301],
addrA_[302],
addrA_[303],
addrA_[304],
addrA_[305],
addrA_[306],
addrA_[307],
addrA_[308],
addrA_[309],
addrA_[310],
addrA_[311],
addrA_[312],
addrA_[313],
addrA_[314],
addrA_[315],
addrA_[316],
addrA_[317],
addrA_[318],
addrA_[319],
addrA_[320],
addrA_[321],
addrA_[322],
addrA_[323],
addrA_[324],
addrA_[325],
addrA_[326],
addrA_[327],
addrA_[328],
addrA_[329],
addrA_[330],
addrA_[331],
addrA_[332],
addrA_[333],
addrA_[334],
addrA_[335],
addrA_[336],
addrA_[337],
addrA_[338],
addrA_[339],
addrA_[340],
addrA_[341],
addrA_[342],
addrA_[343],
addrA_[344],
addrA_[345],
addrA_[346],
addrA_[347],
addrA_[348],
addrA_[349],
addrA_[350],
addrA_[351],
addrA_[352],
addrA_[353],
addrA_[354],
addrA_[355],
addrA_[356],
addrA_[357],
addrA_[358],
addrA_[359],
addrA_[360],
addrA_[361],
addrA_[362],
addrA_[363],
addrA_[364],
addrA_[365],
addrA_[366],
addrA_[367],
addrA_[368],
addrA_[369],
addrA_[370],
addrA_[371],
addrA_[372],
addrA_[373],
addrA_[374],
addrA_[375],
addrA_[376],
addrA_[377],
addrA_[378],
addrA_[379],
addrA_[380],
addrA_[381],
addrA_[382],
addrA_[383],
addrA_[384],
addrA_[385],
addrA_[386],
addrA_[387],
addrA_[388],
addrA_[389],
addrA_[390],
addrA_[391],
addrA_[392],
addrA_[393],
addrA_[394],
addrA_[395],
addrA_[396],
addrA_[397],
addrA_[398],
addrA_[399],
addrA_[400],
addrA_[401],
addrA_[402],
addrA_[403],
addrA_[404],
addrA_[405],
addrA_[406],
addrA_[407],
addrA_[408],
addrA_[409],
addrA_[410],
addrA_[411],
addrA_[412],
addrA_[413],
addrA_[414],
addrA_[415],
addrA_[416],
addrA_[417],
addrA_[418],
addrA_[419],
addrA_[420],
addrA_[421],
addrA_[422],
addrA_[423],
addrA_[424],
addrA_[425],
addrA_[426],
addrA_[427],
addrA_[428],
addrA_[429],
addrA_[430],
addrA_[431],
addrA_[432],
addrA_[433],
addrA_[434],
addrA_[435],
addrA_[436],
addrA_[437],
addrA_[438],
addrA_[439],
addrA_[440],
addrA_[441],
addrA_[442],
addrA_[443],
addrA_[444],
addrA_[445],
addrA_[446],
addrA_[447],
addrA_[448],
addrA_[449],
addrA_[450],
addrA_[451],
addrA_[452],
addrA_[453],
addrA_[454],
addrA_[455],
addrA_[456],
addrA_[457],
addrA_[458],
addrA_[459],
addrA_[460],
addrA_[461],
addrA_[462],
addrA_[463],
addrA_[464],
addrA_[465],
addrA_[466],
addrA_[467],
addrA_[468],
addrA_[469],
addrA_[470],
addrA_[471],
addrA_[472],
addrA_[473],
addrA_[474],
addrA_[475],
addrA_[476],
addrA_[477],
addrA_[478],
addrA_[479],
addrA_[480],
addrA_[481],
addrA_[482],
addrA_[483],
addrA_[484],
addrA_[485],
addrA_[486],
addrA_[487],
addrA_[488],
addrA_[489],
addrA_[490],
addrA_[491],
addrA_[492],
addrA_[493],
addrA_[494],
addrA_[495],
addrA_[496],
addrA_[497],
addrA_[498],
addrA_[499],
addrA_[500],
addrA_[501],
addrA_[502],
addrA_[503],
addrA_[504],
addrA_[505],
addrA_[506],
addrA_[507],
addrA_[508],
addrA_[509],
addrA_[510],
addrA_[511],
addrA_[512],
addrA_[513],
addrA_[514],
addrA_[515],
addrA_[516],
addrA_[517],
addrA_[518],
addrA_[519],
addrA_[520],
addrA_[521],
addrA_[522],
addrA_[523],
addrA_[524],
addrA_[525],
addrA_[526],
addrA_[527],
addrA_[528],
addrA_[529],
addrA_[530],
addrA_[531],
addrA_[532],
addrA_[533],
addrA_[534],
addrA_[535],
addrA_[536],
addrA_[537],
addrA_[538],
addrA_[539],
addrA_[540],
addrA_[541],
addrA_[542],
addrA_[543],
addrA_[544],
addrA_[545],
addrA_[546],
addrA_[547],
addrA_[548],
addrA_[549],
addrA_[550],
addrA_[551],
addrA_[552],
addrA_[553],
addrA_[554],
addrA_[555],
addrA_[556],
addrA_[557],
addrA_[558],
addrA_[559],
addrA_[560],
addrA_[561],
addrA_[562],
addrA_[563],
addrA_[564],
addrA_[565],
addrA_[566],
addrA_[567],
addrA_[568],
addrA_[569],
addrA_[570],
addrA_[571],
addrA_[572],
addrA_[573],
addrA_[574],
addrA_[575],
addrA_[576],
addrA_[577],
addrA_[578],
addrA_[579],
addrA_[580],
addrA_[581],
addrA_[582],
addrA_[583],
addrA_[584],
addrA_[585],
addrA_[586],
addrA_[587],
addrA_[588],
addrA_[589],
addrA_[590],
addrA_[591],
addrA_[592],
addrA_[593],
addrA_[594],
addrA_[595],
addrA_[596],
addrA_[597],
addrA_[598],
addrA_[599],
addrA_[600],
addrA_[601],
addrA_[602],
addrA_[603],
addrA_[604],
addrA_[605],
addrA_[606],
addrA_[607],
addrA_[608],
addrA_[609],
addrA_[610],
addrA_[611],
addrA_[612],
addrA_[613],
addrA_[614],
addrA_[615],
addrA_[616],
addrA_[617],
addrA_[618],
addrA_[619],
addrA_[620],
addrA_[621],
addrA_[622],
addrA_[623],
addrA_[624],
addrA_[625],
addrA_[626],
addrA_[627],
addrA_[628],
addrA_[629],
addrA_[630],
addrA_[631],
addrA_[632],
addrA_[633],
addrA_[634],
addrA_[635],
addrA_[636],
addrA_[637],
addrA_[638],
addrA_[639],
addrA_[640],
addrA_[641],
addrA_[642],
addrA_[643],
addrA_[644],
addrA_[645],
addrA_[646],
addrA_[647],
addrA_[648],
addrA_[649],
addrA_[650],
addrA_[651],
addrA_[652],
addrA_[653],
addrA_[654],
addrA_[655],
addrA_[656],
addrA_[657],
addrA_[658],
addrA_[659],
addrA_[660],
addrA_[661],
addrA_[662],
addrA_[663],
addrA_[664],
addrA_[665],
addrA_[666],
addrA_[667],
addrA_[668],
addrA_[669],
addrA_[670],
addrA_[671],
addrA_[672],
addrA_[673],
addrA_[674],
addrA_[675],
addrA_[676],
addrA_[677],
addrA_[678],
addrA_[679],
addrA_[680],
addrA_[681],
addrA_[682],
addrA_[683],
addrA_[684],
addrA_[685],
addrA_[686],
addrA_[687],
addrA_[688],
addrA_[689],
addrA_[690],
addrA_[691],
addrA_[692],
addrA_[693],
addrA_[694],
addrA_[695],
addrA_[696],
addrA_[697],
addrA_[698],
addrA_[699],
addrA_[700],
addrA_[701],
addrA_[702],
addrA_[703],
addrA_[704],
addrA_[705],
addrA_[706],
addrA_[707],
addrA_[708],
addrA_[709],
addrA_[710],
addrA_[711],
addrA_[712],
addrA_[713],
addrA_[714],
addrA_[715],
addrA_[716],
addrA_[717],
addrA_[718],
addrA_[719],
addrA_[720],
addrA_[721],
addrA_[722],
addrA_[723],
addrA_[724],
addrA_[725],
addrA_[726],
addrA_[727],
addrA_[728],
addrA_[729],
addrA_[730],
addrA_[731],
addrA_[732],
addrA_[733],
addrA_[734],
addrA_[735],
addrA_[736],
addrA_[737],
addrA_[738],
addrA_[739],
addrA_[740],
addrA_[741],
addrA_[742],
addrA_[743],
addrA_[744],
addrA_[745],
addrA_[746],
addrA_[747],
addrA_[748],
addrA_[749],
addrA_[750],
addrA_[751],
addrA_[752],
addrA_[753],
addrA_[754],
addrA_[755],
addrA_[756],
addrA_[757],
addrA_[758],
addrA_[759],
addrA_[760],
addrA_[761],
addrA_[762],
addrA_[763],
addrA_[764],
addrA_[765],
addrA_[766],
addrA_[767],


   doutA[0],
doutA[1],
doutA[2],
doutA[3],
doutA[4],
doutA[5],
doutA[6],
doutA[7],
doutA[8],
doutA[9],
doutA[10],
doutA[11],
doutA[12],
doutA[13],
doutA[14],
doutA[15],
doutA[16],
doutA[17],
doutA[18],
doutA[19],
doutA[20],
doutA[21],
doutA[22],
doutA[23],
doutA[24],
doutA[25],
doutA[26],
doutA[27],
doutA[28],
doutA[29],
doutA[30],
doutA[31],
doutA[32],
doutA[33],
doutA[34],
doutA[35],
doutA[36],
doutA[37],
doutA[38],
doutA[39],
doutA[40],
doutA[41],
doutA[42],
doutA[43],
doutA[44],
doutA[45],
doutA[46],
doutA[47],
doutA[48],
doutA[49],
doutA[50],
doutA[51],
doutA[52],
doutA[53],
doutA[54],
doutA[55],
doutA[56],
doutA[57],
doutA[58],
doutA[59],
doutA[60],
doutA[61],
doutA[62],
doutA[63],
doutA[64],
doutA[65],
doutA[66],
doutA[67],
doutA[68],
doutA[69],
doutA[70],
doutA[71],
doutA[72],
doutA[73],
doutA[74],
doutA[75],
doutA[76],
doutA[77],
doutA[78],
doutA[79],
doutA[80],
doutA[81],
doutA[82],
doutA[83],
doutA[84],
doutA[85],
doutA[86],
doutA[87],
doutA[88],
doutA[89],
doutA[90],
doutA[91],
doutA[92],
doutA[93],
doutA[94],
doutA[95],
doutA[96],
doutA[97],
doutA[98],
doutA[99],
doutA[100],
doutA[101],
doutA[102],
doutA[103],
doutA[104],
doutA[105],
doutA[106],
doutA[107],
doutA[108],
doutA[109],
doutA[110],
doutA[111],
doutA[112],
doutA[113],
doutA[114],
doutA[115],
doutA[116],
doutA[117],
doutA[118],
doutA[119],
doutA[120],
doutA[121],
doutA[122],
doutA[123],
doutA[124],
doutA[125],
doutA[126],
doutA[127],
doutA[128],
doutA[129],
doutA[130],
doutA[131],
doutA[132],
doutA[133],
doutA[134],
doutA[135],
doutA[136],
doutA[137],
doutA[138],
doutA[139],
doutA[140],
doutA[141],
doutA[142],
doutA[143],
doutA[144],
doutA[145],
doutA[146],
doutA[147],
doutA[148],
doutA[149],
doutA[150],
doutA[151],
doutA[152],
doutA[153],
doutA[154],
doutA[155],
doutA[156],
doutA[157],
doutA[158],
doutA[159],
doutA[160],
doutA[161],
doutA[162],
doutA[163],
doutA[164],
doutA[165],
doutA[166],
doutA[167],
doutA[168],
doutA[169],
doutA[170],
doutA[171],
doutA[172],
doutA[173],
doutA[174],
doutA[175],
doutA[176],
doutA[177],
doutA[178],
doutA[179],
doutA[180],
doutA[181],
doutA[182],
doutA[183],
doutA[184],
doutA[185],
doutA[186],
doutA[187],
doutA[188],
doutA[189],
doutA[190],
doutA[191],
doutA[192],
doutA[193],
doutA[194],
doutA[195],
doutA[196],
doutA[197],
doutA[198],
doutA[199],
doutA[200],
doutA[201],
doutA[202],
doutA[203],
doutA[204],
doutA[205],
doutA[206],
doutA[207],
doutA[208],
doutA[209],
doutA[210],
doutA[211],
doutA[212],
doutA[213],
doutA[214],
doutA[215],
doutA[216],
doutA[217],
doutA[218],
doutA[219],
doutA[220],
doutA[221],
doutA[222],
doutA[223],
doutA[224],
doutA[225],
doutA[226],
doutA[227],
doutA[228],
doutA[229],
doutA[230],
doutA[231],
doutA[232],
doutA[233],
doutA[234],
doutA[235],
doutA[236],
doutA[237],
doutA[238],
doutA[239],
doutA[240],
doutA[241],
doutA[242],
doutA[243],
doutA[244],
doutA[245],
doutA[246],
doutA[247],
doutA[248],
doutA[249],
doutA[250],
doutA[251],
doutA[252],
doutA[253],
doutA[254],
doutA[255],
doutA[256],
doutA[257],
doutA[258],
doutA[259],
doutA[260],
doutA[261],
doutA[262],
doutA[263],
doutA[264],
doutA[265],
doutA[266],
doutA[267],
doutA[268],
doutA[269],
doutA[270],
doutA[271],
doutA[272],
doutA[273],
doutA[274],
doutA[275],
doutA[276],
doutA[277],
doutA[278],
doutA[279],
doutA[280],
doutA[281],
doutA[282],
doutA[283],
doutA[284],
doutA[285],
doutA[286],
doutA[287],
doutA[288],
doutA[289],
doutA[290],
doutA[291],
doutA[292],
doutA[293],
doutA[294],
doutA[295],
doutA[296],
doutA[297],
doutA[298],
doutA[299],
doutA[300],
doutA[301],
doutA[302],
doutA[303],
doutA[304],
doutA[305],
doutA[306],
doutA[307],
doutA[308],
doutA[309],
doutA[310],
doutA[311],
doutA[312],
doutA[313],
doutA[314],
doutA[315],
doutA[316],
doutA[317],
doutA[318],
doutA[319],
doutA[320],
doutA[321],
doutA[322],
doutA[323],
doutA[324],
doutA[325],
doutA[326],
doutA[327],
doutA[328],
doutA[329],
doutA[330],
doutA[331],
doutA[332],
doutA[333],
doutA[334],
doutA[335],
doutA[336],
doutA[337],
doutA[338],
doutA[339],
doutA[340],
doutA[341],
doutA[342],
doutA[343],
doutA[344],
doutA[345],
doutA[346],
doutA[347],
doutA[348],
doutA[349],
doutA[350],
doutA[351],
doutA[352],
doutA[353],
doutA[354],
doutA[355],
doutA[356],
doutA[357],
doutA[358],
doutA[359],
doutA[360],
doutA[361],
doutA[362],
doutA[363],
doutA[364],
doutA[365],
doutA[366],
doutA[367],
doutA[368],
doutA[369],
doutA[370],
doutA[371],
doutA[372],
doutA[373],
doutA[374],
doutA[375],
doutA[376],
doutA[377],
doutA[378],
doutA[379],
doutA[380],
doutA[381],
doutA[382],
doutA[383],
doutA[384],
doutA[385],
doutA[386],
doutA[387],
doutA[388],
doutA[389],
doutA[390],
doutA[391],
doutA[392],
doutA[393],
doutA[394],
doutA[395],
doutA[396],
doutA[397],
doutA[398],
doutA[399],
doutA[400],
doutA[401],
doutA[402],
doutA[403],
doutA[404],
doutA[405],
doutA[406],
doutA[407],
doutA[408],
doutA[409],
doutA[410],
doutA[411],
doutA[412],
doutA[413],
doutA[414],
doutA[415],
doutA[416],
doutA[417],
doutA[418],
doutA[419],
doutA[420],
doutA[421],
doutA[422],
doutA[423],
doutA[424],
doutA[425],
doutA[426],
doutA[427],
doutA[428],
doutA[429],
doutA[430],
doutA[431],
doutA[432],
doutA[433],
doutA[434],
doutA[435],
doutA[436],
doutA[437],
doutA[438],
doutA[439],
doutA[440],
doutA[441],
doutA[442],
doutA[443],
doutA[444],
doutA[445],
doutA[446],
doutA[447],
doutA[448],
doutA[449],
doutA[450],
doutA[451],
doutA[452],
doutA[453],
doutA[454],
doutA[455],
doutA[456],
doutA[457],
doutA[458],
doutA[459],
doutA[460],
doutA[461],
doutA[462],
doutA[463],
doutA[464],
doutA[465],
doutA[466],
doutA[467],
doutA[468],
doutA[469],
doutA[470],
doutA[471],
doutA[472],
doutA[473],
doutA[474],
doutA[475],
doutA[476],
doutA[477],
doutA[478],
doutA[479],
doutA[480],
doutA[481],
doutA[482],
doutA[483],
doutA[484],
doutA[485],
doutA[486],
doutA[487],
doutA[488],
doutA[489],
doutA[490],
doutA[491],
doutA[492],
doutA[493],
doutA[494],
doutA[495],
doutA[496],
doutA[497],
doutA[498],
doutA[499],
doutA[500],
doutA[501],
doutA[502],
doutA[503],
doutA[504],
doutA[505],
doutA[506],
doutA[507],
doutA[508],
doutA[509],
doutA[510],
doutA[511],
doutA[512],
doutA[513],
doutA[514],
doutA[515],
doutA[516],
doutA[517],
doutA[518],
doutA[519],
doutA[520],
doutA[521],
doutA[522],
doutA[523],
doutA[524],
doutA[525],
doutA[526],
doutA[527],
doutA[528],
doutA[529],
doutA[530],
doutA[531],
doutA[532],
doutA[533],
doutA[534],
doutA[535],
doutA[536],
doutA[537],
doutA[538],
doutA[539],
doutA[540],
doutA[541],
doutA[542],
doutA[543],
doutA[544],
doutA[545],
doutA[546],
doutA[547],
doutA[548],
doutA[549],
doutA[550],
doutA[551],
doutA[552],
doutA[553],
doutA[554],
doutA[555],
doutA[556],
doutA[557],
doutA[558],
doutA[559],
doutA[560],
doutA[561],
doutA[562],
doutA[563],
doutA[564],
doutA[565],
doutA[566],
doutA[567],
doutA[568],
doutA[569],
doutA[570],
doutA[571],
doutA[572],
doutA[573],
doutA[574],
doutA[575],
doutA[576],
doutA[577],
doutA[578],
doutA[579],
doutA[580],
doutA[581],
doutA[582],
doutA[583],
doutA[584],
doutA[585],
doutA[586],
doutA[587],
doutA[588],
doutA[589],
doutA[590],
doutA[591],
doutA[592],
doutA[593],
doutA[594],
doutA[595],
doutA[596],
doutA[597],
doutA[598],
doutA[599],
doutA[600],
doutA[601],
doutA[602],
doutA[603],
doutA[604],
doutA[605],
doutA[606],
doutA[607],
doutA[608],
doutA[609],
doutA[610],
doutA[611],
doutA[612],
doutA[613],
doutA[614],
doutA[615],
doutA[616],
doutA[617],
doutA[618],
doutA[619],
doutA[620],
doutA[621],
doutA[622],
doutA[623],
doutA[624],
doutA[625],
doutA[626],
doutA[627],
doutA[628],
doutA[629],
doutA[630],
doutA[631],
doutA[632],
doutA[633],
doutA[634],
doutA[635],
doutA[636],
doutA[637],
doutA[638],
doutA[639],
doutA[640],
doutA[641],
doutA[642],
doutA[643],
doutA[644],
doutA[645],
doutA[646],
doutA[647],
doutA[648],
doutA[649],
doutA[650],
doutA[651],
doutA[652],
doutA[653],
doutA[654],
doutA[655],
doutA[656],
doutA[657],
doutA[658],
doutA[659],
doutA[660],
doutA[661],
doutA[662],
doutA[663],
doutA[664],
doutA[665],
doutA[666],
doutA[667],
doutA[668],
doutA[669],
doutA[670],
doutA[671],
doutA[672],
doutA[673],
doutA[674],
doutA[675],
doutA[676],
doutA[677],
doutA[678],
doutA[679],
doutA[680],
doutA[681],
doutA[682],
doutA[683],
doutA[684],
doutA[685],
doutA[686],
doutA[687],
doutA[688],
doutA[689],
doutA[690],
doutA[691],
doutA[692],
doutA[693],
doutA[694],
doutA[695],
doutA[696],
doutA[697],
doutA[698],
doutA[699],
doutA[700],
doutA[701],
doutA[702],
doutA[703],
doutA[704],
doutA[705],
doutA[706],
doutA[707],
doutA[708],
doutA[709],
doutA[710],
doutA[711],
doutA[712],
doutA[713],
doutA[714],
doutA[715],
doutA[716],
doutA[717],
doutA[718],
doutA[719],
doutA[720],
doutA[721],
doutA[722],
doutA[723],
doutA[724],
doutA[725],
doutA[726],
doutA[727],
doutA[728],
doutA[729],
doutA[730],
doutA[731],
doutA[732],
doutA[733],
doutA[734],
doutA[735],
doutA[736],
doutA[737],
doutA[738],
doutA[739],
doutA[740],
doutA[741],
doutA[742],
doutA[743],
doutA[744],
doutA[745],
doutA[746],
doutA[747],
doutA[748],
doutA[749],
doutA[750],
doutA[751],
doutA[752],
doutA[753],
doutA[754],
doutA[755],
doutA[756],
doutA[757],
doutA[758],
doutA[759],
doutA[760],
doutA[761],
doutA[762],
doutA[763],
doutA[764],
doutA[765],
doutA[766],
doutA[767]


   )
begin
if(reset) begin
for(loop_var=0;loop_var<768;loop_var=loop_var+1) begin
weA[loop_var]=0;
addrA[loop_var]=0;
dinA[loop_var]=0;
weA1[loop_var]=0;
addrA1[loop_var]=0;
dinA1[loop_var]=0;
end


for(loop_var=0;loop_var<16;loop_var=loop_var+1) begin
for(loop_var1=0;loop_var1<3;loop_var1=loop_var1+1) begin
for(loop_var2=0;loop_var2<256;loop_var2=loop_var2+1) begin
F[loop_var][loop_var1][loop_var2]=0;
end
end
end


for(loop_var=0;loop_var<16;loop_var=loop_var+1) begin
for(loop_var1=0;loop_var1<3;loop_var1=loop_var1+1) begin
for(loop_var2=0;loop_var2<256;loop_var2=loop_var2+1) begin
B[loop_var][loop_var1][loop_var2]=0;
end
end
end


col_state=10'd0;
row_state=10'd0;

address=10'd0;
address1=4'd0;
out_enable=1'd0;
out=6'd0;
end
else begin
case(state)
`RESET_STATE: begin

end
`GAMMAIN0: begin
for(loop_var=0;loop_var<768;loop_var=loop_var+1) begin
dinA[loop_var]=GAM;
addrA[loop_var]=count[3:0];
weA[loop_var]=1'b1;
end
end

`GAMMAIN1: begin
for(loop_var=0;loop_var<768;loop_var=loop_var+1) begin
dinA[loop_var]=GAM;
addrA[loop_var]=count[3:0];
weA[loop_var]=1'b1;
end
end


`processing_state0: begin

for(loop_var=0;loop_var<768; loop_var=loop_var+1) begin
weA[loop_var]=1'b0;
weA1[loop_var]=1'b0;

end
for(row_state=0;row_state<256; row_state=row_state+1) begin
addrA[( col_row[row_state][0]*10'd2)+{9'd0,alphaCSR[row_state][ col_row[row_state][0]]}]=4'd0;
end

for(row_state=0;row_state<256; row_state=row_state+1) begin
addrA1[(col_row[row_state][2]*10'd2)+{9'd0,alphaCSR[row_state][col_row[row_state][2]]}]=4'd0;
end


end


`processing_state1: begin
for(loop_var=0;loop_var<768; loop_var=loop_var+1) begin
weA[loop_var]=1'b0;
weA1[loop_var]=1'b0;
end


for(row_state=0;row_state<256; row_state=row_state+1) begin

inv_gf(H[row_state][col_row[row_state][0]],inv_val[row_state]);
mul_gf(inv_val[row_state],a_read_FB[3:0],mul_val[row_state]);
addrA[( col_row[row_state][0]*10'd2)+{9'd0,alphaCSR[row_state][ col_row[row_state][0]]}]=mul_val[row_state];
end



for(row_state=0;row_state<256;row_state=row_state+1)
begin
inv_gf(H[row_state][col_row[row_state][2]],inv_val1[row_state]);
mul_gf(inv_val1[row_state],a_read_FB[3:0],mul_val1[row_state]);
addrA1[(col_row[row_state][2]*10'd2)+{9'd0,alphaCSR[row_state][col_row[row_state][2]]}]=mul_val1[row_state];
end





end



`FB_init1: begin

for(loop_var=0;loop_var<768; loop_var=loop_var+1) begin
weA[loop_var]=1'd0;
weA1[loop_var]=1'd0;
end


for(row_state=0;row_state<256; row_state=row_state+1) begin

inv_gf(H[row_state][col_row[row_state][0]],inv_val[row_state]);
mul_gf(inv_val[row_state],a_read_FB[3:0],mul_val[row_state]);
addrA[(col_row[row_state][0]*10'd2)+{9'd0,alphaCSR[row_state][ col_row[row_state][0]]}]=mul_val[row_state];
end



for(row_state=0;row_state<256;row_state=row_state+1)
begin
inv_gf(H[row_state][col_row[row_state][2]],inv_val1[row_state]);
mul_gf(inv_val1[row_state],a_read_FB[3:0],mul_val1[row_state]);
addrA1[(col_row[row_state][2]*10'd2)+{9'd0,alphaCSR[row_state][col_row[row_state][2]]}]=mul_val1[row_state];
end


for(row_state=0;row_state<256;row_state=row_state+1) begin
F[a_write_FB][0][row_state]=doutA[( col_row[row_state][0]*10'd2)+{9'd0,alphaCSR[row_state][ col_row[row_state][0]]}];

B[a_write_FB][2][row_state]=doutA1[(col_row[row_state][2]*10'd2)+{9'd0,alphaCSR[row_state][col_row[row_state][2]]}];
end



end


`F_OUT: begin
out_enable=1;
row_state={6'd0,f_count[11:8]};
col_state={2'd0,f_count[7:0]};

out=F[row_state][0][col_state];
end

`B_OUT: begin
row_state={6'd0,b_count[11:8]};
col_state={2'd0,b_count[7:0]};


out=B[row_state][2][col_state];

if(b_count!=12'b1111_1111_1111) begin
out_enable=1'b1;
end
else
out_enable=1'b0;
end

`END: begin
out_enable=1'b0;

end


default: begin


for(loop_var=0;loop_var<768;loop_var=loop_var+1) begin
addrA[loop_var]=addrA_[loop_var];
end
for(loop_var=0;loop_var<16;loop_var=loop_var+1) begin
for(loop_var1=0;loop_var1<3;loop_var1=loop_var1+1) begin
for(loop_var2=0;loop_var2<256;loop_var2=loop_var2+1) begin
F[loop_var][loop_var1][loop_var2]=F_[loop_var][loop_var1][loop_var2];
end
end
end
for(loop_var=0;loop_var<16;loop_var=loop_var+1) begin
for(loop_var1=0;loop_var1<3;loop_var1=loop_var1+1) begin
for(loop_var2=0;loop_var2<256;loop_var2=loop_var2+1) begin
B[loop_var][loop_var1][loop_var2]=B_[loop_var][loop_var1][loop_var2];
end
end
end


end
endcase
end

end



always@(posedge clk or posedge reset) begin
if(reset)
state=6'd0;
else
state=next_state;
end


always@(posedge clk,posedge reset) begin
if(reset)
begin
for(row2=0;row2<2;row2=row2+1) begin
for(col2=0;col2<384;col2=col2+1) begin
row_col[row2][col2]=0;
end
end
for(row2=0;row2<256;row2=row2+1) begin
for(col2=0;col2<384;col2=col2+1) begin
alphaCSR[row2][col2]=0;
H[row2][col2]=0;
end
end


for(row2=0;row2<256;row2=row2+1) begin
for(col2=0;col2<3;col2=col2+1) begin
col_row[row2][col2]=0;
end
end


end
else begin

alphaCSR[0][0]=0;
alphaCSR[127][0]=1;
alphaCSR[0][1]=0;
alphaCSR[1][1]=1;
alphaCSR[1][2]=0;
alphaCSR[2][2]=1;
alphaCSR[2][3]=0;
alphaCSR[3][3]=1;
alphaCSR[3][4]=0;
alphaCSR[4][4]=1;
alphaCSR[4][5]=0;
alphaCSR[5][5]=1;
alphaCSR[5][6]=0;
alphaCSR[6][6]=1;
alphaCSR[6][7]=0;
alphaCSR[7][7]=1;
alphaCSR[7][8]=0;
alphaCSR[8][8]=1;
alphaCSR[8][9]=0;
alphaCSR[9][9]=1;
alphaCSR[9][10]=0;
alphaCSR[10][10]=1;
alphaCSR[10][11]=0;
alphaCSR[11][11]=1;
alphaCSR[11][12]=0;
alphaCSR[12][12]=1;
alphaCSR[12][13]=0;
alphaCSR[13][13]=1;
alphaCSR[13][14]=0;
alphaCSR[14][14]=1;
alphaCSR[14][15]=0;
alphaCSR[15][15]=1;
alphaCSR[15][16]=0;
alphaCSR[16][16]=1;
alphaCSR[16][17]=0;
alphaCSR[17][17]=1;
alphaCSR[17][18]=0;
alphaCSR[18][18]=1;
alphaCSR[18][19]=0;
alphaCSR[19][19]=1;
alphaCSR[19][20]=0;
alphaCSR[20][20]=1;
alphaCSR[20][21]=0;
alphaCSR[21][21]=1;
alphaCSR[21][22]=0;
alphaCSR[22][22]=1;
alphaCSR[22][23]=0;
alphaCSR[23][23]=1;
alphaCSR[23][24]=0;
alphaCSR[24][24]=1;
alphaCSR[24][25]=0;
alphaCSR[25][25]=1;
alphaCSR[25][26]=0;
alphaCSR[26][26]=1;
alphaCSR[26][27]=0;
alphaCSR[27][27]=1;
alphaCSR[27][28]=0;
alphaCSR[28][28]=1;
alphaCSR[28][29]=0;
alphaCSR[29][29]=1;
alphaCSR[29][30]=0;
alphaCSR[30][30]=1;
alphaCSR[30][31]=0;
alphaCSR[31][31]=1;
alphaCSR[31][32]=0;
alphaCSR[32][32]=1;
alphaCSR[32][33]=0;
alphaCSR[33][33]=1;
alphaCSR[33][34]=0;
alphaCSR[34][34]=1;
alphaCSR[34][35]=0;
alphaCSR[35][35]=1;
alphaCSR[35][36]=0;
alphaCSR[36][36]=1;
alphaCSR[36][37]=0;
alphaCSR[37][37]=1;
alphaCSR[37][38]=0;
alphaCSR[38][38]=1;
alphaCSR[38][39]=0;
alphaCSR[39][39]=1;
alphaCSR[39][40]=0;
alphaCSR[40][40]=1;
alphaCSR[40][41]=0;
alphaCSR[41][41]=1;
alphaCSR[41][42]=0;
alphaCSR[42][42]=1;
alphaCSR[42][43]=0;
alphaCSR[43][43]=1;
alphaCSR[43][44]=0;
alphaCSR[44][44]=1;
alphaCSR[44][45]=0;
alphaCSR[45][45]=1;
alphaCSR[45][46]=0;
alphaCSR[46][46]=1;
alphaCSR[46][47]=0;
alphaCSR[47][47]=1;
alphaCSR[47][48]=0;
alphaCSR[48][48]=1;
alphaCSR[48][49]=0;
alphaCSR[49][49]=1;
alphaCSR[49][50]=0;
alphaCSR[50][50]=1;
alphaCSR[50][51]=0;
alphaCSR[51][51]=1;
alphaCSR[51][52]=0;
alphaCSR[52][52]=1;
alphaCSR[52][53]=0;
alphaCSR[53][53]=1;
alphaCSR[53][54]=0;
alphaCSR[54][54]=1;
alphaCSR[54][55]=0;
alphaCSR[55][55]=1;
alphaCSR[55][56]=0;
alphaCSR[56][56]=1;
alphaCSR[56][57]=0;
alphaCSR[57][57]=1;
alphaCSR[57][58]=0;
alphaCSR[58][58]=1;
alphaCSR[58][59]=0;
alphaCSR[59][59]=1;
alphaCSR[59][60]=0;
alphaCSR[60][60]=1;
alphaCSR[60][61]=0;
alphaCSR[61][61]=1;
alphaCSR[61][62]=0;
alphaCSR[62][62]=1;
alphaCSR[62][63]=0;
alphaCSR[63][63]=1;
alphaCSR[63][64]=0;
alphaCSR[64][64]=1;
alphaCSR[64][65]=0;
alphaCSR[65][65]=1;
alphaCSR[65][66]=0;
alphaCSR[66][66]=1;
alphaCSR[66][67]=0;
alphaCSR[67][67]=1;
alphaCSR[67][68]=0;
alphaCSR[68][68]=1;
alphaCSR[68][69]=0;
alphaCSR[69][69]=1;
alphaCSR[69][70]=0;
alphaCSR[70][70]=1;
alphaCSR[70][71]=0;
alphaCSR[71][71]=1;
alphaCSR[71][72]=0;
alphaCSR[72][72]=1;
alphaCSR[72][73]=0;
alphaCSR[73][73]=1;
alphaCSR[73][74]=0;
alphaCSR[74][74]=1;
alphaCSR[74][75]=0;
alphaCSR[75][75]=1;
alphaCSR[75][76]=0;
alphaCSR[76][76]=1;
alphaCSR[76][77]=0;
alphaCSR[77][77]=1;
alphaCSR[77][78]=0;
alphaCSR[78][78]=1;
alphaCSR[78][79]=0;
alphaCSR[79][79]=1;
alphaCSR[79][80]=0;
alphaCSR[80][80]=1;
alphaCSR[80][81]=0;
alphaCSR[81][81]=1;
alphaCSR[81][82]=0;
alphaCSR[82][82]=1;
alphaCSR[82][83]=0;
alphaCSR[83][83]=1;
alphaCSR[83][84]=0;
alphaCSR[84][84]=1;
alphaCSR[84][85]=0;
alphaCSR[85][85]=1;
alphaCSR[85][86]=0;
alphaCSR[86][86]=1;
alphaCSR[86][87]=0;
alphaCSR[87][87]=1;
alphaCSR[87][88]=0;
alphaCSR[88][88]=1;
alphaCSR[88][89]=0;
alphaCSR[89][89]=1;
alphaCSR[89][90]=0;
alphaCSR[90][90]=1;
alphaCSR[90][91]=0;
alphaCSR[91][91]=1;
alphaCSR[91][92]=0;
alphaCSR[92][92]=1;
alphaCSR[92][93]=0;
alphaCSR[93][93]=1;
alphaCSR[93][94]=0;
alphaCSR[94][94]=1;
alphaCSR[94][95]=0;
alphaCSR[95][95]=1;
alphaCSR[95][96]=0;
alphaCSR[96][96]=1;
alphaCSR[96][97]=0;
alphaCSR[97][97]=1;
alphaCSR[97][98]=0;
alphaCSR[98][98]=1;
alphaCSR[98][99]=0;
alphaCSR[99][99]=1;
alphaCSR[99][100]=0;
alphaCSR[100][100]=1;
alphaCSR[100][101]=0;
alphaCSR[101][101]=1;
alphaCSR[101][102]=0;
alphaCSR[102][102]=1;
alphaCSR[102][103]=0;
alphaCSR[103][103]=1;
alphaCSR[103][104]=0;
alphaCSR[104][104]=1;
alphaCSR[104][105]=0;
alphaCSR[105][105]=1;
alphaCSR[105][106]=0;
alphaCSR[106][106]=1;
alphaCSR[106][107]=0;
alphaCSR[107][107]=1;
alphaCSR[107][108]=0;
alphaCSR[108][108]=1;
alphaCSR[108][109]=0;
alphaCSR[109][109]=1;
alphaCSR[109][110]=0;
alphaCSR[110][110]=1;
alphaCSR[110][111]=0;
alphaCSR[111][111]=1;
alphaCSR[111][112]=0;
alphaCSR[112][112]=1;
alphaCSR[112][113]=0;
alphaCSR[113][113]=1;
alphaCSR[113][114]=0;
alphaCSR[114][114]=1;
alphaCSR[114][115]=0;
alphaCSR[115][115]=1;
alphaCSR[115][116]=0;
alphaCSR[116][116]=1;
alphaCSR[116][117]=0;
alphaCSR[117][117]=1;
alphaCSR[117][118]=0;
alphaCSR[118][118]=1;
alphaCSR[118][119]=0;
alphaCSR[119][119]=1;
alphaCSR[119][120]=0;
alphaCSR[120][120]=1;
alphaCSR[120][121]=0;
alphaCSR[121][121]=1;
alphaCSR[121][122]=0;
alphaCSR[122][122]=1;
alphaCSR[122][123]=0;
alphaCSR[123][123]=1;
alphaCSR[123][124]=0;
alphaCSR[124][124]=1;
alphaCSR[124][125]=0;
alphaCSR[125][125]=1;
alphaCSR[125][126]=0;
alphaCSR[126][126]=1;
alphaCSR[126][127]=0;
alphaCSR[127][127]=1;
alphaCSR[128][128]=0;
alphaCSR[255][128]=1;
alphaCSR[128][129]=0;
alphaCSR[129][129]=1;
alphaCSR[129][130]=0;
alphaCSR[130][130]=1;
alphaCSR[130][131]=0;
alphaCSR[131][131]=1;
alphaCSR[131][132]=0;
alphaCSR[132][132]=1;
alphaCSR[132][133]=0;
alphaCSR[133][133]=1;
alphaCSR[133][134]=0;
alphaCSR[134][134]=1;
alphaCSR[134][135]=0;
alphaCSR[135][135]=1;
alphaCSR[135][136]=0;
alphaCSR[136][136]=1;
alphaCSR[136][137]=0;
alphaCSR[137][137]=1;
alphaCSR[137][138]=0;
alphaCSR[138][138]=1;
alphaCSR[138][139]=0;
alphaCSR[139][139]=1;
alphaCSR[139][140]=0;
alphaCSR[140][140]=1;
alphaCSR[140][141]=0;
alphaCSR[141][141]=1;
alphaCSR[141][142]=0;
alphaCSR[142][142]=1;
alphaCSR[142][143]=0;
alphaCSR[143][143]=1;
alphaCSR[143][144]=0;
alphaCSR[144][144]=1;
alphaCSR[144][145]=0;
alphaCSR[145][145]=1;
alphaCSR[145][146]=0;
alphaCSR[146][146]=1;
alphaCSR[146][147]=0;
alphaCSR[147][147]=1;
alphaCSR[147][148]=0;
alphaCSR[148][148]=1;
alphaCSR[148][149]=0;
alphaCSR[149][149]=1;
alphaCSR[149][150]=0;
alphaCSR[150][150]=1;
alphaCSR[150][151]=0;
alphaCSR[151][151]=1;
alphaCSR[151][152]=0;
alphaCSR[152][152]=1;
alphaCSR[152][153]=0;
alphaCSR[153][153]=1;
alphaCSR[153][154]=0;
alphaCSR[154][154]=1;
alphaCSR[154][155]=0;
alphaCSR[155][155]=1;
alphaCSR[155][156]=0;
alphaCSR[156][156]=1;
alphaCSR[156][157]=0;
alphaCSR[157][157]=1;
alphaCSR[157][158]=0;
alphaCSR[158][158]=1;
alphaCSR[158][159]=0;
alphaCSR[159][159]=1;
alphaCSR[159][160]=0;
alphaCSR[160][160]=1;
alphaCSR[160][161]=0;
alphaCSR[161][161]=1;
alphaCSR[161][162]=0;
alphaCSR[162][162]=1;
alphaCSR[162][163]=0;
alphaCSR[163][163]=1;
alphaCSR[163][164]=0;
alphaCSR[164][164]=1;
alphaCSR[164][165]=0;
alphaCSR[165][165]=1;
alphaCSR[165][166]=0;
alphaCSR[166][166]=1;
alphaCSR[166][167]=0;
alphaCSR[167][167]=1;
alphaCSR[167][168]=0;
alphaCSR[168][168]=1;
alphaCSR[168][169]=0;
alphaCSR[169][169]=1;
alphaCSR[169][170]=0;
alphaCSR[170][170]=1;
alphaCSR[170][171]=0;
alphaCSR[171][171]=1;
alphaCSR[171][172]=0;
alphaCSR[172][172]=1;
alphaCSR[172][173]=0;
alphaCSR[173][173]=1;
alphaCSR[173][174]=0;
alphaCSR[174][174]=1;
alphaCSR[174][175]=0;
alphaCSR[175][175]=1;
alphaCSR[175][176]=0;
alphaCSR[176][176]=1;
alphaCSR[176][177]=0;
alphaCSR[177][177]=1;
alphaCSR[177][178]=0;
alphaCSR[178][178]=1;
alphaCSR[178][179]=0;
alphaCSR[179][179]=1;
alphaCSR[179][180]=0;
alphaCSR[180][180]=1;
alphaCSR[180][181]=0;
alphaCSR[181][181]=1;
alphaCSR[181][182]=0;
alphaCSR[182][182]=1;
alphaCSR[182][183]=0;
alphaCSR[183][183]=1;
alphaCSR[183][184]=0;
alphaCSR[184][184]=1;
alphaCSR[184][185]=0;
alphaCSR[185][185]=1;
alphaCSR[185][186]=0;
alphaCSR[186][186]=1;
alphaCSR[186][187]=0;
alphaCSR[187][187]=1;
alphaCSR[187][188]=0;
alphaCSR[188][188]=1;
alphaCSR[188][189]=0;
alphaCSR[189][189]=1;
alphaCSR[189][190]=0;
alphaCSR[190][190]=1;
alphaCSR[190][191]=0;
alphaCSR[191][191]=1;
alphaCSR[191][192]=0;
alphaCSR[192][192]=1;
alphaCSR[192][193]=0;
alphaCSR[193][193]=1;
alphaCSR[193][194]=0;
alphaCSR[194][194]=1;
alphaCSR[194][195]=0;
alphaCSR[195][195]=1;
alphaCSR[195][196]=0;
alphaCSR[196][196]=1;
alphaCSR[196][197]=0;
alphaCSR[197][197]=1;
alphaCSR[197][198]=0;
alphaCSR[198][198]=1;
alphaCSR[198][199]=0;
alphaCSR[199][199]=1;
alphaCSR[199][200]=0;
alphaCSR[200][200]=1;
alphaCSR[200][201]=0;
alphaCSR[201][201]=1;
alphaCSR[201][202]=0;
alphaCSR[202][202]=1;
alphaCSR[202][203]=0;
alphaCSR[203][203]=1;
alphaCSR[203][204]=0;
alphaCSR[204][204]=1;
alphaCSR[204][205]=0;
alphaCSR[205][205]=1;
alphaCSR[205][206]=0;
alphaCSR[206][206]=1;
alphaCSR[206][207]=0;
alphaCSR[207][207]=1;
alphaCSR[207][208]=0;
alphaCSR[208][208]=1;
alphaCSR[208][209]=0;
alphaCSR[209][209]=1;
alphaCSR[209][210]=0;
alphaCSR[210][210]=1;
alphaCSR[210][211]=0;
alphaCSR[211][211]=1;
alphaCSR[211][212]=0;
alphaCSR[212][212]=1;
alphaCSR[212][213]=0;
alphaCSR[213][213]=1;
alphaCSR[213][214]=0;
alphaCSR[214][214]=1;
alphaCSR[214][215]=0;
alphaCSR[215][215]=1;
alphaCSR[215][216]=0;
alphaCSR[216][216]=1;
alphaCSR[216][217]=0;
alphaCSR[217][217]=1;
alphaCSR[217][218]=0;
alphaCSR[218][218]=1;
alphaCSR[218][219]=0;
alphaCSR[219][219]=1;
alphaCSR[219][220]=0;
alphaCSR[220][220]=1;
alphaCSR[220][221]=0;
alphaCSR[221][221]=1;
alphaCSR[221][222]=0;
alphaCSR[222][222]=1;
alphaCSR[222][223]=0;
alphaCSR[223][223]=1;
alphaCSR[223][224]=0;
alphaCSR[224][224]=1;
alphaCSR[224][225]=0;
alphaCSR[225][225]=1;
alphaCSR[225][226]=0;
alphaCSR[226][226]=1;
alphaCSR[226][227]=0;
alphaCSR[227][227]=1;
alphaCSR[227][228]=0;
alphaCSR[228][228]=1;
alphaCSR[228][229]=0;
alphaCSR[229][229]=1;
alphaCSR[229][230]=0;
alphaCSR[230][230]=1;
alphaCSR[230][231]=0;
alphaCSR[231][231]=1;
alphaCSR[231][232]=0;
alphaCSR[232][232]=1;
alphaCSR[232][233]=0;
alphaCSR[233][233]=1;
alphaCSR[233][234]=0;
alphaCSR[234][234]=1;
alphaCSR[234][235]=0;
alphaCSR[235][235]=1;
alphaCSR[235][236]=0;
alphaCSR[236][236]=1;
alphaCSR[236][237]=0;
alphaCSR[237][237]=1;
alphaCSR[237][238]=0;
alphaCSR[238][238]=1;
alphaCSR[238][239]=0;
alphaCSR[239][239]=1;
alphaCSR[239][240]=0;
alphaCSR[240][240]=1;
alphaCSR[240][241]=0;
alphaCSR[241][241]=1;
alphaCSR[241][242]=0;
alphaCSR[242][242]=1;
alphaCSR[242][243]=0;
alphaCSR[243][243]=1;
alphaCSR[243][244]=0;
alphaCSR[244][244]=1;
alphaCSR[244][245]=0;
alphaCSR[245][245]=1;
alphaCSR[245][246]=0;
alphaCSR[246][246]=1;
alphaCSR[246][247]=0;
alphaCSR[247][247]=1;
alphaCSR[247][248]=0;
alphaCSR[248][248]=1;
alphaCSR[248][249]=0;
alphaCSR[249][249]=1;
alphaCSR[249][250]=0;
alphaCSR[250][250]=1;
alphaCSR[250][251]=0;
alphaCSR[251][251]=1;
alphaCSR[251][252]=0;
alphaCSR[252][252]=1;
alphaCSR[252][253]=0;
alphaCSR[253][253]=1;
alphaCSR[253][254]=0;
alphaCSR[254][254]=1;
alphaCSR[254][255]=0;
alphaCSR[255][255]=1;
alphaCSR[0][256]=0;
alphaCSR[141][256]=1;
alphaCSR[1][257]=0;
alphaCSR[132][257]=1;
alphaCSR[2][258]=0;
alphaCSR[251][258]=1;
alphaCSR[3][259]=0;
alphaCSR[148][259]=1;
alphaCSR[4][260]=0;
alphaCSR[243][260]=1;
alphaCSR[5][261]=0;
alphaCSR[156][261]=1;
alphaCSR[6][262]=0;
alphaCSR[165][262]=1;
alphaCSR[7][263]=0;
alphaCSR[236][263]=1;
alphaCSR[8][264]=0;
alphaCSR[135][264]=1;
alphaCSR[9][265]=0;
alphaCSR[172][265]=1;
alphaCSR[10][266]=0;
alphaCSR[145][266]=1;
alphaCSR[11][267]=0;
alphaCSR[246][267]=1;
alphaCSR[12][268]=0;
alphaCSR[129][268]=1;
alphaCSR[13][269]=0;
alphaCSR[152][269]=1;
alphaCSR[14][270]=0;
alphaCSR[177][270]=1;
alphaCSR[15][271]=0;
alphaCSR[238][271]=1;
alphaCSR[16][272]=0;
alphaCSR[159][272]=1;
alphaCSR[17][273]=0;
alphaCSR[184][273]=1;
alphaCSR[18][274]=0;
alphaCSR[231][274]=1;
alphaCSR[19][275]=0;
alphaCSR[254][275]=1;
alphaCSR[20][276]=0;
alphaCSR[223][276]=1;
alphaCSR[21][277]=0;
alphaCSR[142][277]=1;
alphaCSR[22][278]=0;
alphaCSR[153][278]=1;
alphaCSR[23][279]=0;
alphaCSR[170][279]=1;
alphaCSR[24][280]=0;
alphaCSR[187][280]=1;
alphaCSR[25][281]=0;
alphaCSR[242][281]=1;
alphaCSR[26][282]=0;
alphaCSR[195][282]=1;
alphaCSR[27][283]=0;
alphaCSR[230][283]=1;
alphaCSR[28][284]=0;
alphaCSR[219][284]=1;
alphaCSR[29][285]=0;
alphaCSR[174][285]=1;
alphaCSR[30][286]=0;
alphaCSR[211][286]=1;
alphaCSR[31][287]=0;
alphaCSR[200][287]=1;
alphaCSR[32][288]=0;
alphaCSR[167][288]=1;
alphaCSR[33][289]=0;
alphaCSR[138][289]=1;
alphaCSR[34][290]=0;
alphaCSR[247][290]=1;
alphaCSR[35][291]=0;
alphaCSR[228][291]=1;
alphaCSR[36][292]=0;
alphaCSR[189][292]=1;
alphaCSR[37][293]=0;
alphaCSR[150][293]=1;
alphaCSR[38][294]=0;
alphaCSR[163][294]=1;
alphaCSR[39][295]=0;
alphaCSR[198][295]=1;
alphaCSR[40][296]=0;
alphaCSR[217][296]=1;
alphaCSR[41][297]=0;
alphaCSR[134][297]=1;
alphaCSR[42][298]=0;
alphaCSR[209][298]=1;
alphaCSR[43][299]=0;
alphaCSR[186][299]=1;
alphaCSR[44][300]=0;
alphaCSR[147][300]=1;
alphaCSR[45][301]=0;
alphaCSR[224][301]=1;
alphaCSR[46][302]=0;
alphaCSR[175][302]=1;
alphaCSR[47][303]=0;
alphaCSR[248][303]=1;
alphaCSR[48][304]=0;
alphaCSR[205][304]=1;
alphaCSR[49][305]=0;
alphaCSR[158][305]=1;
alphaCSR[50][306]=0;
alphaCSR[197][306]=1;
alphaCSR[51][307]=0;
alphaCSR[144][307]=1;
alphaCSR[52][308]=0;
alphaCSR[181][308]=1;
alphaCSR[53][309]=0;
alphaCSR[214][309]=1;
alphaCSR[54][310]=0;
alphaCSR[239][310]=1;
alphaCSR[55][311]=0;
alphaCSR[190][311]=1;
alphaCSR[56][312]=0;
alphaCSR[253][312]=1;
alphaCSR[57][313]=0;
alphaCSR[208][313]=1;
alphaCSR[58][314]=0;
alphaCSR[139][314]=1;
alphaCSR[59][315]=0;
alphaCSR[162][315]=1;
alphaCSR[60][316]=0;
alphaCSR[225][316]=1;
alphaCSR[61][317]=0;
alphaCSR[244][317]=1;
alphaCSR[62][318]=0;
alphaCSR[203][318]=1;
alphaCSR[63][319]=0;
alphaCSR[178][319]=1;
alphaCSR[64][320]=0;
alphaCSR[133][320]=1;
alphaCSR[65][321]=0;
alphaCSR[194][321]=1;
alphaCSR[66][322]=0;
alphaCSR[155][322]=1;
alphaCSR[67][323]=0;
alphaCSR[212][323]=1;
alphaCSR[68][324]=0;
alphaCSR[255][324]=1;
alphaCSR[69][325]=0;
alphaCSR[149][325]=1;
alphaCSR[70][326]=0;
alphaCSR[136][326]=1;
alphaCSR[71][327]=0;
alphaCSR[183][327]=1;
alphaCSR[72][328]=0;
alphaCSR[221][328]=1;
alphaCSR[73][329]=0;
alphaCSR[250][329]=1;
alphaCSR[74][330]=0;
alphaCSR[168][330]=1;
alphaCSR[75][331]=0;
alphaCSR[215][331]=1;
alphaCSR[76][332]=0;
alphaCSR[226][332]=1;
alphaCSR[77][333]=0;
alphaCSR[234][333]=1;
alphaCSR[78][334]=0;
alphaCSR[128][334]=1;
alphaCSR[79][335]=0;
alphaCSR[196][335]=1;
alphaCSR[80][336]=0;
alphaCSR[140][336]=1;
alphaCSR[81][337]=0;
alphaCSR[173][337]=1;
alphaCSR[82][338]=0;
alphaCSR[182][338]=1;
alphaCSR[83][339]=0;
alphaCSR[154][339]=1;
alphaCSR[84][340]=0;
alphaCSR[202][340]=1;
alphaCSR[85][341]=0;
alphaCSR[191][341]=1;
alphaCSR[86][342]=0;
alphaCSR[131][342]=1;
alphaCSR[87][343]=0;
alphaCSR[169][343]=1;
alphaCSR[88][344]=0;
alphaCSR[161][344]=1;
alphaCSR[89][345]=0;
alphaCSR[180][345]=1;
alphaCSR[90][346]=0;
alphaCSR[232][346]=1;
alphaCSR[91][347]=0;
alphaCSR[245][347]=1;
alphaCSR[92][348]=0;
alphaCSR[216][348]=1;
alphaCSR[93][349]=0;
alphaCSR[192][349]=1;
alphaCSR[94][350]=0;
alphaCSR[143][350]=1;
alphaCSR[95][351]=0;
alphaCSR[164][351]=1;
alphaCSR[96][352]=0;
alphaCSR[252][352]=1;
alphaCSR[97][353]=0;
alphaCSR[176][353]=1;
alphaCSR[98][354]=0;
alphaCSR[233][354]=1;
alphaCSR[99][355]=0;
alphaCSR[137][355]=1;
alphaCSR[100][356]=0;
alphaCSR[157][356]=1;
alphaCSR[101][357]=0;
alphaCSR[188][357]=1;
alphaCSR[102][358]=0;
alphaCSR[220][358]=1;
alphaCSR[103][359]=0;
alphaCSR[130][359]=1;
alphaCSR[104][360]=0;
alphaCSR[206][360]=1;
alphaCSR[105][361]=0;
alphaCSR[237][361]=1;
alphaCSR[106][362]=0;
alphaCSR[229][362]=1;
alphaCSR[107][363]=0;
alphaCSR[146][363]=1;
alphaCSR[108][364]=0;
alphaCSR[201][364]=1;
alphaCSR[109][365]=0;
alphaCSR[249][365]=1;
alphaCSR[110][366]=0;
alphaCSR[241][366]=1;
alphaCSR[111][367]=0;
alphaCSR[151][367]=1;
alphaCSR[112][368]=0;
alphaCSR[210][368]=1;
alphaCSR[113][369]=0;
alphaCSR[235][369]=1;
alphaCSR[114][370]=0;
alphaCSR[193][370]=1;
alphaCSR[115][371]=0;
alphaCSR[160][371]=1;
alphaCSR[116][372]=0;
alphaCSR[222][372]=1;
alphaCSR[117][373]=0;
alphaCSR[199][373]=1;
alphaCSR[118][374]=0;
alphaCSR[171][374]=1;
alphaCSR[119][375]=0;
alphaCSR[207][375]=1;
alphaCSR[120][376]=0;
alphaCSR[179][376]=1;
alphaCSR[121][377]=0;
alphaCSR[218][377]=1;
alphaCSR[122][378]=0;
alphaCSR[166][378]=1;
alphaCSR[123][379]=0;
alphaCSR[240][379]=1;
alphaCSR[124][380]=0;
alphaCSR[227][380]=1;
alphaCSR[125][381]=0;
alphaCSR[185][381]=1;
alphaCSR[126][382]=0;
alphaCSR[204][382]=1;
alphaCSR[127][383]=0;
alphaCSR[213][383]=1;
//*/


row_col[0][0]=0;
row_col[1][0]=127;
row_col[0][1]=0;
row_col[1][1]=1;
row_col[0][2]=1;
row_col[1][2]=2;
row_col[0][3]=2;
row_col[1][3]=3;
row_col[0][4]=3;
row_col[1][4]=4;
row_col[0][5]=4;
row_col[1][5]=5;
row_col[0][6]=5;
row_col[1][6]=6;
row_col[0][7]=6;
row_col[1][7]=7;
row_col[0][8]=7;
row_col[1][8]=8;
row_col[0][9]=8;
row_col[1][9]=9;
row_col[0][10]=9;
row_col[1][10]=10;
row_col[0][11]=10;
row_col[1][11]=11;
row_col[0][12]=11;
row_col[1][12]=12;
row_col[0][13]=12;
row_col[1][13]=13;
row_col[0][14]=13;
row_col[1][14]=14;
row_col[0][15]=14;
row_col[1][15]=15;
row_col[0][16]=15;
row_col[1][16]=16;
row_col[0][17]=16;
row_col[1][17]=17;
row_col[0][18]=17;
row_col[1][18]=18;
row_col[0][19]=18;
row_col[1][19]=19;
row_col[0][20]=19;
row_col[1][20]=20;
row_col[0][21]=20;
row_col[1][21]=21;
row_col[0][22]=21;
row_col[1][22]=22;
row_col[0][23]=22;
row_col[1][23]=23;
row_col[0][24]=23;
row_col[1][24]=24;
row_col[0][25]=24;
row_col[1][25]=25;
row_col[0][26]=25;
row_col[1][26]=26;
row_col[0][27]=26;
row_col[1][27]=27;
row_col[0][28]=27;
row_col[1][28]=28;
row_col[0][29]=28;
row_col[1][29]=29;
row_col[0][30]=29;
row_col[1][30]=30;
row_col[0][31]=30;
row_col[1][31]=31;
row_col[0][32]=31;
row_col[1][32]=32;
row_col[0][33]=32;
row_col[1][33]=33;
row_col[0][34]=33;
row_col[1][34]=34;
row_col[0][35]=34;
row_col[1][35]=35;
row_col[0][36]=35;
row_col[1][36]=36;
row_col[0][37]=36;
row_col[1][37]=37;
row_col[0][38]=37;
row_col[1][38]=38;
row_col[0][39]=38;
row_col[1][39]=39;
row_col[0][40]=39;
row_col[1][40]=40;
row_col[0][41]=40;
row_col[1][41]=41;
row_col[0][42]=41;
row_col[1][42]=42;
row_col[0][43]=42;
row_col[1][43]=43;
row_col[0][44]=43;
row_col[1][44]=44;
row_col[0][45]=44;
row_col[1][45]=45;
row_col[0][46]=45;
row_col[1][46]=46;
row_col[0][47]=46;
row_col[1][47]=47;
row_col[0][48]=47;
row_col[1][48]=48;
row_col[0][49]=48;
row_col[1][49]=49;
row_col[0][50]=49;
row_col[1][50]=50;
row_col[0][51]=50;
row_col[1][51]=51;
row_col[0][52]=51;
row_col[1][52]=52;
row_col[0][53]=52;
row_col[1][53]=53;
row_col[0][54]=53;
row_col[1][54]=54;
row_col[0][55]=54;
row_col[1][55]=55;
row_col[0][56]=55;
row_col[1][56]=56;
row_col[0][57]=56;
row_col[1][57]=57;
row_col[0][58]=57;
row_col[1][58]=58;
row_col[0][59]=58;
row_col[1][59]=59;
row_col[0][60]=59;
row_col[1][60]=60;
row_col[0][61]=60;
row_col[1][61]=61;
row_col[0][62]=61;
row_col[1][62]=62;
row_col[0][63]=62;
row_col[1][63]=63;
row_col[0][64]=63;
row_col[1][64]=64;
row_col[0][65]=64;
row_col[1][65]=65;
row_col[0][66]=65;
row_col[1][66]=66;
row_col[0][67]=66;
row_col[1][67]=67;
row_col[0][68]=67;
row_col[1][68]=68;
row_col[0][69]=68;
row_col[1][69]=69;
row_col[0][70]=69;
row_col[1][70]=70;
row_col[0][71]=70;
row_col[1][71]=71;
row_col[0][72]=71;
row_col[1][72]=72;
row_col[0][73]=72;
row_col[1][73]=73;
row_col[0][74]=73;
row_col[1][74]=74;
row_col[0][75]=74;
row_col[1][75]=75;
row_col[0][76]=75;
row_col[1][76]=76;
row_col[0][77]=76;
row_col[1][77]=77;
row_col[0][78]=77;
row_col[1][78]=78;
row_col[0][79]=78;
row_col[1][79]=79;
row_col[0][80]=79;
row_col[1][80]=80;
row_col[0][81]=80;
row_col[1][81]=81;
row_col[0][82]=81;
row_col[1][82]=82;
row_col[0][83]=82;
row_col[1][83]=83;
row_col[0][84]=83;
row_col[1][84]=84;
row_col[0][85]=84;
row_col[1][85]=85;
row_col[0][86]=85;
row_col[1][86]=86;
row_col[0][87]=86;
row_col[1][87]=87;
row_col[0][88]=87;
row_col[1][88]=88;
row_col[0][89]=88;
row_col[1][89]=89;
row_col[0][90]=89;
row_col[1][90]=90;
row_col[0][91]=90;
row_col[1][91]=91;
row_col[0][92]=91;
row_col[1][92]=92;
row_col[0][93]=92;
row_col[1][93]=93;
row_col[0][94]=93;
row_col[1][94]=94;
row_col[0][95]=94;
row_col[1][95]=95;
row_col[0][96]=95;
row_col[1][96]=96;
row_col[0][97]=96;
row_col[1][97]=97;
row_col[0][98]=97;
row_col[1][98]=98;
row_col[0][99]=98;
row_col[1][99]=99;
row_col[0][100]=99;
row_col[1][100]=100;
row_col[0][101]=100;
row_col[1][101]=101;
row_col[0][102]=101;
row_col[1][102]=102;
row_col[0][103]=102;
row_col[1][103]=103;
row_col[0][104]=103;
row_col[1][104]=104;
row_col[0][105]=104;
row_col[1][105]=105;
row_col[0][106]=105;
row_col[1][106]=106;
row_col[0][107]=106;
row_col[1][107]=107;
row_col[0][108]=107;
row_col[1][108]=108;
row_col[0][109]=108;
row_col[1][109]=109;
row_col[0][110]=109;
row_col[1][110]=110;
row_col[0][111]=110;
row_col[1][111]=111;
row_col[0][112]=111;
row_col[1][112]=112;
row_col[0][113]=112;
row_col[1][113]=113;
row_col[0][114]=113;
row_col[1][114]=114;
row_col[0][115]=114;
row_col[1][115]=115;
row_col[0][116]=115;
row_col[1][116]=116;
row_col[0][117]=116;
row_col[1][117]=117;
row_col[0][118]=117;
row_col[1][118]=118;
row_col[0][119]=118;
row_col[1][119]=119;
row_col[0][120]=119;
row_col[1][120]=120;
row_col[0][121]=120;
row_col[1][121]=121;
row_col[0][122]=121;
row_col[1][122]=122;
row_col[0][123]=122;
row_col[1][123]=123;
row_col[0][124]=123;
row_col[1][124]=124;
row_col[0][125]=124;
row_col[1][125]=125;
row_col[0][126]=125;
row_col[1][126]=126;
row_col[0][127]=126;
row_col[1][127]=127;
row_col[0][128]=128;
row_col[1][128]=255;
row_col[0][129]=128;
row_col[1][129]=129;
row_col[0][130]=129;
row_col[1][130]=130;
row_col[0][131]=130;
row_col[1][131]=131;
row_col[0][132]=131;
row_col[1][132]=132;
row_col[0][133]=132;
row_col[1][133]=133;
row_col[0][134]=133;
row_col[1][134]=134;
row_col[0][135]=134;
row_col[1][135]=135;
row_col[0][136]=135;
row_col[1][136]=136;
row_col[0][137]=136;
row_col[1][137]=137;
row_col[0][138]=137;
row_col[1][138]=138;
row_col[0][139]=138;
row_col[1][139]=139;
row_col[0][140]=139;
row_col[1][140]=140;
row_col[0][141]=140;
row_col[1][141]=141;
row_col[0][142]=141;
row_col[1][142]=142;
row_col[0][143]=142;
row_col[1][143]=143;
row_col[0][144]=143;
row_col[1][144]=144;
row_col[0][145]=144;
row_col[1][145]=145;
row_col[0][146]=145;
row_col[1][146]=146;
row_col[0][147]=146;
row_col[1][147]=147;
row_col[0][148]=147;
row_col[1][148]=148;
row_col[0][149]=148;
row_col[1][149]=149;
row_col[0][150]=149;
row_col[1][150]=150;
row_col[0][151]=150;
row_col[1][151]=151;
row_col[0][152]=151;
row_col[1][152]=152;
row_col[0][153]=152;
row_col[1][153]=153;
row_col[0][154]=153;
row_col[1][154]=154;
row_col[0][155]=154;
row_col[1][155]=155;
row_col[0][156]=155;
row_col[1][156]=156;
row_col[0][157]=156;
row_col[1][157]=157;
row_col[0][158]=157;
row_col[1][158]=158;
row_col[0][159]=158;
row_col[1][159]=159;
row_col[0][160]=159;
row_col[1][160]=160;
row_col[0][161]=160;
row_col[1][161]=161;
row_col[0][162]=161;
row_col[1][162]=162;
row_col[0][163]=162;
row_col[1][163]=163;
row_col[0][164]=163;
row_col[1][164]=164;
row_col[0][165]=164;
row_col[1][165]=165;
row_col[0][166]=165;
row_col[1][166]=166;
row_col[0][167]=166;
row_col[1][167]=167;
row_col[0][168]=167;
row_col[1][168]=168;
row_col[0][169]=168;
row_col[1][169]=169;
row_col[0][170]=169;
row_col[1][170]=170;
row_col[0][171]=170;
row_col[1][171]=171;
row_col[0][172]=171;
row_col[1][172]=172;
row_col[0][173]=172;
row_col[1][173]=173;
row_col[0][174]=173;
row_col[1][174]=174;
row_col[0][175]=174;
row_col[1][175]=175;
row_col[0][176]=175;
row_col[1][176]=176;
row_col[0][177]=176;
row_col[1][177]=177;
row_col[0][178]=177;
row_col[1][178]=178;
row_col[0][179]=178;
row_col[1][179]=179;
row_col[0][180]=179;
row_col[1][180]=180;
row_col[0][181]=180;
row_col[1][181]=181;
row_col[0][182]=181;
row_col[1][182]=182;
row_col[0][183]=182;
row_col[1][183]=183;
row_col[0][184]=183;
row_col[1][184]=184;
row_col[0][185]=184;
row_col[1][185]=185;
row_col[0][186]=185;
row_col[1][186]=186;
row_col[0][187]=186;
row_col[1][187]=187;
row_col[0][188]=187;
row_col[1][188]=188;
row_col[0][189]=188;
row_col[1][189]=189;
row_col[0][190]=189;
row_col[1][190]=190;
row_col[0][191]=190;
row_col[1][191]=191;
row_col[0][192]=191;
row_col[1][192]=192;
row_col[0][193]=192;
row_col[1][193]=193;
row_col[0][194]=193;
row_col[1][194]=194;
row_col[0][195]=194;
row_col[1][195]=195;
row_col[0][196]=195;
row_col[1][196]=196;
row_col[0][197]=196;
row_col[1][197]=197;
row_col[0][198]=197;
row_col[1][198]=198;
row_col[0][199]=198;
row_col[1][199]=199;
row_col[0][200]=199;
row_col[1][200]=200;
row_col[0][201]=200;
row_col[1][201]=201;
row_col[0][202]=201;
row_col[1][202]=202;
row_col[0][203]=202;
row_col[1][203]=203;
row_col[0][204]=203;
row_col[1][204]=204;
row_col[0][205]=204;
row_col[1][205]=205;
row_col[0][206]=205;
row_col[1][206]=206;
row_col[0][207]=206;
row_col[1][207]=207;
row_col[0][208]=207;
row_col[1][208]=208;
row_col[0][209]=208;
row_col[1][209]=209;
row_col[0][210]=209;
row_col[1][210]=210;
row_col[0][211]=210;
row_col[1][211]=211;
row_col[0][212]=211;
row_col[1][212]=212;
row_col[0][213]=212;
row_col[1][213]=213;
row_col[0][214]=213;
row_col[1][214]=214;
row_col[0][215]=214;
row_col[1][215]=215;
row_col[0][216]=215;
row_col[1][216]=216;
row_col[0][217]=216;
row_col[1][217]=217;
row_col[0][218]=217;
row_col[1][218]=218;
row_col[0][219]=218;
row_col[1][219]=219;
row_col[0][220]=219;
row_col[1][220]=220;
row_col[0][221]=220;
row_col[1][221]=221;
row_col[0][222]=221;
row_col[1][222]=222;
row_col[0][223]=222;
row_col[1][223]=223;
row_col[0][224]=223;
row_col[1][224]=224;
row_col[0][225]=224;
row_col[1][225]=225;
row_col[0][226]=225;
row_col[1][226]=226;
row_col[0][227]=226;
row_col[1][227]=227;
row_col[0][228]=227;
row_col[1][228]=228;
row_col[0][229]=228;
row_col[1][229]=229;
row_col[0][230]=229;
row_col[1][230]=230;
row_col[0][231]=230;
row_col[1][231]=231;
row_col[0][232]=231;
row_col[1][232]=232;
row_col[0][233]=232;
row_col[1][233]=233;
row_col[0][234]=233;
row_col[1][234]=234;
row_col[0][235]=234;
row_col[1][235]=235;
row_col[0][236]=235;
row_col[1][236]=236;
row_col[0][237]=236;
row_col[1][237]=237;
row_col[0][238]=237;
row_col[1][238]=238;
row_col[0][239]=238;
row_col[1][239]=239;
row_col[0][240]=239;
row_col[1][240]=240;
row_col[0][241]=240;
row_col[1][241]=241;
row_col[0][242]=241;
row_col[1][242]=242;
row_col[0][243]=242;
row_col[1][243]=243;
row_col[0][244]=243;
row_col[1][244]=244;
row_col[0][245]=244;
row_col[1][245]=245;
row_col[0][246]=245;
row_col[1][246]=246;
row_col[0][247]=246;
row_col[1][247]=247;
row_col[0][248]=247;
row_col[1][248]=248;
row_col[0][249]=248;
row_col[1][249]=249;
row_col[0][250]=249;
row_col[1][250]=250;
row_col[0][251]=250;
row_col[1][251]=251;
row_col[0][252]=251;
row_col[1][252]=252;
row_col[0][253]=252;
row_col[1][253]=253;
row_col[0][254]=253;
row_col[1][254]=254;
row_col[0][255]=254;
row_col[1][255]=255;
row_col[0][256]=0;
row_col[1][256]=141;
row_col[0][257]=1;
row_col[1][257]=132;
row_col[0][258]=2;
row_col[1][258]=251;
row_col[0][259]=3;
row_col[1][259]=148;
row_col[0][260]=4;
row_col[1][260]=243;
row_col[0][261]=5;
row_col[1][261]=156;
row_col[0][262]=6;
row_col[1][262]=165;
row_col[0][263]=7;
row_col[1][263]=236;
row_col[0][264]=8;
row_col[1][264]=135;
row_col[0][265]=9;
row_col[1][265]=172;
row_col[0][266]=10;
row_col[1][266]=145;
row_col[0][267]=11;
row_col[1][267]=246;
row_col[0][268]=12;
row_col[1][268]=129;
row_col[0][269]=13;
row_col[1][269]=152;
row_col[0][270]=14;
row_col[1][270]=177;
row_col[0][271]=15;
row_col[1][271]=238;
row_col[0][272]=16;
row_col[1][272]=159;
row_col[0][273]=17;
row_col[1][273]=184;
row_col[0][274]=18;
row_col[1][274]=231;
row_col[0][275]=19;
row_col[1][275]=254;
row_col[0][276]=20;
row_col[1][276]=223;
row_col[0][277]=21;
row_col[1][277]=142;
row_col[0][278]=22;
row_col[1][278]=153;
row_col[0][279]=23;
row_col[1][279]=170;
row_col[0][280]=24;
row_col[1][280]=187;
row_col[0][281]=25;
row_col[1][281]=242;
row_col[0][282]=26;
row_col[1][282]=195;
row_col[0][283]=27;
row_col[1][283]=230;
row_col[0][284]=28;
row_col[1][284]=219;
row_col[0][285]=29;
row_col[1][285]=174;
row_col[0][286]=30;
row_col[1][286]=211;
row_col[0][287]=31;
row_col[1][287]=200;
row_col[0][288]=32;
row_col[1][288]=167;
row_col[0][289]=33;
row_col[1][289]=138;
row_col[0][290]=34;
row_col[1][290]=247;
row_col[0][291]=35;
row_col[1][291]=228;
row_col[0][292]=36;
row_col[1][292]=189;
row_col[0][293]=37;
row_col[1][293]=150;
row_col[0][294]=38;
row_col[1][294]=163;
row_col[0][295]=39;
row_col[1][295]=198;
row_col[0][296]=40;
row_col[1][296]=217;
row_col[0][297]=41;
row_col[1][297]=134;
row_col[0][298]=42;
row_col[1][298]=209;
row_col[0][299]=43;
row_col[1][299]=186;
row_col[0][300]=44;
row_col[1][300]=147;
row_col[0][301]=45;
row_col[1][301]=224;
row_col[0][302]=46;
row_col[1][302]=175;
row_col[0][303]=47;
row_col[1][303]=248;
row_col[0][304]=48;
row_col[1][304]=205;
row_col[0][305]=49;
row_col[1][305]=158;
row_col[0][306]=50;
row_col[1][306]=197;
row_col[0][307]=51;
row_col[1][307]=144;
row_col[0][308]=52;
row_col[1][308]=181;
row_col[0][309]=53;
row_col[1][309]=214;
row_col[0][310]=54;
row_col[1][310]=239;
row_col[0][311]=55;
row_col[1][311]=190;
row_col[0][312]=56;
row_col[1][312]=253;
row_col[0][313]=57;
row_col[1][313]=208;
row_col[0][314]=58;
row_col[1][314]=139;
row_col[0][315]=59;
row_col[1][315]=162;
row_col[0][316]=60;
row_col[1][316]=225;
row_col[0][317]=61;
row_col[1][317]=244;
row_col[0][318]=62;
row_col[1][318]=203;
row_col[0][319]=63;
row_col[1][319]=178;
row_col[0][320]=64;
row_col[1][320]=133;
row_col[0][321]=65;
row_col[1][321]=194;
row_col[0][322]=66;
row_col[1][322]=155;
row_col[0][323]=67;
row_col[1][323]=212;
row_col[0][324]=68;
row_col[1][324]=255;
row_col[0][325]=69;
row_col[1][325]=149;
row_col[0][326]=70;
row_col[1][326]=136;
row_col[0][327]=71;
row_col[1][327]=183;
row_col[0][328]=72;
row_col[1][328]=221;
row_col[0][329]=73;
row_col[1][329]=250;
row_col[0][330]=74;
row_col[1][330]=168;
row_col[0][331]=75;
row_col[1][331]=215;
row_col[0][332]=76;
row_col[1][332]=226;
row_col[0][333]=77;
row_col[1][333]=234;
row_col[0][334]=78;
row_col[1][334]=128;
row_col[0][335]=79;
row_col[1][335]=196;
row_col[0][336]=80;
row_col[1][336]=140;
row_col[0][337]=81;
row_col[1][337]=173;
row_col[0][338]=82;
row_col[1][338]=182;
row_col[0][339]=83;
row_col[1][339]=154;
row_col[0][340]=84;
row_col[1][340]=202;
row_col[0][341]=85;
row_col[1][341]=191;
row_col[0][342]=86;
row_col[1][342]=131;
row_col[0][343]=87;
row_col[1][343]=169;
row_col[0][344]=88;
row_col[1][344]=161;
row_col[0][345]=89;
row_col[1][345]=180;
row_col[0][346]=90;
row_col[1][346]=232;
row_col[0][347]=91;
row_col[1][347]=245;
row_col[0][348]=92;
row_col[1][348]=216;
row_col[0][349]=93;
row_col[1][349]=192;
row_col[0][350]=94;
row_col[1][350]=143;
row_col[0][351]=95;
row_col[1][351]=164;
row_col[0][352]=96;
row_col[1][352]=252;
row_col[0][353]=97;
row_col[1][353]=176;
row_col[0][354]=98;
row_col[1][354]=233;
row_col[0][355]=99;
row_col[1][355]=137;
row_col[0][356]=100;
row_col[1][356]=157;
row_col[0][357]=101;
row_col[1][357]=188;
row_col[0][358]=102;
row_col[1][358]=220;
row_col[0][359]=103;
row_col[1][359]=130;
row_col[0][360]=104;
row_col[1][360]=206;
row_col[0][361]=105;
row_col[1][361]=237;
row_col[0][362]=106;
row_col[1][362]=229;
row_col[0][363]=107;
row_col[1][363]=146;
row_col[0][364]=108;
row_col[1][364]=201;
row_col[0][365]=109;
row_col[1][365]=249;
row_col[0][366]=110;
row_col[1][366]=241;
row_col[0][367]=111;
row_col[1][367]=151;
row_col[0][368]=112;
row_col[1][368]=210;
row_col[0][369]=113;
row_col[1][369]=235;
row_col[0][370]=114;
row_col[1][370]=193;
row_col[0][371]=115;
row_col[1][371]=160;
row_col[0][372]=116;
row_col[1][372]=222;
row_col[0][373]=117;
row_col[1][373]=199;
row_col[0][374]=118;
row_col[1][374]=171;
row_col[0][375]=119;
row_col[1][375]=207;
row_col[0][376]=120;
row_col[1][376]=179;
row_col[0][377]=121;
row_col[1][377]=218;
row_col[0][378]=122;
row_col[1][378]=166;
row_col[0][379]=123;
row_col[1][379]=240;
row_col[0][380]=124;
row_col[1][380]=227;
row_col[0][381]=125;
row_col[1][381]=185;
row_col[0][382]=126;
row_col[1][382]=204;
row_col[0][383]=127;
row_col[1][383]=213;



col_row[0][0]=0;
col_row[0][1]=1;
col_row[0][2]=256;
col_row[1][0]=1;
col_row[1][1]=2;
col_row[1][2]=257;
col_row[2][0]=2;
col_row[2][1]=3;
col_row[2][2]=258;
col_row[3][0]=3;
col_row[3][1]=4;
col_row[3][2]=259;
col_row[4][0]=4;
col_row[4][1]=5;
col_row[4][2]=260;
col_row[5][0]=5;
col_row[5][1]=6;
col_row[5][2]=261;
col_row[6][0]=6;
col_row[6][1]=7;
col_row[6][2]=262;
col_row[7][0]=7;
col_row[7][1]=8;
col_row[7][2]=263;
col_row[8][0]=8;
col_row[8][1]=9;
col_row[8][2]=264;
col_row[9][0]=9;
col_row[9][1]=10;
col_row[9][2]=265;
col_row[10][0]=10;
col_row[10][1]=11;
col_row[10][2]=266;
col_row[11][0]=11;
col_row[11][1]=12;
col_row[11][2]=267;
col_row[12][0]=12;
col_row[12][1]=13;
col_row[12][2]=268;
col_row[13][0]=13;
col_row[13][1]=14;
col_row[13][2]=269;
col_row[14][0]=14;
col_row[14][1]=15;
col_row[14][2]=270;
col_row[15][0]=15;
col_row[15][1]=16;
col_row[15][2]=271;
col_row[16][0]=16;
col_row[16][1]=17;
col_row[16][2]=272;
col_row[17][0]=17;
col_row[17][1]=18;
col_row[17][2]=273;
col_row[18][0]=18;
col_row[18][1]=19;
col_row[18][2]=274;
col_row[19][0]=19;
col_row[19][1]=20;
col_row[19][2]=275;
col_row[20][0]=20;
col_row[20][1]=21;
col_row[20][2]=276;
col_row[21][0]=21;
col_row[21][1]=22;
col_row[21][2]=277;
col_row[22][0]=22;
col_row[22][1]=23;
col_row[22][2]=278;
col_row[23][0]=23;
col_row[23][1]=24;
col_row[23][2]=279;
col_row[24][0]=24;
col_row[24][1]=25;
col_row[24][2]=280;
col_row[25][0]=25;
col_row[25][1]=26;
col_row[25][2]=281;
col_row[26][0]=26;
col_row[26][1]=27;
col_row[26][2]=282;
col_row[27][0]=27;
col_row[27][1]=28;
col_row[27][2]=283;
col_row[28][0]=28;
col_row[28][1]=29;
col_row[28][2]=284;
col_row[29][0]=29;
col_row[29][1]=30;
col_row[29][2]=285;
col_row[30][0]=30;
col_row[30][1]=31;
col_row[30][2]=286;
col_row[31][0]=31;
col_row[31][1]=32;
col_row[31][2]=287;
col_row[32][0]=32;
col_row[32][1]=33;
col_row[32][2]=288;
col_row[33][0]=33;
col_row[33][1]=34;
col_row[33][2]=289;
col_row[34][0]=34;
col_row[34][1]=35;
col_row[34][2]=290;
col_row[35][0]=35;
col_row[35][1]=36;
col_row[35][2]=291;
col_row[36][0]=36;
col_row[36][1]=37;
col_row[36][2]=292;
col_row[37][0]=37;
col_row[37][1]=38;
col_row[37][2]=293;
col_row[38][0]=38;
col_row[38][1]=39;
col_row[38][2]=294;
col_row[39][0]=39;
col_row[39][1]=40;
col_row[39][2]=295;
col_row[40][0]=40;
col_row[40][1]=41;
col_row[40][2]=296;
col_row[41][0]=41;
col_row[41][1]=42;
col_row[41][2]=297;
col_row[42][0]=42;
col_row[42][1]=43;
col_row[42][2]=298;
col_row[43][0]=43;
col_row[43][1]=44;
col_row[43][2]=299;
col_row[44][0]=44;
col_row[44][1]=45;
col_row[44][2]=300;
col_row[45][0]=45;
col_row[45][1]=46;
col_row[45][2]=301;
col_row[46][0]=46;
col_row[46][1]=47;
col_row[46][2]=302;
col_row[47][0]=47;
col_row[47][1]=48;
col_row[47][2]=303;
col_row[48][0]=48;
col_row[48][1]=49;
col_row[48][2]=304;
col_row[49][0]=49;
col_row[49][1]=50;
col_row[49][2]=305;
col_row[50][0]=50;
col_row[50][1]=51;
col_row[50][2]=306;
col_row[51][0]=51;
col_row[51][1]=52;
col_row[51][2]=307;
col_row[52][0]=52;
col_row[52][1]=53;
col_row[52][2]=308;
col_row[53][0]=53;
col_row[53][1]=54;
col_row[53][2]=309;
col_row[54][0]=54;
col_row[54][1]=55;
col_row[54][2]=310;
col_row[55][0]=55;
col_row[55][1]=56;
col_row[55][2]=311;
col_row[56][0]=56;
col_row[56][1]=57;
col_row[56][2]=312;
col_row[57][0]=57;
col_row[57][1]=58;
col_row[57][2]=313;
col_row[58][0]=58;
col_row[58][1]=59;
col_row[58][2]=314;
col_row[59][0]=59;
col_row[59][1]=60;
col_row[59][2]=315;
col_row[60][0]=60;
col_row[60][1]=61;
col_row[60][2]=316;
col_row[61][0]=61;
col_row[61][1]=62;
col_row[61][2]=317;
col_row[62][0]=62;
col_row[62][1]=63;
col_row[62][2]=318;
col_row[63][0]=63;
col_row[63][1]=64;
col_row[63][2]=319;
col_row[64][0]=64;
col_row[64][1]=65;
col_row[64][2]=320;
col_row[65][0]=65;
col_row[65][1]=66;
col_row[65][2]=321;
col_row[66][0]=66;
col_row[66][1]=67;
col_row[66][2]=322;
col_row[67][0]=67;
col_row[67][1]=68;
col_row[67][2]=323;
col_row[68][0]=68;
col_row[68][1]=69;
col_row[68][2]=324;
col_row[69][0]=69;
col_row[69][1]=70;
col_row[69][2]=325;
col_row[70][0]=70;
col_row[70][1]=71;
col_row[70][2]=326;
col_row[71][0]=71;
col_row[71][1]=72;
col_row[71][2]=327;
col_row[72][0]=72;
col_row[72][1]=73;
col_row[72][2]=328;
col_row[73][0]=73;
col_row[73][1]=74;
col_row[73][2]=329;
col_row[74][0]=74;
col_row[74][1]=75;
col_row[74][2]=330;
col_row[75][0]=75;
col_row[75][1]=76;
col_row[75][2]=331;
col_row[76][0]=76;
col_row[76][1]=77;
col_row[76][2]=332;
col_row[77][0]=77;
col_row[77][1]=78;
col_row[77][2]=333;
col_row[78][0]=78;
col_row[78][1]=79;
col_row[78][2]=334;
col_row[79][0]=79;
col_row[79][1]=80;
col_row[79][2]=335;
col_row[80][0]=80;
col_row[80][1]=81;
col_row[80][2]=336;
col_row[81][0]=81;
col_row[81][1]=82;
col_row[81][2]=337;
col_row[82][0]=82;
col_row[82][1]=83;
col_row[82][2]=338;
col_row[83][0]=83;
col_row[83][1]=84;
col_row[83][2]=339;
col_row[84][0]=84;
col_row[84][1]=85;
col_row[84][2]=340;
col_row[85][0]=85;
col_row[85][1]=86;
col_row[85][2]=341;
col_row[86][0]=86;
col_row[86][1]=87;
col_row[86][2]=342;
col_row[87][0]=87;
col_row[87][1]=88;
col_row[87][2]=343;
col_row[88][0]=88;
col_row[88][1]=89;
col_row[88][2]=344;
col_row[89][0]=89;
col_row[89][1]=90;
col_row[89][2]=345;
col_row[90][0]=90;
col_row[90][1]=91;
col_row[90][2]=346;
col_row[91][0]=91;
col_row[91][1]=92;
col_row[91][2]=347;
col_row[92][0]=92;
col_row[92][1]=93;
col_row[92][2]=348;
col_row[93][0]=93;
col_row[93][1]=94;
col_row[93][2]=349;
col_row[94][0]=94;
col_row[94][1]=95;
col_row[94][2]=350;
col_row[95][0]=95;
col_row[95][1]=96;
col_row[95][2]=351;
col_row[96][0]=96;
col_row[96][1]=97;
col_row[96][2]=352;
col_row[97][0]=97;
col_row[97][1]=98;
col_row[97][2]=353;
col_row[98][0]=98;
col_row[98][1]=99;
col_row[98][2]=354;
col_row[99][0]=99;
col_row[99][1]=100;
col_row[99][2]=355;
col_row[100][0]=100;
col_row[100][1]=101;
col_row[100][2]=356;
col_row[101][0]=101;
col_row[101][1]=102;
col_row[101][2]=357;
col_row[102][0]=102;
col_row[102][1]=103;
col_row[102][2]=358;
col_row[103][0]=103;
col_row[103][1]=104;
col_row[103][2]=359;
col_row[104][0]=104;
col_row[104][1]=105;
col_row[104][2]=360;
col_row[105][0]=105;
col_row[105][1]=106;
col_row[105][2]=361;
col_row[106][0]=106;
col_row[106][1]=107;
col_row[106][2]=362;
col_row[107][0]=107;
col_row[107][1]=108;
col_row[107][2]=363;
col_row[108][0]=108;
col_row[108][1]=109;
col_row[108][2]=364;
col_row[109][0]=109;
col_row[109][1]=110;
col_row[109][2]=365;
col_row[110][0]=110;
col_row[110][1]=111;
col_row[110][2]=366;
col_row[111][0]=111;
col_row[111][1]=112;
col_row[111][2]=367;
col_row[112][0]=112;
col_row[112][1]=113;
col_row[112][2]=368;
col_row[113][0]=113;
col_row[113][1]=114;
col_row[113][2]=369;
col_row[114][0]=114;
col_row[114][1]=115;
col_row[114][2]=370;
col_row[115][0]=115;
col_row[115][1]=116;
col_row[115][2]=371;
col_row[116][0]=116;
col_row[116][1]=117;
col_row[116][2]=372;
col_row[117][0]=117;
col_row[117][1]=118;
col_row[117][2]=373;
col_row[118][0]=118;
col_row[118][1]=119;
col_row[118][2]=374;
col_row[119][0]=119;
col_row[119][1]=120;
col_row[119][2]=375;
col_row[120][0]=120;
col_row[120][1]=121;
col_row[120][2]=376;
col_row[121][0]=121;
col_row[121][1]=122;
col_row[121][2]=377;
col_row[122][0]=122;
col_row[122][1]=123;
col_row[122][2]=378;
col_row[123][0]=123;
col_row[123][1]=124;
col_row[123][2]=379;
col_row[124][0]=124;
col_row[124][1]=125;
col_row[124][2]=380;
col_row[125][0]=125;
col_row[125][1]=126;
col_row[125][2]=381;
col_row[126][0]=126;
col_row[126][1]=127;
col_row[126][2]=382;
col_row[127][0]=0;
col_row[127][1]=127;
col_row[127][2]=383;
col_row[128][0]=128;
col_row[128][1]=129;
col_row[128][2]=334;
col_row[129][0]=129;
col_row[129][1]=130;
col_row[129][2]=268;
col_row[130][0]=130;
col_row[130][1]=131;
col_row[130][2]=359;
col_row[131][0]=131;
col_row[131][1]=132;
col_row[131][2]=342;
col_row[132][0]=132;
col_row[132][1]=133;
col_row[132][2]=257;
col_row[133][0]=133;
col_row[133][1]=134;
col_row[133][2]=320;
col_row[134][0]=134;
col_row[134][1]=135;
col_row[134][2]=297;
col_row[135][0]=135;
col_row[135][1]=136;
col_row[135][2]=264;
col_row[136][0]=136;
col_row[136][1]=137;
col_row[136][2]=326;
col_row[137][0]=137;
col_row[137][1]=138;
col_row[137][2]=355;
col_row[138][0]=138;
col_row[138][1]=139;
col_row[138][2]=289;
col_row[139][0]=139;
col_row[139][1]=140;
col_row[139][2]=314;
col_row[140][0]=140;
col_row[140][1]=141;
col_row[140][2]=336;
col_row[141][0]=141;
col_row[141][1]=142;
col_row[141][2]=256;
col_row[142][0]=142;
col_row[142][1]=143;
col_row[142][2]=277;
col_row[143][0]=143;
col_row[143][1]=144;
col_row[143][2]=350;
col_row[144][0]=144;
col_row[144][1]=145;
col_row[144][2]=307;
col_row[145][0]=145;
col_row[145][1]=146;
col_row[145][2]=266;
col_row[146][0]=146;
col_row[146][1]=147;
col_row[146][2]=363;
col_row[147][0]=147;
col_row[147][1]=148;
col_row[147][2]=300;
col_row[148][0]=148;
col_row[148][1]=149;
col_row[148][2]=259;
col_row[149][0]=149;
col_row[149][1]=150;
col_row[149][2]=325;
col_row[150][0]=150;
col_row[150][1]=151;
col_row[150][2]=293;
col_row[151][0]=151;
col_row[151][1]=152;
col_row[151][2]=367;
col_row[152][0]=152;
col_row[152][1]=153;
col_row[152][2]=269;
col_row[153][0]=153;
col_row[153][1]=154;
col_row[153][2]=278;
col_row[154][0]=154;
col_row[154][1]=155;
col_row[154][2]=339;
col_row[155][0]=155;
col_row[155][1]=156;
col_row[155][2]=322;
col_row[156][0]=156;
col_row[156][1]=157;
col_row[156][2]=261;
col_row[157][0]=157;
col_row[157][1]=158;
col_row[157][2]=356;
col_row[158][0]=158;
col_row[158][1]=159;
col_row[158][2]=305;
col_row[159][0]=159;
col_row[159][1]=160;
col_row[159][2]=272;
col_row[160][0]=160;
col_row[160][1]=161;
col_row[160][2]=371;
col_row[161][0]=161;
col_row[161][1]=162;
col_row[161][2]=344;
col_row[162][0]=162;
col_row[162][1]=163;
col_row[162][2]=315;
col_row[163][0]=163;
col_row[163][1]=164;
col_row[163][2]=294;
col_row[164][0]=164;
col_row[164][1]=165;
col_row[164][2]=351;
col_row[165][0]=165;
col_row[165][1]=166;
col_row[165][2]=262;
col_row[166][0]=166;
col_row[166][1]=167;
col_row[166][2]=378;
col_row[167][0]=167;
col_row[167][1]=168;
col_row[167][2]=288;
col_row[168][0]=168;
col_row[168][1]=169;
col_row[168][2]=330;
col_row[169][0]=169;
col_row[169][1]=170;
col_row[169][2]=343;
col_row[170][0]=170;
col_row[170][1]=171;
col_row[170][2]=279;
col_row[171][0]=171;
col_row[171][1]=172;
col_row[171][2]=374;
col_row[172][0]=172;
col_row[172][1]=173;
col_row[172][2]=265;
col_row[173][0]=173;
col_row[173][1]=174;
col_row[173][2]=337;
col_row[174][0]=174;
col_row[174][1]=175;
col_row[174][2]=285;
col_row[175][0]=175;
col_row[175][1]=176;
col_row[175][2]=302;
col_row[176][0]=176;
col_row[176][1]=177;
col_row[176][2]=353;
col_row[177][0]=177;
col_row[177][1]=178;
col_row[177][2]=270;
col_row[178][0]=178;
col_row[178][1]=179;
col_row[178][2]=319;
col_row[179][0]=179;
col_row[179][1]=180;
col_row[179][2]=376;
col_row[180][0]=180;
col_row[180][1]=181;
col_row[180][2]=345;
col_row[181][0]=181;
col_row[181][1]=182;
col_row[181][2]=308;
col_row[182][0]=182;
col_row[182][1]=183;
col_row[182][2]=338;
col_row[183][0]=183;
col_row[183][1]=184;
col_row[183][2]=327;
col_row[184][0]=184;
col_row[184][1]=185;
col_row[184][2]=273;
col_row[185][0]=185;
col_row[185][1]=186;
col_row[185][2]=381;
col_row[186][0]=186;
col_row[186][1]=187;
col_row[186][2]=299;
col_row[187][0]=187;
col_row[187][1]=188;
col_row[187][2]=280;
col_row[188][0]=188;
col_row[188][1]=189;
col_row[188][2]=357;
col_row[189][0]=189;
col_row[189][1]=190;
col_row[189][2]=292;
col_row[190][0]=190;
col_row[190][1]=191;
col_row[190][2]=311;
col_row[191][0]=191;
col_row[191][1]=192;
col_row[191][2]=341;
col_row[192][0]=192;
col_row[192][1]=193;
col_row[192][2]=349;
col_row[193][0]=193;
col_row[193][1]=194;
col_row[193][2]=370;
col_row[194][0]=194;
col_row[194][1]=195;
col_row[194][2]=321;
col_row[195][0]=195;
col_row[195][1]=196;
col_row[195][2]=282;
col_row[196][0]=196;
col_row[196][1]=197;
col_row[196][2]=335;
col_row[197][0]=197;
col_row[197][1]=198;
col_row[197][2]=306;
col_row[198][0]=198;
col_row[198][1]=199;
col_row[198][2]=295;
col_row[199][0]=199;
col_row[199][1]=200;
col_row[199][2]=373;
col_row[200][0]=200;
col_row[200][1]=201;
col_row[200][2]=287;
col_row[201][0]=201;
col_row[201][1]=202;
col_row[201][2]=364;
col_row[202][0]=202;
col_row[202][1]=203;
col_row[202][2]=340;
col_row[203][0]=203;
col_row[203][1]=204;
col_row[203][2]=318;
col_row[204][0]=204;
col_row[204][1]=205;
col_row[204][2]=382;
col_row[205][0]=205;
col_row[205][1]=206;
col_row[205][2]=304;
col_row[206][0]=206;
col_row[206][1]=207;
col_row[206][2]=360;
col_row[207][0]=207;
col_row[207][1]=208;
col_row[207][2]=375;
col_row[208][0]=208;
col_row[208][1]=209;
col_row[208][2]=313;
col_row[209][0]=209;
col_row[209][1]=210;
col_row[209][2]=298;
col_row[210][0]=210;
col_row[210][1]=211;
col_row[210][2]=368;
col_row[211][0]=211;
col_row[211][1]=212;
col_row[211][2]=286;
col_row[212][0]=212;
col_row[212][1]=213;
col_row[212][2]=323;
col_row[213][0]=213;
col_row[213][1]=214;
col_row[213][2]=383;
col_row[214][0]=214;
col_row[214][1]=215;
col_row[214][2]=309;
col_row[215][0]=215;
col_row[215][1]=216;
col_row[215][2]=331;
col_row[216][0]=216;
col_row[216][1]=217;
col_row[216][2]=348;
col_row[217][0]=217;
col_row[217][1]=218;
col_row[217][2]=296;
col_row[218][0]=218;
col_row[218][1]=219;
col_row[218][2]=377;
col_row[219][0]=219;
col_row[219][1]=220;
col_row[219][2]=284;
col_row[220][0]=220;
col_row[220][1]=221;
col_row[220][2]=358;
col_row[221][0]=221;
col_row[221][1]=222;
col_row[221][2]=328;
col_row[222][0]=222;
col_row[222][1]=223;
col_row[222][2]=372;
col_row[223][0]=223;
col_row[223][1]=224;
col_row[223][2]=276;
col_row[224][0]=224;
col_row[224][1]=225;
col_row[224][2]=301;
col_row[225][0]=225;
col_row[225][1]=226;
col_row[225][2]=316;
col_row[226][0]=226;
col_row[226][1]=227;
col_row[226][2]=332;
col_row[227][0]=227;
col_row[227][1]=228;
col_row[227][2]=380;
col_row[228][0]=228;
col_row[228][1]=229;
col_row[228][2]=291;
col_row[229][0]=229;
col_row[229][1]=230;
col_row[229][2]=362;
col_row[230][0]=230;
col_row[230][1]=231;
col_row[230][2]=283;
col_row[231][0]=231;
col_row[231][1]=232;
col_row[231][2]=274;
col_row[232][0]=232;
col_row[232][1]=233;
col_row[232][2]=346;
col_row[233][0]=233;
col_row[233][1]=234;
col_row[233][2]=354;
col_row[234][0]=234;
col_row[234][1]=235;
col_row[234][2]=333;
col_row[235][0]=235;
col_row[235][1]=236;
col_row[235][2]=369;
col_row[236][0]=236;
col_row[236][1]=237;
col_row[236][2]=263;
col_row[237][0]=237;
col_row[237][1]=238;
col_row[237][2]=361;
col_row[238][0]=238;
col_row[238][1]=239;
col_row[238][2]=271;
col_row[239][0]=239;
col_row[239][1]=240;
col_row[239][2]=310;
col_row[240][0]=240;
col_row[240][1]=241;
col_row[240][2]=379;
col_row[241][0]=241;
col_row[241][1]=242;
col_row[241][2]=366;
col_row[242][0]=242;
col_row[242][1]=243;
col_row[242][2]=281;
col_row[243][0]=243;
col_row[243][1]=244;
col_row[243][2]=260;
col_row[244][0]=244;
col_row[244][1]=245;
col_row[244][2]=317;
col_row[245][0]=245;
col_row[245][1]=246;
col_row[245][2]=347;
col_row[246][0]=246;
col_row[246][1]=247;
col_row[246][2]=267;
col_row[247][0]=247;
col_row[247][1]=248;
col_row[247][2]=290;
col_row[248][0]=248;
col_row[248][1]=249;
col_row[248][2]=303;
col_row[249][0]=249;
col_row[249][1]=250;
col_row[249][2]=365;
col_row[250][0]=250;
col_row[250][1]=251;
col_row[250][2]=329;
col_row[251][0]=251;
col_row[251][1]=252;
col_row[251][2]=258;
col_row[252][0]=252;
col_row[252][1]=253;
col_row[252][2]=352;
col_row[253][0]=253;
col_row[253][1]=254;
col_row[253][2]=312;
col_row[254][0]=254;
col_row[254][1]=255;
col_row[254][2]=275;
col_row[255][0]=128;
col_row[255][1]=255;
col_row[255][2]=324;


H[0][0]=1;
H[0][1]=8;
H[0][256]=9;
H[1][1]=9;
H[1][2]=1;
H[1][257]=8;
H[2][2]=8;
H[2][3]=1;
H[2][258]=9;
H[3][3]=1;
H[3][4]=1;
H[3][259]=8;
H[4][4]=8;
H[4][5]=9;
H[4][260]=1;
H[5][5]=1;
H[5][6]=11;
H[5][261]=1;
H[6][6]=1;
H[6][7]=1;
H[6][262]=10;
H[7][7]=1;
H[7][8]=14;
H[7][263]=8;
H[8][8]=1;
H[8][9]=9;
H[8][264]=8;
H[9][9]=3;
H[9][10]=1;
H[9][265]=11;
H[10][10]=1;
H[10][11]=1;
H[10][266]=11;
H[11][11]=10;
H[11][12]=1;
H[11][267]=1;
H[12][12]=8;
H[12][13]=9;
H[12][268]=1;
H[13][13]=1;
H[13][14]=10;
H[13][269]=1;
H[14][14]=1;
H[14][15]=8;
H[14][270]=1;
H[15][15]=1;
H[15][16]=1;
H[15][271]=8;
H[16][16]=1;
H[16][17]=1;
H[16][272]=10;
H[17][17]=8;
H[17][18]=1;
H[17][273]=7;
H[18][18]=8;
H[18][19]=9;
H[18][274]=1;
H[19][19]=8;
H[19][20]=1;
H[19][275]=1;
H[20][20]=1;
H[20][21]=8;
H[20][276]=14;
H[21][21]=9;
H[21][22]=8;
H[21][277]=1;
H[22][22]=1;
H[22][23]=9;
H[22][278]=8;
H[23][23]=1;
H[23][24]=9;
H[23][279]=9;
H[24][24]=8;
H[24][25]=9;
H[24][280]=1;
H[25][25]=11;
H[25][26]=1;
H[25][281]=1;
H[26][26]=11;
H[26][27]=1;
H[26][282]=1;
H[27][27]=10;
H[27][28]=1;
H[27][283]=1;
H[28][28]=8;
H[28][29]=1;
H[28][284]=1;
H[29][29]=1;
H[29][30]=3;
H[29][285]=11;
H[30][30]=11;
H[30][31]=3;
H[30][286]=1;
H[31][31]=8;
H[31][32]=1;
H[31][287]=14;
H[32][32]=8;
H[32][33]=1;
H[32][288]=9;
H[33][33]=1;
H[33][34]=10;
H[33][289]=1;
H[34][34]=1;
H[34][35]=1;
H[34][290]=8;
H[35][35]=11;
H[35][36]=3;
H[35][291]=1;
H[36][36]=1;
H[36][37]=1;
H[36][292]=10;
H[37][37]=8;
H[37][38]=9;
H[37][293]=1;
H[38][38]=1;
H[38][39]=1;
H[38][294]=11;
H[39][39]=10;
H[39][40]=1;
H[39][295]=1;
H[40][40]=7;
H[40][41]=1;
H[40][296]=7;
H[41][41]=8;
H[41][42]=1;
H[41][297]=1;
H[42][42]=1;
H[42][43]=10;
H[42][298]=1;
H[43][43]=1;
H[43][44]=9;
H[43][299]=8;
H[44][44]=8;
H[44][45]=9;
H[44][300]=1;
H[45][45]=1;
H[45][46]=1;
H[45][301]=8;
H[46][46]=1;
H[46][47]=1;
H[46][302]=10;
H[47][47]=10;
H[47][48]=1;
H[47][303]=1;
H[48][48]=11;
H[48][49]=1;
H[48][304]=1;
H[49][49]=1;
H[49][50]=8;
H[49][305]=9;
H[50][50]=1;
H[50][51]=11;
H[50][306]=3;
H[51][51]=3;
H[51][52]=1;
H[51][307]=11;
H[52][52]=8;
H[52][53]=1;
H[52][308]=1;
H[53][53]=1;
H[53][54]=11;
H[53][309]=1;
H[54][54]=8;
H[54][55]=1;
H[54][310]=1;
H[55][55]=1;
H[55][56]=9;
H[55][311]=8;
H[56][56]=1;
H[56][57]=8;
H[56][312]=1;
H[57][57]=8;
H[57][58]=9;
H[57][313]=1;
H[58][58]=8;
H[58][59]=1;
H[58][314]=7;
H[59][59]=1;
H[59][60]=10;
H[59][315]=1;
H[60][60]=9;
H[60][61]=1;
H[60][316]=8;
H[61][61]=10;
H[61][62]=1;
H[61][317]=1;
H[62][62]=8;
H[62][63]=14;
H[62][318]=1;
H[63][63]=1;
H[63][64]=10;
H[63][319]=1;
H[64][64]=1;
H[64][65]=10;
H[64][320]=1;
H[65][65]=8;
H[65][66]=1;
H[65][321]=1;
H[66][66]=1;
H[66][67]=8;
H[66][322]=9;
H[67][67]=8;
H[67][68]=1;
H[67][323]=1;
H[68][68]=1;
H[68][69]=11;
H[68][324]=3;
H[69][69]=8;
H[69][70]=7;
H[69][325]=1;
H[70][70]=1;
H[70][71]=1;
H[70][326]=8;
H[71][71]=8;
H[71][72]=14;
H[71][327]=1;
H[72][72]=11;
H[72][73]=1;
H[72][328]=1;
H[73][73]=1;
H[73][74]=3;
H[73][329]=11;
H[74][74]=1;
H[74][75]=1;
H[74][330]=10;
H[75][75]=1;
H[75][76]=8;
H[75][331]=1;
H[76][76]=1;
H[76][77]=1;
H[76][332]=11;
H[77][77]=1;
H[77][78]=10;
H[77][333]=1;
H[78][78]=11;
H[78][79]=1;
H[78][334]=1;
H[79][79]=9;
H[79][80]=6;
H[79][335]=1;
H[80][80]=1;
H[80][81]=11;
H[80][336]=1;
H[81][81]=1;
H[81][82]=10;
H[81][337]=1;
H[82][82]=9;
H[82][83]=1;
H[82][338]=1;
H[83][83]=1;
H[83][84]=1;
H[83][339]=9;
H[84][84]=1;
H[84][85]=8;
H[84][340]=1;
H[85][85]=7;
H[85][86]=7;
H[85][341]=1;
H[86][86]=1;
H[86][87]=10;
H[86][342]=1;
H[87][87]=8;
H[87][88]=1;
H[87][343]=9;
H[88][88]=1;
H[88][89]=8;
H[88][344]=14;
H[89][89]=8;
H[89][90]=1;
H[89][345]=1;
H[90][90]=1;
H[90][91]=9;
H[90][346]=1;
H[91][91]=14;
H[91][92]=8;
H[91][347]=1;
H[92][92]=1;
H[92][93]=1;
H[92][348]=8;
H[93][93]=1;
H[93][94]=6;
H[93][349]=9;
H[94][94]=1;
H[94][95]=10;
H[94][350]=1;
H[95][95]=1;
H[95][96]=8;
H[95][351]=1;
H[96][96]=10;
H[96][97]=1;
H[96][352]=1;
H[97][97]=1;
H[97][98]=1;
H[97][353]=10;
H[98][98]=1;
H[98][99]=1;
H[98][354]=8;
H[99][99]=1;
H[99][100]=8;
H[99][355]=1;
H[100][100]=8;
H[100][101]=14;
H[100][356]=1;
H[101][101]=11;
H[101][102]=1;
H[101][357]=3;
H[102][102]=1;
H[102][103]=1;
H[102][358]=11;
H[103][103]=1;
H[103][104]=10;
H[103][359]=1;
H[104][104]=9;
H[104][105]=1;
H[104][360]=9;
H[105][105]=11;
H[105][106]=1;
H[105][361]=1;
H[106][106]=8;
H[106][107]=7;
H[106][362]=1;
H[107][107]=1;
H[107][108]=8;
H[107][363]=7;
H[108][108]=1;
H[108][109]=8;
H[108][364]=14;
H[109][109]=1;
H[109][110]=1;
H[109][365]=10;
H[110][110]=8;
H[110][111]=1;
H[110][366]=1;
H[111][111]=1;
H[111][112]=11;
H[111][367]=1;
H[112][112]=8;
H[112][113]=1;
H[112][368]=9;
H[113][113]=1;
H[113][114]=8;
H[113][369]=9;
H[114][114]=1;
H[114][115]=1;
H[114][370]=10;
H[115][115]=10;
H[115][116]=1;
H[115][371]=1;
H[116][116]=1;
H[116][117]=1;
H[116][372]=11;
H[117][117]=14;
H[117][118]=8;
H[117][373]=1;
H[118][118]=1;
H[118][119]=8;
H[118][374]=7;
H[119][119]=10;
H[119][120]=1;
H[119][375]=1;
H[120][120]=11;
H[120][121]=1;
H[120][376]=3;
H[121][121]=1;
H[121][122]=9;
H[121][377]=1;
H[122][122]=1;
H[122][123]=9;
H[122][378]=8;
H[123][123]=11;
H[123][124]=1;
H[123][379]=1;
H[124][124]=8;
H[124][125]=1;
H[124][380]=1;
H[125][125]=1;
H[125][126]=8;
H[125][381]=1;
H[126][126]=1;
H[126][127]=10;
H[126][382]=1;
H[127][0]=1;
H[127][127]=10;
H[127][383]=1;
H[128][128]=1;
H[128][129]=9;
H[128][334]=8;
H[129][129]=8;
H[129][130]=9;
H[129][268]=1;
H[130][130]=3;
H[130][131]=11;
H[130][359]=1;
H[131][131]=1;
H[131][132]=9;
H[131][342]=8;
H[132][132]=1;
H[132][133]=1;
H[132][257]=11;
H[133][133]=1;
H[133][134]=8;
H[133][320]=14;
H[134][134]=1;
H[134][135]=3;
H[134][297]=11;
H[135][135]=8;
H[135][136]=1;
H[135][264]=14;
H[136][136]=9;
H[136][137]=8;
H[136][326]=1;
H[137][137]=11;
H[137][138]=1;
H[137][355]=1;
H[138][138]=11;
H[138][139]=1;
H[138][289]=3;
H[139][139]=11;
H[139][140]=1;
H[139][314]=1;
H[140][140]=1;
H[140][141]=8;
H[140][336]=1;
H[141][141]=1;
H[141][142]=1;
H[141][256]=10;
H[142][142]=1;
H[142][143]=1;
H[142][277]=8;
H[143][143]=10;
H[143][144]=1;
H[143][350]=1;
H[144][144]=11;
H[144][145]=1;
H[144][307]=1;
H[145][145]=1;
H[145][146]=1;
H[145][266]=8;
H[146][146]=11;
H[146][147]=1;
H[146][363]=1;
H[147][147]=11;
H[147][148]=3;
H[147][300]=1;
H[148][148]=1;
H[148][149]=8;
H[148][259]=9;
H[149][149]=1;
H[149][150]=8;
H[149][325]=9;
H[150][150]=1;
H[150][151]=10;
H[150][293]=1;
H[151][151]=1;
H[151][152]=8;
H[151][367]=1;
H[152][152]=1;
H[152][153]=10;
H[152][269]=1;
H[153][153]=1;
H[153][154]=1;
H[153][278]=10;
H[154][154]=8;
H[154][155]=14;
H[154][339]=1;
H[155][155]=1;
H[155][156]=10;
H[155][322]=1;
H[156][156]=1;
H[156][157]=1;
H[156][261]=11;
H[157][157]=1;
H[157][158]=1;
H[157][356]=10;
H[158][158]=10;
H[158][159]=1;
H[158][305]=1;
H[159][159]=6;
H[159][160]=9;
H[159][272]=1;
H[160][160]=1;
H[160][161]=10;
H[160][371]=1;
H[161][161]=8;
H[161][162]=1;
H[161][344]=1;
H[162][162]=1;
H[162][163]=10;
H[162][315]=1;
H[163][163]=14;
H[163][164]=1;
H[163][294]=8;
H[164][164]=1;
H[164][165]=6;
H[164][351]=9;
H[165][165]=9;
H[165][166]=1;
H[165][262]=1;
H[166][166]=1;
H[166][167]=11;
H[166][378]=1;
H[167][167]=7;
H[167][168]=1;
H[167][288]=6;
H[168][168]=9;
H[168][169]=6;
H[168][330]=1;
H[169][169]=1;
H[169][170]=1;
H[169][343]=10;
H[170][170]=1;
H[170][171]=1;
H[170][279]=8;
H[171][171]=1;
H[171][172]=10;
H[171][374]=1;
H[172][172]=1;
H[172][173]=8;
H[172][265]=1;
H[173][173]=1;
H[173][174]=1;
H[173][337]=8;
H[174][174]=9;
H[174][175]=1;
H[174][285]=8;
H[175][175]=1;
H[175][176]=1;
H[175][302]=10;
H[176][176]=9;
H[176][177]=1;
H[176][353]=9;
H[177][177]=1;
H[177][178]=1;
H[177][270]=11;
H[178][178]=1;
H[178][179]=8;
H[178][319]=1;
H[179][179]=7;
H[179][180]=7;
H[179][376]=1;
H[180][180]=1;
H[180][181]=1;
H[180][345]=9;
H[181][181]=1;
H[181][182]=1;
H[181][308]=8;
H[182][182]=9;
H[182][183]=1;
H[182][338]=8;
H[183][183]=8;
H[183][184]=9;
H[183][327]=1;
H[184][184]=1;
H[184][185]=7;
H[184][273]=7;
H[185][185]=1;
H[185][186]=8;
H[185][381]=1;
H[186][186]=1;
H[186][187]=1;
H[186][299]=10;
H[187][187]=9;
H[187][188]=1;
H[187][280]=1;
H[188][188]=9;
H[188][189]=8;
H[188][357]=1;
H[189][189]=1;
H[189][190]=10;
H[189][292]=1;
H[190][190]=1;
H[190][191]=11;
H[190][311]=1;
H[191][191]=1;
H[191][192]=1;
H[191][341]=10;
H[192][192]=8;
H[192][193]=1;
H[192][349]=1;
H[193][193]=1;
H[193][194]=8;
H[193][370]=14;
H[194][194]=1;
H[194][195]=1;
H[194][321]=11;
H[195][195]=1;
H[195][196]=9;
H[195][282]=8;
H[196][196]=11;
H[196][197]=1;
H[196][335]=1;
H[197][197]=1;
H[197][198]=1;
H[197][306]=10;
H[198][198]=1;
H[198][199]=11;
H[198][295]=3;
H[199][199]=1;
H[199][200]=10;
H[199][373]=1;
H[200][200]=1;
H[200][201]=10;
H[200][287]=1;
H[201][201]=6;
H[201][202]=9;
H[201][364]=1;
H[202][202]=7;
H[202][203]=1;
H[202][340]=6;
H[203][203]=9;
H[203][204]=8;
H[203][318]=1;
H[204][204]=1;
H[204][205]=8;
H[204][382]=1;
H[205][205]=1;
H[205][206]=9;
H[205][304]=8;
H[206][206]=8;
H[206][207]=1;
H[206][360]=7;
H[207][207]=1;
H[207][208]=11;
H[207][375]=3;
H[208][208]=1;
H[208][209]=8;
H[208][313]=9;
H[209][209]=1;
H[209][210]=1;
H[209][298]=11;
H[210][210]=9;
H[210][211]=1;
H[210][368]=8;
H[211][211]=1;
H[211][212]=10;
H[211][286]=1;
H[212][212]=1;
H[212][213]=11;
H[212][323]=1;
H[213][213]=8;
H[213][214]=1;
H[213][383]=7;
H[214][214]=1;
H[214][215]=8;
H[214][309]=9;
H[215][215]=10;
H[215][216]=1;
H[215][331]=1;
H[216][216]=1;
H[216][217]=11;
H[216][348]=1;
H[217][217]=8;
H[217][218]=1;
H[217][296]=1;
H[218][218]=7;
H[218][219]=7;
H[218][377]=1;
H[219][219]=1;
H[219][220]=1;
H[219][284]=8;
H[220][220]=7;
H[220][221]=7;
H[220][358]=1;
H[221][221]=9;
H[221][222]=1;
H[221][328]=9;
H[222][222]=1;
H[222][223]=8;
H[222][372]=1;
H[223][223]=1;
H[223][224]=1;
H[223][276]=9;
H[224][224]=6;
H[224][225]=9;
H[224][301]=1;
H[225][225]=1;
H[225][226]=6;
H[225][316]=7;
H[226][226]=9;
H[226][227]=6;
H[226][332]=1;
H[227][227]=1;
H[227][228]=10;
H[227][380]=1;
H[228][228]=1;
H[228][229]=1;
H[228][291]=9;
H[229][229]=10;
H[229][230]=1;
H[229][362]=1;
H[230][230]=1;
H[230][231]=9;
H[230][283]=8;
H[231][231]=1;
H[231][232]=1;
H[231][274]=9;
H[232][232]=1;
H[232][233]=6;
H[232][346]=9;
H[233][233]=1;
H[233][234]=1;
H[233][354]=10;
H[234][234]=1;
H[234][235]=9;
H[234][333]=1;
H[235][235]=1;
H[235][236]=1;
H[235][369]=8;
H[236][236]=1;
H[236][237]=9;
H[236][263]=1;
H[237][237]=1;
H[237][238]=1;
H[237][361]=8;
H[238][238]=9;
H[238][239]=1;
H[238][271]=1;
H[239][239]=1;
H[239][240]=1;
H[239][310]=10;
H[240][240]=1;
H[240][241]=9;
H[240][379]=8;
H[241][241]=1;
H[241][242]=11;
H[241][366]=3;
H[242][242]=7;
H[242][243]=7;
H[242][281]=1;
H[243][243]=11;
H[243][244]=1;
H[243][260]=3;
H[244][244]=9;
H[244][245]=1;
H[244][317]=9;
H[245][245]=1;
H[245][246]=11;
H[245][347]=1;
H[246][246]=1;
H[246][247]=11;
H[246][267]=1;
H[247][247]=8;
H[247][248]=1;
H[247][290]=1;
H[248][248]=1;
H[248][249]=1;
H[248][303]=11;
H[249][249]=7;
H[249][250]=7;
H[249][365]=1;
H[250][250]=9;
H[250][251]=9;
H[250][329]=1;
H[251][251]=3;
H[251][252]=11;
H[251][258]=1;
H[252][252]=6;
H[252][253]=1;
H[252][352]=7;
H[253][253]=9;
H[253][254]=1;
H[253][312]=9;
H[254][254]=9;
H[254][255]=1;
H[254][275]=8;
H[255][128]=8;
H[255][255]=1;
H[255][324]=1;




end

end



endmodule
