`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 24.01.2020 18:13:04
// Design Name:
// Module Name: test
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module simulation();
reg clk,reset;
//reg [5:0]in;
reg [5:0]beta;
wire[5:0]vout;
wire vout_en;
//integer handle1;
vn rgr(clk,reset,beta,vout,vout_en);
initial
clk=1'b0;
initial
reset=0;

initial
#110 reset=1;
initial
#120 reset=0;

initial
begin
#100 beta=6'd0;
#470 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd8;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd9;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd9;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd9;
#400 beta=6'd9;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd8;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd8;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd9;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd9;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd9;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd9;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd9;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd9;
#400 beta=6'd9;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd8;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd8;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd2;
#400 beta=6'd8;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd2;
#400 beta=6'd8;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd8;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd9;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd9;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd9;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd10;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd9;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd9;
#400 beta=6'd8;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd9;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd9;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd9;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd8;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd8;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd9;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd9;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd9;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd9;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd0;
#400 beta=6'd8;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd9;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd1;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd1;
#400 beta=6'd6;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd7;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd3;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd7;
#400 beta=6'd2;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd2;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd7;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd5;
#400 beta=6'd7;
#400 beta=6'd6;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd8;
#400 beta=6'd5;
#400 beta=6'd3;
#400 beta=6'd0;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd0;
#400 beta=6'd1;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd8;
#400 beta=6'd9;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd8;
#400 beta=6'd9;
#400 beta=6'd8;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd1;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd0;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd1;
#400 beta=6'd1;
#400 beta=6'd3;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd3;
#400 beta=6'd2;
#400 beta=6'd0;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd4;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd6;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd5;
#400 beta=6'd6;
#400 beta=6'd2;
#400 beta=6'd2;
#400 beta=6'd4;
#400 beta=6'd6;

end
initial
begin
forever
#200 clk=~clk;
end
endmodule
//create_clock -period 12.000 -name clk -waveform {0.000 6.000} -add [get_ports clk]
//create_clock -period 12.000 -name clk -waveform {0.000 6.000} -add [get_ports clk]
